
module b15 ( BE_n, \Address[29] , \Address[28] , \Address[27] , 
        \Address[26] , \Address[25] , \Address[24] , \Address[23] , 
        \Address[22] , \Address[21] , \Address[20] , \Address[19] , 
        \Address[18] , \Address[17] , \Address[16] , \Address[15] , 
        \Address[14] , \Address[13] , \Address[12] , \Address[11] , 
        \Address[10] , \Address[9] , \Address[8] , \Address[7] , \Address[6] , 
        \Address[5] , \Address[4] , \Address[3] , \Address[2] , \Address[1] , 
        \Address[0] , W_R_n, D_C_n, M_IO_n, ADS_n, \Datai[31] , 
        \Datai[30] , \Datai[29] , \Datai[28] , \Datai[27] , \Datai[26] , 
        \Datai[25] , \Datai[24] , \Datai[23] , \Datai[22] , \Datai[21] , 
        \Datai[20] , \Datai[19] , \Datai[18] , \Datai[17] , \Datai[16] , 
        \Datai[15] , \Datai[14] , \Datai[13] , \Datai[12] , \Datai[11] , 
        \Datai[10] , \Datai[9] , \Datai[8] , \Datai[7] , \Datai[6] , 
        \Datai[5] , \Datai[4] , \Datai[3] , \Datai[2] , \Datai[1] , \Datai[0] , 
        \Datao[31] , \Datao[30] , \Datao[29] , \Datao[28] , 
        \Datao[27] , \Datao[26] , \Datao[25] , \Datao[24] , \Datao[23] , 
        \Datao[22] , \Datao[21] , \Datao[20] , \Datao[19] , \Datao[18] , 
        \Datao[17] , \Datao[16] , \Datao[15] , \Datao[14] , \Datao[13] , 
        \Datao[12] , \Datao[11] , \Datao[10] , \Datao[9] , \Datao[8] , 
        \Datao[7] , \Datao[6] , \Datao[5] , \Datao[4] , \Datao[3] , \Datao[2] , 
        \Datao[1] , \Datao[0] , CLOCK, NA_n, BS16_n, READY_n, HOLD, RESET );
  output [3:0] BE_n;
  input \Datai[31] , \Datai[30] , \Datai[29] , \Datai[28] , \Datai[27] ,
         \Datai[26] , \Datai[25] , \Datai[24] , \Datai[23] , \Datai[22] ,
         \Datai[21] , \Datai[20] , \Datai[19] , \Datai[18] , \Datai[17] ,
         \Datai[16] , \Datai[15] , \Datai[14] , \Datai[13] , \Datai[12] ,
         \Datai[11] , \Datai[10] , \Datai[9] , \Datai[8] , \Datai[7] ,
         \Datai[6] , \Datai[5] , \Datai[4] , \Datai[3] , \Datai[2] ,
         \Datai[1] , \Datai[0] , CLOCK, NA_n, BS16_n, READY_n, HOLD, RESET;
  output \Address[29] , \Address[28] , \Address[27] , \Address[26] ,
         \Address[25] , \Address[24] , \Address[23] , \Address[22] ,
         \Address[21] , \Address[20] , \Address[19] , \Address[18] ,
         \Address[17] , \Address[16] , \Address[15] , \Address[14] ,
         \Address[13] , \Address[12] , \Address[11] , \Address[10] ,
         \Address[9] , \Address[8] , \Address[7] , \Address[6] , \Address[5] ,
         \Address[4] , \Address[3] , \Address[2] , \Address[1] , \Address[0] ,
         W_R_n, D_C_n, M_IO_n, ADS_n, \Datao[31] , \Datao[30] , \Datao[29] ,
         \Datao[28] , \Datao[27] , \Datao[26] , \Datao[25] , \Datao[24] ,
         \Datao[23] , \Datao[22] , \Datao[21] , \Datao[20] , \Datao[19] ,
         \Datao[18] , \Datao[17] , \Datao[16] , \Datao[15] , \Datao[14] ,
         \Datao[13] , \Datao[12] , \Datao[11] , \Datao[10] , \Datao[9] ,
         \Datao[8] , \Datao[7] , \Datao[6] , \Datao[5] , \Datao[4] ,
         \Datao[3] , \Datao[2] , \Datao[1] , \Datao[0] ;
  wire   StateBS16, RequestPending, MemoryFetch, ReadRequest, CodeFetch,
         \InstQueue[15][7] , \InstQueue[15][6] , \InstQueue[15][5] ,
         \InstQueue[15][4] , \InstQueue[15][3] , \InstQueue[15][2] ,
         \InstQueue[15][1] , \InstQueue[15][0] , \InstQueue[14][7] ,
         \InstQueue[14][6] , \InstQueue[14][5] , \InstQueue[14][4] ,
         \InstQueue[14][3] , \InstQueue[14][2] , \InstQueue[14][1] ,
         \InstQueue[14][0] , \InstQueue[13][7] , \InstQueue[13][6] ,
         \InstQueue[13][5] , \InstQueue[13][4] , \InstQueue[13][3] ,
         \InstQueue[13][2] , \InstQueue[13][1] , \InstQueue[13][0] ,
         \InstQueue[12][7] , \InstQueue[12][6] , \InstQueue[12][5] ,
         \InstQueue[12][4] , \InstQueue[12][3] , \InstQueue[12][2] ,
         \InstQueue[12][1] , \InstQueue[12][0] , \InstQueue[11][7] ,
         \InstQueue[11][6] , \InstQueue[11][5] , \InstQueue[11][4] ,
         \InstQueue[11][3] , \InstQueue[11][2] , \InstQueue[11][1] ,
         \InstQueue[11][0] , \InstQueue[10][7] , \InstQueue[10][6] ,
         \InstQueue[10][5] , \InstQueue[10][4] , \InstQueue[10][3] ,
         \InstQueue[10][2] , \InstQueue[10][1] , \InstQueue[10][0] ,
         \InstQueue[9][7] , \InstQueue[9][6] , \InstQueue[9][5] ,
         \InstQueue[9][4] , \InstQueue[9][3] , \InstQueue[9][2] ,
         \InstQueue[9][1] , \InstQueue[9][0] , \InstQueue[8][7] ,
         \InstQueue[8][6] , \InstQueue[8][5] , \InstQueue[8][4] ,
         \InstQueue[8][3] , \InstQueue[8][2] , \InstQueue[8][1] ,
         \InstQueue[8][0] , \InstQueue[7][7] , \InstQueue[7][6] ,
         \InstQueue[7][5] , \InstQueue[7][4] , \InstQueue[7][3] ,
         \InstQueue[7][2] , \InstQueue[7][1] , \InstQueue[7][0] ,
         \InstQueue[6][7] , \InstQueue[6][6] , \InstQueue[6][5] ,
         \InstQueue[6][4] , \InstQueue[6][3] , \InstQueue[6][2] ,
         \InstQueue[6][1] , \InstQueue[6][0] , \InstQueue[5][7] ,
         \InstQueue[5][6] , \InstQueue[5][5] , \InstQueue[5][4] ,
         \InstQueue[5][3] , \InstQueue[5][2] , \InstQueue[5][1] ,
         \InstQueue[5][0] , \InstQueue[4][7] , \InstQueue[4][6] ,
         \InstQueue[4][5] , \InstQueue[4][4] , \InstQueue[4][3] ,
         \InstQueue[4][2] , \InstQueue[4][1] , \InstQueue[4][0] ,
         \InstQueue[3][7] , \InstQueue[3][6] , \InstQueue[3][5] ,
         \InstQueue[3][4] , \InstQueue[3][3] , \InstQueue[3][2] ,
         \InstQueue[3][1] , \InstQueue[3][0] , \InstQueue[2][7] ,
         \InstQueue[2][6] , \InstQueue[2][5] , \InstQueue[2][4] ,
         \InstQueue[2][3] , \InstQueue[2][2] , \InstQueue[2][1] ,
         \InstQueue[2][0] , \InstQueue[1][7] , \InstQueue[1][6] ,
         \InstQueue[1][5] , \InstQueue[1][4] , \InstQueue[1][3] ,
         \InstQueue[1][2] , \InstQueue[1][1] , \InstQueue[1][0] , More, Flush,
         N1009, N1351, N1753, N1868, N1989, N2884, N3678, N4154, N4186, N4187,
         N4188, \C1/DATA1_29 , \C1/DATA1_28 , \C1/DATA1_27 , \C1/DATA1_26 ,
         \C1/DATA1_25 , \C1/DATA1_24 , \C1/DATA1_23 , \C1/DATA1_22 ,
         \C1/DATA1_21 , \C1/DATA1_20 , \C1/DATA1_19 , \C1/DATA1_18 ,
         \C1/DATA1_17 , \C1/DATA1_16 , \C1/DATA2_30 , \C1/DATA2_29 ,
         \C1/DATA2_28 , \C1/DATA2_27 , \C1/DATA2_26 , \C1/DATA2_25 ,
         \C1/DATA2_24 , \C1/DATA2_23 , \C1/DATA2_22 , \C1/DATA2_21 ,
         \C1/DATA2_20 , \C1/DATA2_19 , \C1/DATA2_18 , \C1/DATA2_17 ,
         \C1/DATA2_16 , \C1/DATA2_15 , \C1/DATA2_14 , \C1/DATA2_13 ,
         \C1/DATA2_12 , \C1/DATA2_11 , \C1/DATA2_10 , \C1/DATA2_9 ,
         \C1/DATA2_8 , \C1/DATA2_7 , \C1/DATA2_6 , \C1/DATA2_5 , \C1/DATA2_4 ,
         \C1/DATA2_3 , \C1/DATA2_2 , \C1/DATA2_1 , \C1/DATA2_0 , n1660, n1661,
         n1662, n1663, n1664, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, \DP_OP_560J1_146_4463/n14 ,
         \DP_OP_560J1_146_4463/n13 , \DP_OP_560J1_146_4463/n12 ,
         \DP_OP_560J1_146_4463/n11 , \DP_OP_560J1_146_4463/n10 ,
         \DP_OP_560J1_146_4463/n9 , \DP_OP_560J1_146_4463/n8 ,
         \DP_OP_560J1_146_4463/n7 , \DP_OP_560J1_146_4463/n6 ,
         \DP_OP_560J1_146_4463/n5 , \DP_OP_560J1_146_4463/n4 ,
         \DP_OP_560J1_146_4463/n3 , \DP_OP_560J1_146_4463/n2 ,
         \DP_OP_560J1_146_4463/n1 , \DP_OP_469J1_133_8416/n123 ,
         \DP_OP_469J1_133_8416/n122 , \DP_OP_469J1_133_8416/n121 ,
         \DP_OP_469J1_133_8416/n120 , \DP_OP_469J1_133_8416/n119 ,
         \DP_OP_469J1_133_8416/n118 , \DP_OP_469J1_133_8416/n117 ,
         \DP_OP_469J1_133_8416/n116 , n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291;
  wire   [29:0] Address;
  wire   [31:0] Datai;
  wire   [31:0] Datao;
  wire   [2:0] State;
  wire   [31:0] DataWidth;
  wire   [31:0] rEIP;
  wire   [3:0] ByteEnable;
  wire   [3:0] State2;
  wire   [4:0] InstQueueRd_Addr;
  wire   [31:0] InstAddrPointer;
  wire   [31:0] PhyAddrPointer;
  wire   [31:0] EAX;
  wire   [31:0] EBX;
  assign \Datao[31]  = 1'b0;

  DFFARX1 RequestPending_reg ( .D(n2077), .CLK(CLOCK), .RSTB(n5284), .Q(
        RequestPending) );
  DFFARX1 \State_reg[2]  ( .D(n2074), .CLK(CLOCK), .RSTB(n5282), .Q(State[2]), 
        .QN(n5207) );
  DFFARX1 \State_reg[1]  ( .D(n2075), .CLK(CLOCK), .RSTB(n5277), .Q(State[1]), 
        .QN(n5178) );
  DFFARX1 \State_reg[0]  ( .D(n2076), .CLK(CLOCK), .RSTB(n5282), .Q(State[0]), 
        .QN(n5202) );
  DFFARX1 \Address_reg[0]  ( .D(n1702), .CLK(CLOCK), .RSTB(n5290), .Q(
        Address[0]) );
  DFFARX1 \Address_reg[1]  ( .D(n1701), .CLK(CLOCK), .RSTB(n5291), .Q(
        Address[1]) );
  DFFARX1 \Address_reg[2]  ( .D(n1700), .CLK(CLOCK), .RSTB(n5279), .Q(
        Address[2]) );
  DFFARX1 \Address_reg[3]  ( .D(n1699), .CLK(CLOCK), .RSTB(n5286), .Q(
        Address[3]) );
  DFFARX1 \Address_reg[4]  ( .D(n1698), .CLK(CLOCK), .RSTB(n5284), .Q(
        Address[4]) );
  DFFARX1 \Address_reg[5]  ( .D(n1697), .CLK(CLOCK), .RSTB(n5284), .Q(
        Address[5]) );
  DFFARX1 \Address_reg[6]  ( .D(n1696), .CLK(CLOCK), .RSTB(n5285), .Q(
        Address[6]) );
  DFFARX1 \Address_reg[7]  ( .D(n1695), .CLK(CLOCK), .RSTB(n5288), .Q(
        Address[7]) );
  DFFARX1 \Address_reg[8]  ( .D(n1694), .CLK(CLOCK), .RSTB(n5278), .Q(
        Address[8]) );
  DFFARX1 \Address_reg[9]  ( .D(n1693), .CLK(CLOCK), .RSTB(n5283), .Q(
        Address[9]) );
  DFFARX1 \Address_reg[10]  ( .D(n1692), .CLK(CLOCK), .RSTB(n5287), .Q(
        Address[10]) );
  DFFARX1 \Address_reg[11]  ( .D(n1691), .CLK(CLOCK), .RSTB(n5282), .Q(
        Address[11]) );
  DFFARX1 \Address_reg[12]  ( .D(n1690), .CLK(CLOCK), .RSTB(n5278), .Q(
        Address[12]) );
  DFFARX1 \Address_reg[13]  ( .D(n1689), .CLK(CLOCK), .RSTB(n5277), .Q(
        Address[13]) );
  DFFARX1 \Address_reg[14]  ( .D(n1688), .CLK(CLOCK), .RSTB(n5288), .Q(
        Address[14]) );
  DFFARX1 \Address_reg[15]  ( .D(n1687), .CLK(CLOCK), .RSTB(n5278), .Q(
        Address[15]) );
  DFFARX1 \Address_reg[16]  ( .D(n1686), .CLK(CLOCK), .RSTB(n5277), .Q(
        Address[16]) );
  DFFARX1 \Address_reg[17]  ( .D(n1685), .CLK(CLOCK), .RSTB(n5279), .Q(
        Address[17]) );
  DFFARX1 \Address_reg[18]  ( .D(n1684), .CLK(CLOCK), .RSTB(n5284), .Q(
        Address[18]) );
  DFFARX1 \Address_reg[19]  ( .D(n1683), .CLK(CLOCK), .RSTB(n5280), .Q(
        Address[19]) );
  DFFARX1 \Address_reg[20]  ( .D(n1682), .CLK(CLOCK), .RSTB(n5281), .Q(
        Address[20]) );
  DFFARX1 \Address_reg[21]  ( .D(n1681), .CLK(CLOCK), .RSTB(n5286), .Q(
        Address[21]) );
  DFFARX1 \Address_reg[22]  ( .D(n1680), .CLK(CLOCK), .RSTB(n5277), .Q(
        Address[22]) );
  DFFARX1 \Address_reg[23]  ( .D(n1679), .CLK(CLOCK), .RSTB(n5288), .Q(
        Address[23]) );
  DFFARX1 \Address_reg[24]  ( .D(n1678), .CLK(CLOCK), .RSTB(n5288), .Q(
        Address[24]) );
  DFFARX1 \Address_reg[25]  ( .D(n1677), .CLK(CLOCK), .RSTB(n5288), .Q(
        Address[25]) );
  DFFARX1 \Address_reg[26]  ( .D(n1676), .CLK(CLOCK), .RSTB(n5288), .Q(
        Address[26]) );
  DFFARX1 \Address_reg[27]  ( .D(n1675), .CLK(CLOCK), .RSTB(n5288), .Q(
        Address[27]) );
  DFFARX1 \Address_reg[28]  ( .D(n1674), .CLK(CLOCK), .RSTB(n5288), .Q(
        Address[28]) );
  DFFARX1 \Address_reg[29]  ( .D(n1673), .CLK(CLOCK), .RSTB(n5288), .Q(
        Address[29]) );
  DFFARX1 \DataWidth_reg[0]  ( .D(n1704), .CLK(CLOCK), .RSTB(n5280), .Q(
        DataWidth[0]), .QN(n5250) );
  DFFARX1 StateBS16_reg ( .D(n2073), .CLK(CLOCK), .RSTB(n5288), .Q(StateBS16), 
        .QN(n5203) );
  DFFARX1 \State2_reg[2]  ( .D(n2066), .CLK(CLOCK), .RSTB(n5285), .Q(State2[2]), .QN(n5236) );
  DFFARX1 Flush_reg ( .D(n2030), .CLK(CLOCK), .RSTB(n5287), .Q(Flush), .QN(
        n5208) );
  DFFARX1 \EAX_reg[0]  ( .D(n1990), .CLK(CLOCK), .RSTB(n5287), .Q(EAX[0]) );
  DFFARX1 \EAX_reg[1]  ( .D(n1989), .CLK(CLOCK), .RSTB(n5283), .Q(EAX[1]) );
  DFFARX1 \EAX_reg[2]  ( .D(n1988), .CLK(CLOCK), .RSTB(n5289), .Q(EAX[2]) );
  DFFARX1 \EAX_reg[3]  ( .D(n1987), .CLK(CLOCK), .RSTB(n5286), .Q(EAX[3]) );
  DFFARX1 \EAX_reg[4]  ( .D(n1986), .CLK(CLOCK), .RSTB(n5285), .Q(EAX[4]) );
  DFFARX1 \EAX_reg[5]  ( .D(n1985), .CLK(CLOCK), .RSTB(n5284), .Q(EAX[5]) );
  DFFARX1 \EAX_reg[6]  ( .D(n1984), .CLK(CLOCK), .RSTB(n5286), .Q(EAX[6]) );
  DFFARX1 \EAX_reg[7]  ( .D(n1983), .CLK(CLOCK), .RSTB(n5291), .Q(EAX[7]) );
  DFFARX1 \EAX_reg[8]  ( .D(n1982), .CLK(CLOCK), .RSTB(n5290), .Q(EAX[8]) );
  DFFARX1 \EAX_reg[9]  ( .D(n1981), .CLK(CLOCK), .RSTB(n5283), .Q(EAX[9]) );
  DFFARX1 \EAX_reg[10]  ( .D(n1980), .CLK(CLOCK), .RSTB(n5279), .Q(EAX[10]) );
  DFFARX1 \EAX_reg[11]  ( .D(n1979), .CLK(CLOCK), .RSTB(n5277), .Q(EAX[11]) );
  DFFARX1 \EAX_reg[12]  ( .D(n1978), .CLK(CLOCK), .RSTB(n5287), .Q(EAX[12]) );
  DFFARX1 \EAX_reg[13]  ( .D(n1977), .CLK(CLOCK), .RSTB(n5277), .Q(EAX[13]) );
  DFFARX1 \EAX_reg[14]  ( .D(n1976), .CLK(CLOCK), .RSTB(n5278), .Q(EAX[14]) );
  DFFARX1 \EAX_reg[15]  ( .D(n1975), .CLK(CLOCK), .RSTB(n5278), .Q(EAX[15]) );
  DFFARX1 \EAX_reg[16]  ( .D(n1974), .CLK(CLOCK), .RSTB(n5281), .Q(EAX[16]) );
  DFFARX1 \EAX_reg[17]  ( .D(n1973), .CLK(CLOCK), .RSTB(n5281), .Q(EAX[17]) );
  DFFARX1 \EAX_reg[18]  ( .D(n1972), .CLK(CLOCK), .RSTB(n5280), .Q(EAX[18]) );
  DFFARX1 \EAX_reg[19]  ( .D(n1971), .CLK(CLOCK), .RSTB(n5286), .Q(EAX[19]) );
  DFFARX1 \EAX_reg[20]  ( .D(n1970), .CLK(CLOCK), .RSTB(n5279), .Q(EAX[20]) );
  DFFARX1 \EAX_reg[21]  ( .D(n1969), .CLK(CLOCK), .RSTB(n5277), .Q(EAX[21]) );
  DFFARX1 \EAX_reg[22]  ( .D(n1968), .CLK(CLOCK), .RSTB(n5278), .Q(EAX[22]) );
  DFFARX1 \EAX_reg[23]  ( .D(n1967), .CLK(CLOCK), .RSTB(n5289), .Q(EAX[23]) );
  DFFARX1 \EAX_reg[24]  ( .D(n1966), .CLK(CLOCK), .RSTB(n5281), .Q(EAX[24]) );
  DFFARX1 \EAX_reg[25]  ( .D(n1965), .CLK(CLOCK), .RSTB(n5282), .Q(EAX[25]) );
  DFFARX1 \EAX_reg[26]  ( .D(n1964), .CLK(CLOCK), .RSTB(n5280), .Q(EAX[26]) );
  DFFARX1 \EAX_reg[27]  ( .D(n1963), .CLK(CLOCK), .RSTB(n5282), .Q(EAX[27]) );
  DFFARX1 \EAX_reg[28]  ( .D(n1962), .CLK(CLOCK), .RSTB(n5288), .Q(EAX[28]) );
  DFFARX1 \EAX_reg[29]  ( .D(n1961), .CLK(CLOCK), .RSTB(n5291), .Q(EAX[29]) );
  DFFARX1 \EAX_reg[30]  ( .D(n1960), .CLK(CLOCK), .RSTB(n5287), .Q(EAX[30]), 
        .QN(n5262) );
  DFFARX1 \EAX_reg[31]  ( .D(n1959), .CLK(CLOCK), .RSTB(n5283), .Q(EAX[31]) );
  DFFARX1 More_reg ( .D(n2029), .CLK(CLOCK), .RSTB(n5283), .Q(More) );
  DFFARX1 \uWord_reg[0]  ( .D(n1958), .CLK(CLOCK), .RSTB(n5277), .Q(
        \C1/DATA2_16 ) );
  DFFARX1 \uWord_reg[1]  ( .D(n1957), .CLK(CLOCK), .RSTB(n5287), .Q(
        \C1/DATA2_17 ) );
  DFFARX1 \uWord_reg[2]  ( .D(n1956), .CLK(CLOCK), .RSTB(n5282), .Q(
        \C1/DATA2_18 ) );
  DFFARX1 \uWord_reg[3]  ( .D(n1955), .CLK(CLOCK), .RSTB(n5285), .Q(
        \C1/DATA2_19 ) );
  DFFARX1 \uWord_reg[4]  ( .D(n1954), .CLK(CLOCK), .RSTB(n5290), .Q(
        \C1/DATA2_20 ) );
  DFFARX1 \uWord_reg[5]  ( .D(n1953), .CLK(CLOCK), .RSTB(n5284), .Q(
        \C1/DATA2_21 ) );
  DFFARX1 \uWord_reg[6]  ( .D(n1952), .CLK(CLOCK), .RSTB(n5278), .Q(
        \C1/DATA2_22 ) );
  DFFARX1 \uWord_reg[7]  ( .D(n1951), .CLK(CLOCK), .RSTB(n5282), .Q(
        \C1/DATA2_23 ) );
  DFFARX1 \uWord_reg[8]  ( .D(n1950), .CLK(CLOCK), .RSTB(n5289), .Q(
        \C1/DATA2_24 ) );
  DFFARX1 \uWord_reg[9]  ( .D(n1949), .CLK(CLOCK), .RSTB(n5278), .Q(
        \C1/DATA2_25 ) );
  DFFARX1 \uWord_reg[10]  ( .D(n1948), .CLK(CLOCK), .RSTB(n5282), .Q(
        \C1/DATA2_26 ) );
  DFFARX1 \uWord_reg[11]  ( .D(n1947), .CLK(CLOCK), .RSTB(n5280), .Q(
        \C1/DATA2_27 ) );
  DFFARX1 \uWord_reg[12]  ( .D(n1946), .CLK(CLOCK), .RSTB(n5281), .Q(
        \C1/DATA2_28 ) );
  DFFARX1 \uWord_reg[13]  ( .D(n1945), .CLK(CLOCK), .RSTB(n5280), .Q(
        \C1/DATA2_29 ) );
  DFFARX1 \uWord_reg[14]  ( .D(n1944), .CLK(CLOCK), .RSTB(n5291), .Q(
        \C1/DATA2_30 ) );
  DFFARX1 \lWord_reg[0]  ( .D(n1943), .CLK(CLOCK), .RSTB(n5285), .Q(
        \C1/DATA2_0 ) );
  DFFARX1 \lWord_reg[1]  ( .D(n1942), .CLK(CLOCK), .RSTB(n5284), .Q(
        \C1/DATA2_1 ) );
  DFFARX1 \lWord_reg[2]  ( .D(n1941), .CLK(CLOCK), .RSTB(n5286), .Q(
        \C1/DATA2_2 ) );
  DFFARX1 \lWord_reg[3]  ( .D(n1940), .CLK(CLOCK), .RSTB(n5291), .Q(
        \C1/DATA2_3 ) );
  DFFARX1 \lWord_reg[4]  ( .D(n1939), .CLK(CLOCK), .RSTB(n5290), .Q(
        \C1/DATA2_4 ) );
  DFFARX1 \lWord_reg[5]  ( .D(n1938), .CLK(CLOCK), .RSTB(n5285), .Q(
        \C1/DATA2_5 ) );
  DFFARX1 \lWord_reg[6]  ( .D(n1937), .CLK(CLOCK), .RSTB(n5279), .Q(
        \C1/DATA2_6 ) );
  DFFARX1 \lWord_reg[7]  ( .D(n1936), .CLK(CLOCK), .RSTB(n5289), .Q(
        \C1/DATA2_7 ) );
  DFFARX1 \lWord_reg[8]  ( .D(n1935), .CLK(CLOCK), .RSTB(n5280), .Q(
        \C1/DATA2_8 ) );
  DFFARX1 \lWord_reg[9]  ( .D(n1934), .CLK(CLOCK), .RSTB(n5279), .Q(
        \C1/DATA2_9 ) );
  DFFARX1 \lWord_reg[10]  ( .D(n1933), .CLK(CLOCK), .RSTB(n5289), .Q(
        \C1/DATA2_10 ) );
  DFFARX1 \lWord_reg[11]  ( .D(n1932), .CLK(CLOCK), .RSTB(n5281), .Q(
        \C1/DATA2_11 ) );
  DFFARX1 \lWord_reg[12]  ( .D(n1931), .CLK(CLOCK), .RSTB(n5280), .Q(
        \C1/DATA2_12 ) );
  DFFARX1 \lWord_reg[13]  ( .D(n1930), .CLK(CLOCK), .RSTB(n5285), .Q(
        \C1/DATA2_13 ) );
  DFFARX1 \lWord_reg[14]  ( .D(n1929), .CLK(CLOCK), .RSTB(n5279), .Q(
        \C1/DATA2_14 ) );
  DFFARX1 \lWord_reg[15]  ( .D(n1928), .CLK(CLOCK), .RSTB(n5277), .Q(
        \C1/DATA2_15 ) );
  DFFARX1 \State2_reg[0]  ( .D(n2068), .CLK(CLOCK), .RSTB(n5279), .Q(State2[0]), .QN(n5176) );
  DFFARX1 \State2_reg[1]  ( .D(n2067), .CLK(CLOCK), .RSTB(n5279), .Q(State2[1]), .QN(n5242) );
  DFFARX1 \State2_reg[3]  ( .D(n2072), .CLK(CLOCK), .RSTB(n5281), .Q(State2[3]), .QN(n5179) );
  DFFARX1 CodeFetch_reg ( .D(n2034), .CLK(CLOCK), .RSTB(n5280), .Q(CodeFetch), 
        .QN(n5197) );
  DFFARX1 D_C_n_reg ( .D(n1670), .CLK(CLOCK), .RSTB(n5279), .Q(D_C_n) );
  DFFARX1 MemoryFetch_reg ( .D(n2032), .CLK(CLOCK), .RSTB(n5277), .Q(
        MemoryFetch) );
  DFFARX1 M_IO_n_reg ( .D(n1672), .CLK(CLOCK), .RSTB(n5278), .Q(M_IO_n) );
  DFFARX1 ReadRequest_reg ( .D(n2031), .CLK(CLOCK), .RSTB(n5288), .Q(
        ReadRequest), .QN(n5251) );
  DFFARX1 W_R_n_reg ( .D(n1671), .CLK(CLOCK), .RSTB(n5279), .Q(W_R_n) );
  DFFARX1 \InstQueueWr_Addr_reg[0]  ( .D(n2024), .CLK(CLOCK), .RSTB(n5282), 
        .Q(N1351), .QN(n5199) );
  DFFARX1 \Datao_reg[0]  ( .D(n1927), .CLK(CLOCK), .RSTB(n5288), .Q(Datao[0])
         );
  DFFARX1 \Datao_reg[1]  ( .D(n1926), .CLK(CLOCK), .RSTB(n5290), .Q(Datao[1])
         );
  DFFARX1 \Datao_reg[2]  ( .D(n1925), .CLK(CLOCK), .RSTB(n5287), .Q(Datao[2])
         );
  DFFARX1 \Datao_reg[3]  ( .D(n1924), .CLK(CLOCK), .RSTB(n5277), .Q(Datao[3])
         );
  DFFARX1 \Datao_reg[4]  ( .D(n1923), .CLK(CLOCK), .RSTB(n5277), .Q(Datao[4])
         );
  DFFARX1 \Datao_reg[5]  ( .D(n1922), .CLK(CLOCK), .RSTB(n5277), .Q(Datao[5])
         );
  DFFARX1 \Datao_reg[6]  ( .D(n1921), .CLK(CLOCK), .RSTB(n5277), .Q(Datao[6])
         );
  DFFARX1 \Datao_reg[7]  ( .D(n1920), .CLK(CLOCK), .RSTB(n5277), .Q(Datao[7])
         );
  DFFARX1 \Datao_reg[8]  ( .D(n1919), .CLK(CLOCK), .RSTB(n5277), .Q(Datao[8])
         );
  DFFARX1 \Datao_reg[9]  ( .D(n1918), .CLK(CLOCK), .RSTB(n5277), .Q(Datao[9])
         );
  DFFARX1 \Datao_reg[10]  ( .D(n1917), .CLK(CLOCK), .RSTB(n5277), .Q(Datao[10]) );
  DFFARX1 \Datao_reg[11]  ( .D(n1916), .CLK(CLOCK), .RSTB(n5277), .Q(Datao[11]) );
  DFFARX1 \Datao_reg[12]  ( .D(n1915), .CLK(CLOCK), .RSTB(n5277), .Q(Datao[12]) );
  DFFARX1 \Datao_reg[13]  ( .D(n1914), .CLK(CLOCK), .RSTB(n5277), .Q(Datao[13]) );
  DFFARX1 \Datao_reg[14]  ( .D(n1913), .CLK(CLOCK), .RSTB(n5277), .Q(Datao[14]) );
  DFFARX1 \Datao_reg[15]  ( .D(n1912), .CLK(CLOCK), .RSTB(n5278), .Q(Datao[15]) );
  DFFARX1 \Datao_reg[16]  ( .D(n1911), .CLK(CLOCK), .RSTB(n5277), .Q(Datao[16]) );
  DFFARX1 \Datao_reg[17]  ( .D(n1910), .CLK(CLOCK), .RSTB(n5282), .Q(Datao[17]) );
  DFFARX1 \Datao_reg[18]  ( .D(n1909), .CLK(CLOCK), .RSTB(n5288), .Q(Datao[18]) );
  DFFARX1 \Datao_reg[19]  ( .D(n1908), .CLK(CLOCK), .RSTB(n5277), .Q(Datao[19]) );
  DFFARX1 \Datao_reg[20]  ( .D(n1907), .CLK(CLOCK), .RSTB(n5287), .Q(Datao[20]) );
  DFFARX1 \Datao_reg[21]  ( .D(n1906), .CLK(CLOCK), .RSTB(n5283), .Q(Datao[21]) );
  DFFARX1 \Datao_reg[22]  ( .D(n1905), .CLK(CLOCK), .RSTB(n5285), .Q(Datao[22]) );
  DFFARX1 \Datao_reg[23]  ( .D(n1904), .CLK(CLOCK), .RSTB(n5284), .Q(Datao[23]) );
  DFFARX1 \Datao_reg[24]  ( .D(n1903), .CLK(CLOCK), .RSTB(n5286), .Q(Datao[24]) );
  DFFARX1 \Datao_reg[25]  ( .D(n1902), .CLK(CLOCK), .RSTB(n5291), .Q(Datao[25]) );
  DFFARX1 \Datao_reg[26]  ( .D(n1901), .CLK(CLOCK), .RSTB(n5290), .Q(Datao[26]) );
  DFFARX1 \Datao_reg[27]  ( .D(n1900), .CLK(CLOCK), .RSTB(n5289), .Q(Datao[27]) );
  DFFARX1 \Datao_reg[28]  ( .D(n1899), .CLK(CLOCK), .RSTB(n5287), .Q(Datao[28]) );
  DFFARX1 \Datao_reg[29]  ( .D(n1898), .CLK(CLOCK), .RSTB(n5283), .Q(Datao[29]) );
  DFFARX1 \Datao_reg[30]  ( .D(n1897), .CLK(CLOCK), .RSTB(n5285), .Q(Datao[30]) );
  DFFARX1 \EBX_reg[0]  ( .D(n1888), .CLK(CLOCK), .RSTB(n5291), .Q(EBX[0]) );
  DFFARX1 \EBX_reg[1]  ( .D(n1887), .CLK(CLOCK), .RSTB(n5291), .Q(EBX[1]) );
  DFFARX1 \EBX_reg[2]  ( .D(n1886), .CLK(CLOCK), .RSTB(n5291), .Q(EBX[2]) );
  DFFARX1 \EBX_reg[3]  ( .D(n1885), .CLK(CLOCK), .RSTB(n5291), .Q(EBX[3]) );
  DFFARX1 \EBX_reg[4]  ( .D(n1884), .CLK(CLOCK), .RSTB(n5291), .Q(EBX[4]) );
  DFFARX1 \EBX_reg[5]  ( .D(n1883), .CLK(CLOCK), .RSTB(n5291), .Q(EBX[5]) );
  DFFARX1 \EBX_reg[6]  ( .D(n1882), .CLK(CLOCK), .RSTB(n5291), .Q(EBX[6]) );
  DFFARX1 \EBX_reg[7]  ( .D(n1881), .CLK(CLOCK), .RSTB(n5283), .Q(EBX[7]) );
  DFFARX1 \EBX_reg[8]  ( .D(n1880), .CLK(CLOCK), .RSTB(n5285), .Q(EBX[8]) );
  DFFARX1 \EBX_reg[9]  ( .D(n1879), .CLK(CLOCK), .RSTB(n5284), .Q(EBX[9]) );
  DFFARX1 \EBX_reg[10]  ( .D(n1878), .CLK(CLOCK), .RSTB(n5286), .Q(EBX[10]) );
  DFFARX1 \EBX_reg[11]  ( .D(n1877), .CLK(CLOCK), .RSTB(n5291), .Q(EBX[11]) );
  DFFARX1 \EBX_reg[12]  ( .D(n1876), .CLK(CLOCK), .RSTB(n5290), .Q(EBX[12]) );
  DFFARX1 \EBX_reg[13]  ( .D(n1875), .CLK(CLOCK), .RSTB(n5290), .Q(EBX[13]) );
  DFFARX1 \EBX_reg[14]  ( .D(n1874), .CLK(CLOCK), .RSTB(n5287), .Q(EBX[14]) );
  DFFARX1 \EBX_reg[15]  ( .D(n1873), .CLK(CLOCK), .RSTB(n5289), .Q(EBX[15]) );
  DFFARX1 \EBX_reg[16]  ( .D(n1872), .CLK(CLOCK), .RSTB(n5280), .Q(EBX[16]) );
  DFFARX1 \EBX_reg[17]  ( .D(n1871), .CLK(CLOCK), .RSTB(n5283), .Q(EBX[17]) );
  DFFARX1 \EBX_reg[18]  ( .D(n1870), .CLK(CLOCK), .RSTB(n5278), .Q(EBX[18]) );
  DFFARX1 \EBX_reg[19]  ( .D(n1869), .CLK(CLOCK), .RSTB(n5283), .Q(EBX[19]) );
  DFFARX1 \EBX_reg[20]  ( .D(n1868), .CLK(CLOCK), .RSTB(n5285), .Q(EBX[20]) );
  DFFARX1 \EBX_reg[21]  ( .D(n1867), .CLK(CLOCK), .RSTB(n5284), .Q(EBX[21]) );
  DFFARX1 \EBX_reg[22]  ( .D(n1866), .CLK(CLOCK), .RSTB(n5286), .Q(EBX[22]) );
  DFFARX1 \EBX_reg[23]  ( .D(n1865), .CLK(CLOCK), .RSTB(n5291), .Q(EBX[23]) );
  DFFARX1 \EBX_reg[24]  ( .D(n1864), .CLK(CLOCK), .RSTB(n5290), .Q(EBX[24]) );
  DFFARX1 \EBX_reg[25]  ( .D(n1863), .CLK(CLOCK), .RSTB(n5289), .Q(EBX[25]) );
  DFFARX1 \EBX_reg[26]  ( .D(n1862), .CLK(CLOCK), .RSTB(n5289), .Q(EBX[26]) );
  DFFARX1 \EBX_reg[27]  ( .D(n1861), .CLK(CLOCK), .RSTB(n5287), .Q(EBX[27]) );
  DFFARX1 \EBX_reg[28]  ( .D(n1860), .CLK(CLOCK), .RSTB(n5285), .Q(EBX[28]) );
  DFFARX1 \EBX_reg[29]  ( .D(n1859), .CLK(CLOCK), .RSTB(n5282), .Q(EBX[29]) );
  DFFARX1 \EBX_reg[30]  ( .D(n1858), .CLK(CLOCK), .RSTB(n5281), .Q(EBX[30]) );
  DFFARX1 \EBX_reg[31]  ( .D(n1857), .CLK(CLOCK), .RSTB(n5291), .Q(N1989) );
  DFFARX1 \PhyAddrPointer_reg[0]  ( .D(n1736), .CLK(CLOCK), .RSTB(n5288), .Q(
        N1009), .QN(n5196) );
  DFFARX1 \rEIP_reg[0]  ( .D(n2065), .CLK(CLOCK), .RSTB(n5291), .Q(rEIP[0]) );
  DFFARX1 \InstAddrPointer_reg[0]  ( .D(n2021), .CLK(CLOCK), .RSTB(n5289), .Q(
        N1868), .QN(n5204) );
  DFFARX1 \InstQueueRd_Addr_reg[0]  ( .D(n2028), .CLK(CLOCK), .RSTB(n5286), 
        .Q(N2884), .QN(n5183) );
  DFFARX1 \PhyAddrPointer_reg[1]  ( .D(n1735), .CLK(CLOCK), .RSTB(n5281), .Q(
        PhyAddrPointer[1]), .QN(n5201) );
  DFFARX1 \rEIP_reg[1]  ( .D(n2064), .CLK(CLOCK), .RSTB(n5289), .Q(N4154), 
        .QN(n5190) );
  DFFARX1 \InstAddrPointer_reg[1]  ( .D(n2020), .CLK(CLOCK), .RSTB(n5280), .Q(
        InstAddrPointer[1]), .QN(n5185) );
  DFFARX1 \InstQueueRd_Addr_reg[1]  ( .D(n2027), .CLK(CLOCK), .RSTB(n5281), 
        .Q(InstQueueRd_Addr[1]), .QN(n5177) );
  DFFARX1 \InstQueueRd_Addr_reg[2]  ( .D(n2026), .CLK(CLOCK), .RSTB(n5288), 
        .Q(InstQueueRd_Addr[2]), .QN(n5180) );
  DFFARX1 \InstQueueRd_Addr_reg[3]  ( .D(n2025), .CLK(CLOCK), .RSTB(n5290), 
        .Q(InstQueueRd_Addr[3]), .QN(n5206) );
  DFFARX1 \PhyAddrPointer_reg[2]  ( .D(n1734), .CLK(CLOCK), .RSTB(n5285), .Q(
        PhyAddrPointer[2]), .QN(n5214) );
  DFFARX1 \rEIP_reg[2]  ( .D(n2063), .CLK(CLOCK), .RSTB(n5284), .Q(rEIP[2]) );
  DFFARX1 \InstAddrPointer_reg[2]  ( .D(n2019), .CLK(CLOCK), .RSTB(n5280), .Q(
        InstAddrPointer[2]) );
  DFFARX1 \PhyAddrPointer_reg[3]  ( .D(n1733), .CLK(CLOCK), .RSTB(n5283), .Q(
        PhyAddrPointer[3]), .QN(n5253) );
  DFFARX1 \rEIP_reg[3]  ( .D(n2062), .CLK(CLOCK), .RSTB(n5287), .Q(rEIP[3]), 
        .QN(n5217) );
  DFFARX1 \InstAddrPointer_reg[3]  ( .D(n2018), .CLK(CLOCK), .RSTB(n5281), .Q(
        InstAddrPointer[3]), .QN(n5222) );
  DFFARX1 \PhyAddrPointer_reg[4]  ( .D(n1732), .CLK(CLOCK), .RSTB(n5291), .Q(
        PhyAddrPointer[4]) );
  DFFARX1 \rEIP_reg[4]  ( .D(n2061), .CLK(CLOCK), .RSTB(n5290), .Q(rEIP[4]) );
  DFFARX1 \InstAddrPointer_reg[4]  ( .D(n2017), .CLK(CLOCK), .RSTB(n5277), .Q(
        InstAddrPointer[4]) );
  DFFARX1 \PhyAddrPointer_reg[5]  ( .D(n1731), .CLK(CLOCK), .RSTB(n5284), .Q(
        PhyAddrPointer[5]), .QN(n5181) );
  DFFARX1 \rEIP_reg[5]  ( .D(n2060), .CLK(CLOCK), .RSTB(n5286), .Q(rEIP[5]), 
        .QN(n5260) );
  DFFARX1 \InstAddrPointer_reg[5]  ( .D(n2016), .CLK(CLOCK), .RSTB(n5282), .Q(
        InstAddrPointer[5]), .QN(n5205) );
  DFFARX1 \PhyAddrPointer_reg[6]  ( .D(n1730), .CLK(CLOCK), .RSTB(n5283), .Q(
        PhyAddrPointer[6]), .QN(n5184) );
  DFFARX1 \rEIP_reg[6]  ( .D(n2059), .CLK(CLOCK), .RSTB(n5285), .Q(rEIP[6]), 
        .QN(n5261) );
  DFFARX1 \InstAddrPointer_reg[6]  ( .D(n2015), .CLK(CLOCK), .RSTB(n5278), .Q(
        InstAddrPointer[6]) );
  DFFARX1 \PhyAddrPointer_reg[7]  ( .D(n1729), .CLK(CLOCK), .RSTB(n5287), .Q(
        PhyAddrPointer[7]) );
  DFFARX1 \rEIP_reg[7]  ( .D(n2058), .CLK(CLOCK), .RSTB(n5279), .Q(rEIP[7]) );
  DFFARX1 \InstAddrPointer_reg[7]  ( .D(n2014), .CLK(CLOCK), .RSTB(n5288), .Q(
        InstAddrPointer[7]), .QN(n5209) );
  DFFARX1 \PhyAddrPointer_reg[8]  ( .D(n1728), .CLK(CLOCK), .RSTB(n5290), .Q(
        PhyAddrPointer[8]), .QN(n5189) );
  DFFARX1 \rEIP_reg[8]  ( .D(n2057), .CLK(CLOCK), .RSTB(n5291), .Q(rEIP[8]), 
        .QN(n5259) );
  DFFARX1 \InstAddrPointer_reg[8]  ( .D(n2013), .CLK(CLOCK), .RSTB(n5286), .Q(
        InstAddrPointer[8]), .QN(n5225) );
  DFFARX1 \PhyAddrPointer_reg[9]  ( .D(n1727), .CLK(CLOCK), .RSTB(n5279), .Q(
        PhyAddrPointer[9]) );
  DFFARX1 \rEIP_reg[9]  ( .D(n2056), .CLK(CLOCK), .RSTB(n5289), .Q(rEIP[9]) );
  DFFARX1 \InstAddrPointer_reg[9]  ( .D(n2012), .CLK(CLOCK), .RSTB(n5281), .Q(
        InstAddrPointer[9]), .QN(n5218) );
  DFFARX1 \PhyAddrPointer_reg[10]  ( .D(n1726), .CLK(CLOCK), .RSTB(n5288), .Q(
        PhyAddrPointer[10]), .QN(n5195) );
  DFFARX1 \rEIP_reg[10]  ( .D(n2055), .CLK(CLOCK), .RSTB(n5284), .Q(rEIP[10]), 
        .QN(n5258) );
  DFFARX1 \InstAddrPointer_reg[10]  ( .D(n2011), .CLK(CLOCK), .RSTB(n5289), 
        .Q(InstAddrPointer[10]), .QN(n5229) );
  DFFARX1 \PhyAddrPointer_reg[11]  ( .D(n1725), .CLK(CLOCK), .RSTB(n5277), .Q(
        PhyAddrPointer[11]) );
  DFFARX1 \rEIP_reg[11]  ( .D(n2054), .CLK(CLOCK), .RSTB(n5278), .Q(rEIP[11])
         );
  DFFARX1 \InstAddrPointer_reg[11]  ( .D(n2010), .CLK(CLOCK), .RSTB(n5291), 
        .Q(InstAddrPointer[11]), .QN(n5219) );
  DFFARX1 \PhyAddrPointer_reg[12]  ( .D(n1724), .CLK(CLOCK), .RSTB(n5279), .Q(
        PhyAddrPointer[12]), .QN(n5194) );
  DFFARX1 \rEIP_reg[12]  ( .D(n2053), .CLK(CLOCK), .RSTB(n5280), .Q(rEIP[12]), 
        .QN(n5257) );
  DFFARX1 \InstAddrPointer_reg[12]  ( .D(n2009), .CLK(CLOCK), .RSTB(n5281), 
        .Q(InstAddrPointer[12]), .QN(n5228) );
  DFFARX1 \PhyAddrPointer_reg[13]  ( .D(n1723), .CLK(CLOCK), .RSTB(n5282), .Q(
        PhyAddrPointer[13]) );
  DFFARX1 \rEIP_reg[13]  ( .D(n2052), .CLK(CLOCK), .RSTB(n5288), .Q(rEIP[13])
         );
  DFFARX1 \InstAddrPointer_reg[13]  ( .D(n2008), .CLK(CLOCK), .RSTB(n5282), 
        .Q(InstAddrPointer[13]), .QN(n5220) );
  DFFARX1 \PhyAddrPointer_reg[14]  ( .D(n1722), .CLK(CLOCK), .RSTB(n5283), .Q(
        PhyAddrPointer[14]), .QN(n5193) );
  DFFARX1 \rEIP_reg[14]  ( .D(n2051), .CLK(CLOCK), .RSTB(n5287), .Q(rEIP[14]), 
        .QN(n5256) );
  DFFARX1 \InstAddrPointer_reg[14]  ( .D(n2007), .CLK(CLOCK), .RSTB(n5288), 
        .Q(InstAddrPointer[14]), .QN(n5227) );
  DFFARX1 \PhyAddrPointer_reg[15]  ( .D(n1721), .CLK(CLOCK), .RSTB(n5286), .Q(
        PhyAddrPointer[15]) );
  DFFARX1 \rEIP_reg[15]  ( .D(n2050), .CLK(CLOCK), .RSTB(n5291), .Q(rEIP[15])
         );
  DFFARX1 \InstAddrPointer_reg[15]  ( .D(n2006), .CLK(CLOCK), .RSTB(n5287), 
        .Q(InstAddrPointer[15]), .QN(n5221) );
  DFFARX1 \PhyAddrPointer_reg[16]  ( .D(n1720), .CLK(CLOCK), .RSTB(n5284), .Q(
        PhyAddrPointer[16]), .QN(n5192) );
  DFFARX1 \rEIP_reg[16]  ( .D(n2049), .CLK(CLOCK), .RSTB(n5285), .Q(rEIP[16]), 
        .QN(n5255) );
  DFFARX1 \InstAddrPointer_reg[16]  ( .D(n2005), .CLK(CLOCK), .RSTB(n5283), 
        .Q(InstAddrPointer[16]), .QN(n5226) );
  DFFARX1 \PhyAddrPointer_reg[17]  ( .D(n1719), .CLK(CLOCK), .RSTB(n5285), .Q(
        PhyAddrPointer[17]), .QN(n5241) );
  DFFARX1 \rEIP_reg[17]  ( .D(n2048), .CLK(CLOCK), .RSTB(n5284), .Q(rEIP[17])
         );
  DFFARX1 \InstAddrPointer_reg[17]  ( .D(n2004), .CLK(CLOCK), .RSTB(n5290), 
        .Q(InstAddrPointer[17]), .QN(n5234) );
  DFFARX1 \PhyAddrPointer_reg[18]  ( .D(n1718), .CLK(CLOCK), .RSTB(n5281), .Q(
        PhyAddrPointer[18]), .QN(n5191) );
  DFFARX1 \rEIP_reg[18]  ( .D(n2047), .CLK(CLOCK), .RSTB(n5289), .Q(rEIP[18]), 
        .QN(n5254) );
  DFFARX1 \InstAddrPointer_reg[18]  ( .D(n2003), .CLK(CLOCK), .RSTB(n5278), 
        .Q(InstAddrPointer[18]), .QN(n5238) );
  DFFARX1 \PhyAddrPointer_reg[19]  ( .D(n1717), .CLK(CLOCK), .RSTB(n5289), .Q(
        PhyAddrPointer[19]) );
  DFFARX1 \rEIP_reg[19]  ( .D(n2046), .CLK(CLOCK), .RSTB(n5289), .Q(rEIP[19])
         );
  DFFARX1 \InstAddrPointer_reg[19]  ( .D(n2002), .CLK(CLOCK), .RSTB(n5286), 
        .Q(InstAddrPointer[19]), .QN(n5235) );
  DFFARX1 \PhyAddrPointer_reg[20]  ( .D(n1716), .CLK(CLOCK), .RSTB(n5289), .Q(
        PhyAddrPointer[20]), .QN(n5247) );
  DFFARX1 \rEIP_reg[20]  ( .D(n2045), .CLK(CLOCK), .RSTB(n5289), .Q(rEIP[20])
         );
  DFFARX1 \InstAddrPointer_reg[20]  ( .D(n2001), .CLK(CLOCK), .RSTB(n5282), 
        .Q(InstAddrPointer[20]), .QN(n5215) );
  DFFARX1 \PhyAddrPointer_reg[21]  ( .D(n1715), .CLK(CLOCK), .RSTB(n5289), .Q(
        PhyAddrPointer[21]) );
  DFFARX1 \rEIP_reg[21]  ( .D(n2044), .CLK(CLOCK), .RSTB(n5289), .Q(rEIP[21]), 
        .QN(n5188) );
  DFFARX1 \InstAddrPointer_reg[21]  ( .D(n2000), .CLK(CLOCK), .RSTB(n5278), 
        .Q(InstAddrPointer[21]), .QN(n5210) );
  DFFARX1 \PhyAddrPointer_reg[22]  ( .D(n1714), .CLK(CLOCK), .RSTB(n5289), .Q(
        PhyAddrPointer[22]), .QN(n5246) );
  DFFARX1 \rEIP_reg[22]  ( .D(n2043), .CLK(CLOCK), .RSTB(n5289), .Q(rEIP[22])
         );
  DFFARX1 \InstAddrPointer_reg[22]  ( .D(n1999), .CLK(CLOCK), .RSTB(n5277), 
        .Q(InstAddrPointer[22]), .QN(n5231) );
  DFFARX1 \PhyAddrPointer_reg[23]  ( .D(n1713), .CLK(CLOCK), .RSTB(n5289), .Q(
        PhyAddrPointer[23]) );
  DFFARX1 \rEIP_reg[23]  ( .D(n2042), .CLK(CLOCK), .RSTB(n5289), .Q(rEIP[23]), 
        .QN(n5216) );
  DFFARX1 \InstAddrPointer_reg[23]  ( .D(n1998), .CLK(CLOCK), .RSTB(n5279), 
        .Q(InstAddrPointer[23]), .QN(n5211) );
  DFFARX1 \PhyAddrPointer_reg[24]  ( .D(n1712), .CLK(CLOCK), .RSTB(n5289), .Q(
        PhyAddrPointer[24]), .QN(n5245) );
  DFFARX1 \rEIP_reg[24]  ( .D(n2041), .CLK(CLOCK), .RSTB(n5289), .Q(rEIP[24])
         );
  DFFARX1 \InstAddrPointer_reg[24]  ( .D(n1997), .CLK(CLOCK), .RSTB(n5280), 
        .Q(InstAddrPointer[24]), .QN(n5232) );
  DFFARX1 \PhyAddrPointer_reg[25]  ( .D(n1711), .CLK(CLOCK), .RSTB(n5290), .Q(
        PhyAddrPointer[25]) );
  DFFARX1 \rEIP_reg[25]  ( .D(n2040), .CLK(CLOCK), .RSTB(n5290), .Q(rEIP[25]), 
        .QN(n5187) );
  DFFARX1 \InstAddrPointer_reg[25]  ( .D(n1996), .CLK(CLOCK), .RSTB(n5281), 
        .Q(InstAddrPointer[25]), .QN(n5212) );
  DFFARX1 \PhyAddrPointer_reg[26]  ( .D(n1710), .CLK(CLOCK), .RSTB(n5290), .Q(
        PhyAddrPointer[26]), .QN(n5244) );
  DFFARX1 \rEIP_reg[26]  ( .D(n2039), .CLK(CLOCK), .RSTB(n5290), .Q(rEIP[26])
         );
  DFFARX1 \InstAddrPointer_reg[26]  ( .D(n1995), .CLK(CLOCK), .RSTB(n5289), 
        .Q(InstAddrPointer[26]), .QN(n5233) );
  DFFARX1 \PhyAddrPointer_reg[27]  ( .D(n1709), .CLK(CLOCK), .RSTB(n5290), .Q(
        PhyAddrPointer[27]) );
  DFFARX1 \rEIP_reg[27]  ( .D(n2038), .CLK(CLOCK), .RSTB(n5290), .Q(rEIP[27]), 
        .QN(n5186) );
  DFFARX1 \InstAddrPointer_reg[27]  ( .D(n1994), .CLK(CLOCK), .RSTB(n5290), 
        .Q(InstAddrPointer[27]), .QN(n5213) );
  DFFARX1 \PhyAddrPointer_reg[28]  ( .D(n1708), .CLK(CLOCK), .RSTB(n5290), .Q(
        PhyAddrPointer[28]), .QN(n5243) );
  DFFARX1 \rEIP_reg[28]  ( .D(n2037), .CLK(CLOCK), .RSTB(n5290), .Q(rEIP[28])
         );
  DFFARX1 \InstAddrPointer_reg[28]  ( .D(n1993), .CLK(CLOCK), .RSTB(n5291), 
        .Q(InstAddrPointer[28]), .QN(n5237) );
  DFFARX1 \PhyAddrPointer_reg[29]  ( .D(n1707), .CLK(CLOCK), .RSTB(n5290), .Q(
        PhyAddrPointer[29]), .QN(n5240) );
  DFFARX1 \rEIP_reg[29]  ( .D(n2036), .CLK(CLOCK), .RSTB(n5290), .Q(rEIP[29])
         );
  DFFARX1 \InstAddrPointer_reg[29]  ( .D(n1992), .CLK(CLOCK), .RSTB(n5290), 
        .Q(InstAddrPointer[29]), .QN(n5223) );
  DFFARX1 \PhyAddrPointer_reg[30]  ( .D(n1706), .CLK(CLOCK), .RSTB(n5291), .Q(
        PhyAddrPointer[30]) );
  DFFARX1 \rEIP_reg[30]  ( .D(n2035), .CLK(CLOCK), .RSTB(n5291), .Q(rEIP[30])
         );
  DFFARX1 \InstAddrPointer_reg[30]  ( .D(n1991), .CLK(CLOCK), .RSTB(n5291), 
        .Q(InstAddrPointer[30]), .QN(n5230) );
  DFFARX1 \PhyAddrPointer_reg[31]  ( .D(n1705), .CLK(CLOCK), .RSTB(n5281), .Q(
        PhyAddrPointer[31]), .QN(n5239) );
  DFFARX1 \rEIP_reg[31]  ( .D(n2071), .CLK(CLOCK), .RSTB(n5291), .Q(rEIP[31]), 
        .QN(n5248) );
  DFFARX1 \InstAddrPointer_reg[31]  ( .D(n2070), .CLK(CLOCK), .RSTB(n5290), 
        .Q(N3678), .QN(n5224) );
  DFFARX1 \InstQueueWr_Addr_reg[1]  ( .D(n2023), .CLK(CLOCK), .RSTB(n5284), 
        .Q(N4188), .QN(n5182) );
  DFFARX1 \InstQueueWr_Addr_reg[2]  ( .D(n2022), .CLK(CLOCK), .RSTB(n5286), 
        .Q(N4187), .QN(n5198) );
  DFFARX1 \InstQueueWr_Addr_reg[3]  ( .D(n2033), .CLK(CLOCK), .RSTB(n5291), 
        .Q(N4186), .QN(n5200) );
  DFFARX1 \InstQueue_reg[3][0]  ( .D(n1840), .CLK(CLOCK), .RSTB(n5290), .Q(
        \InstQueue[3][0] ) );
  DFFARX1 \InstQueue_reg[3][1]  ( .D(n1839), .CLK(CLOCK), .RSTB(n5291), .Q(
        \InstQueue[3][1] ) );
  DFFARX1 \InstQueue_reg[3][2]  ( .D(n1838), .CLK(CLOCK), .RSTB(n5288), .Q(
        \InstQueue[3][2] ) );
  DFFARX1 \InstQueue_reg[3][3]  ( .D(n1837), .CLK(CLOCK), .RSTB(n5290), .Q(
        \InstQueue[3][3] ) );
  DFFARX1 \InstQueue_reg[3][4]  ( .D(n1836), .CLK(CLOCK), .RSTB(n5289), .Q(
        \InstQueue[3][4] ) );
  DFFARX1 \InstQueue_reg[3][5]  ( .D(n1835), .CLK(CLOCK), .RSTB(n5278), .Q(
        \InstQueue[3][5] ) );
  DFFARX1 \InstQueue_reg[3][6]  ( .D(n1834), .CLK(CLOCK), .RSTB(n5278), .Q(
        \InstQueue[3][6] ) );
  DFFARX1 \InstQueue_reg[3][7]  ( .D(n1833), .CLK(CLOCK), .RSTB(n5278), .Q(
        \InstQueue[3][7] ) );
  DFFARX1 \InstQueue_reg[4][0]  ( .D(n1832), .CLK(CLOCK), .RSTB(n5278), .Q(
        \InstQueue[4][0] ) );
  DFFARX1 \InstQueue_reg[4][1]  ( .D(n1831), .CLK(CLOCK), .RSTB(n5278), .Q(
        \InstQueue[4][1] ) );
  DFFARX1 \InstQueue_reg[4][2]  ( .D(n1830), .CLK(CLOCK), .RSTB(n5278), .Q(
        \InstQueue[4][2] ) );
  DFFARX1 \InstQueue_reg[4][3]  ( .D(n1829), .CLK(CLOCK), .RSTB(n5278), .Q(
        \InstQueue[4][3] ) );
  DFFARX1 \InstQueue_reg[4][4]  ( .D(n1828), .CLK(CLOCK), .RSTB(n5278), .Q(
        \InstQueue[4][4] ) );
  DFFARX1 \InstQueue_reg[4][5]  ( .D(n1827), .CLK(CLOCK), .RSTB(n5278), .Q(
        \InstQueue[4][5] ) );
  DFFARX1 \InstQueue_reg[4][6]  ( .D(n1826), .CLK(CLOCK), .RSTB(n5278), .Q(
        \InstQueue[4][6] ) );
  DFFARX1 \InstQueue_reg[4][7]  ( .D(n1825), .CLK(CLOCK), .RSTB(n5278), .Q(
        \InstQueue[4][7] ) );
  DFFARX1 \InstQueue_reg[5][0]  ( .D(n1824), .CLK(CLOCK), .RSTB(n5278), .Q(
        \InstQueue[5][0] ), .QN(n5276) );
  DFFARX1 \InstQueue_reg[5][1]  ( .D(n1823), .CLK(CLOCK), .RSTB(n5279), .Q(
        \InstQueue[5][1] ), .QN(n5275) );
  DFFARX1 \InstQueue_reg[5][2]  ( .D(n1822), .CLK(CLOCK), .RSTB(n5279), .Q(
        \InstQueue[5][2] ), .QN(n5274) );
  DFFARX1 \InstQueue_reg[5][3]  ( .D(n1821), .CLK(CLOCK), .RSTB(n5279), .Q(
        \InstQueue[5][3] ), .QN(n5270) );
  DFFARX1 \InstQueue_reg[5][4]  ( .D(n1820), .CLK(CLOCK), .RSTB(n5279), .Q(
        \InstQueue[5][4] ), .QN(n5273) );
  DFFARX1 \InstQueue_reg[5][5]  ( .D(n1819), .CLK(CLOCK), .RSTB(n5279), .Q(
        \InstQueue[5][5] ), .QN(n5272) );
  DFFARX1 \InstQueue_reg[5][6]  ( .D(n1818), .CLK(CLOCK), .RSTB(n5279), .Q(
        \InstQueue[5][6] ), .QN(n5271) );
  DFFARX1 \InstQueue_reg[5][7]  ( .D(n1817), .CLK(CLOCK), .RSTB(n5279), .Q(
        \InstQueue[5][7] ) );
  DFFARX1 \InstQueue_reg[6][0]  ( .D(n1816), .CLK(CLOCK), .RSTB(n5279), .Q(
        \InstQueue[6][0] ) );
  DFFARX1 \InstQueue_reg[6][1]  ( .D(n1815), .CLK(CLOCK), .RSTB(n5279), .Q(
        \InstQueue[6][1] ) );
  DFFARX1 \InstQueue_reg[6][2]  ( .D(n1814), .CLK(CLOCK), .RSTB(n5279), .Q(
        \InstQueue[6][2] ) );
  DFFARX1 \InstQueue_reg[6][3]  ( .D(n1813), .CLK(CLOCK), .RSTB(n5279), .Q(
        \InstQueue[6][3] ) );
  DFFARX1 \InstQueue_reg[6][4]  ( .D(n1812), .CLK(CLOCK), .RSTB(n5279), .Q(
        \InstQueue[6][4] ) );
  DFFARX1 \InstQueue_reg[6][5]  ( .D(n1811), .CLK(CLOCK), .RSTB(n5280), .Q(
        \InstQueue[6][5] ) );
  DFFARX1 \InstQueue_reg[6][6]  ( .D(n1810), .CLK(CLOCK), .RSTB(n5280), .Q(
        \InstQueue[6][6] ) );
  DFFARX1 \InstQueue_reg[6][7]  ( .D(n1809), .CLK(CLOCK), .RSTB(n5280), .Q(
        \InstQueue[6][7] ) );
  DFFARX1 \InstQueue_reg[7][0]  ( .D(n1808), .CLK(CLOCK), .RSTB(n5280), .Q(
        \InstQueue[7][0] ) );
  DFFARX1 \InstQueue_reg[7][1]  ( .D(n1807), .CLK(CLOCK), .RSTB(n5280), .Q(
        \InstQueue[7][1] ) );
  DFFARX1 \InstQueue_reg[7][2]  ( .D(n1806), .CLK(CLOCK), .RSTB(n5280), .Q(
        \InstQueue[7][2] ) );
  DFFARX1 \InstQueue_reg[7][3]  ( .D(n1805), .CLK(CLOCK), .RSTB(n5280), .Q(
        \InstQueue[7][3] ) );
  DFFARX1 \InstQueue_reg[7][4]  ( .D(n1804), .CLK(CLOCK), .RSTB(n5280), .Q(
        \InstQueue[7][4] ) );
  DFFARX1 \InstQueue_reg[7][5]  ( .D(n1803), .CLK(CLOCK), .RSTB(n5280), .Q(
        \InstQueue[7][5] ) );
  DFFARX1 \InstQueue_reg[7][6]  ( .D(n1802), .CLK(CLOCK), .RSTB(n5280), .Q(
        \InstQueue[7][6] ) );
  DFFARX1 \InstQueue_reg[7][7]  ( .D(n1801), .CLK(CLOCK), .RSTB(n5280), .Q(
        \InstQueue[7][7] ) );
  DFFARX1 \InstQueue_reg[8][0]  ( .D(n1800), .CLK(CLOCK), .RSTB(n5280), .Q(
        \InstQueue[8][0] ) );
  DFFARX1 \InstQueue_reg[8][1]  ( .D(n1799), .CLK(CLOCK), .RSTB(n5281), .Q(
        \InstQueue[8][1] ) );
  DFFARX1 \InstQueue_reg[8][2]  ( .D(n1798), .CLK(CLOCK), .RSTB(n5281), .Q(
        \InstQueue[8][2] ) );
  DFFARX1 \InstQueue_reg[8][3]  ( .D(n1797), .CLK(CLOCK), .RSTB(n5281), .Q(
        \InstQueue[8][3] ) );
  DFFARX1 \InstQueue_reg[8][4]  ( .D(n1796), .CLK(CLOCK), .RSTB(n5281), .Q(
        \InstQueue[8][4] ) );
  DFFARX1 \InstQueue_reg[8][5]  ( .D(n1795), .CLK(CLOCK), .RSTB(n5281), .Q(
        \InstQueue[8][5] ) );
  DFFARX1 \InstQueue_reg[8][6]  ( .D(n1794), .CLK(CLOCK), .RSTB(n5281), .Q(
        \InstQueue[8][6] ) );
  DFFARX1 \InstQueue_reg[8][7]  ( .D(n1793), .CLK(CLOCK), .RSTB(n5281), .Q(
        \InstQueue[8][7] ) );
  DFFARX1 \InstQueue_reg[9][0]  ( .D(n1792), .CLK(CLOCK), .RSTB(n5281), .Q(
        \InstQueue[9][0] ), .QN(n5269) );
  DFFARX1 \InstQueue_reg[9][1]  ( .D(n1791), .CLK(CLOCK), .RSTB(n5281), .Q(
        \InstQueue[9][1] ), .QN(n5268) );
  DFFARX1 \InstQueue_reg[9][2]  ( .D(n1790), .CLK(CLOCK), .RSTB(n5281), .Q(
        \InstQueue[9][2] ), .QN(n5267) );
  DFFARX1 \InstQueue_reg[9][3]  ( .D(n1789), .CLK(CLOCK), .RSTB(n5281), .Q(
        \InstQueue[9][3] ), .QN(n5263) );
  DFFARX1 \InstQueue_reg[9][4]  ( .D(n1788), .CLK(CLOCK), .RSTB(n5281), .Q(
        \InstQueue[9][4] ), .QN(n5266) );
  DFFARX1 \InstQueue_reg[9][5]  ( .D(n1787), .CLK(CLOCK), .RSTB(n5282), .Q(
        \InstQueue[9][5] ), .QN(n5265) );
  DFFARX1 \InstQueue_reg[9][6]  ( .D(n1786), .CLK(CLOCK), .RSTB(n5282), .Q(
        \InstQueue[9][6] ), .QN(n5264) );
  DFFARX1 \InstQueue_reg[9][7]  ( .D(n1785), .CLK(CLOCK), .RSTB(n5282), .Q(
        \InstQueue[9][7] ) );
  DFFARX1 \InstQueue_reg[10][0]  ( .D(n1784), .CLK(CLOCK), .RSTB(n5282), .Q(
        \InstQueue[10][0] ) );
  DFFARX1 \InstQueue_reg[10][1]  ( .D(n1783), .CLK(CLOCK), .RSTB(n5282), .Q(
        \InstQueue[10][1] ) );
  DFFARX1 \InstQueue_reg[10][2]  ( .D(n1782), .CLK(CLOCK), .RSTB(n5282), .Q(
        \InstQueue[10][2] ) );
  DFFARX1 \InstQueue_reg[10][3]  ( .D(n1781), .CLK(CLOCK), .RSTB(n5282), .Q(
        \InstQueue[10][3] ) );
  DFFARX1 \InstQueue_reg[10][4]  ( .D(n1780), .CLK(CLOCK), .RSTB(n5282), .Q(
        \InstQueue[10][4] ) );
  DFFARX1 \InstQueue_reg[10][5]  ( .D(n1779), .CLK(CLOCK), .RSTB(n5282), .Q(
        \InstQueue[10][5] ) );
  DFFARX1 \InstQueue_reg[10][6]  ( .D(n1778), .CLK(CLOCK), .RSTB(n5282), .Q(
        \InstQueue[10][6] ) );
  DFFARX1 \InstQueue_reg[10][7]  ( .D(n1777), .CLK(CLOCK), .RSTB(n5282), .Q(
        \InstQueue[10][7] ) );
  DFFARX1 \InstQueue_reg[11][0]  ( .D(n1776), .CLK(CLOCK), .RSTB(n5282), .Q(
        \InstQueue[11][0] ) );
  DFFARX1 \InstQueue_reg[11][1]  ( .D(n1775), .CLK(CLOCK), .RSTB(n5283), .Q(
        \InstQueue[11][1] ) );
  DFFARX1 \InstQueue_reg[11][2]  ( .D(n1774), .CLK(CLOCK), .RSTB(n5283), .Q(
        \InstQueue[11][2] ) );
  DFFARX1 \InstQueue_reg[11][3]  ( .D(n1773), .CLK(CLOCK), .RSTB(n5283), .Q(
        \InstQueue[11][3] ) );
  DFFARX1 \InstQueue_reg[11][4]  ( .D(n1772), .CLK(CLOCK), .RSTB(n5283), .Q(
        \InstQueue[11][4] ) );
  DFFARX1 \InstQueue_reg[11][5]  ( .D(n1771), .CLK(CLOCK), .RSTB(n5283), .Q(
        \InstQueue[11][5] ) );
  DFFARX1 \InstQueue_reg[11][6]  ( .D(n1770), .CLK(CLOCK), .RSTB(n5283), .Q(
        \InstQueue[11][6] ) );
  DFFARX1 \InstQueue_reg[11][7]  ( .D(n1769), .CLK(CLOCK), .RSTB(n5283), .Q(
        \InstQueue[11][7] ) );
  DFFARX1 \InstQueue_reg[2][0]  ( .D(n1848), .CLK(CLOCK), .RSTB(n5283), .Q(
        \InstQueue[2][0] ) );
  DFFARX1 \InstQueue_reg[2][1]  ( .D(n1847), .CLK(CLOCK), .RSTB(n5283), .Q(
        \InstQueue[2][1] ) );
  DFFARX1 \InstQueue_reg[2][2]  ( .D(n1846), .CLK(CLOCK), .RSTB(n5283), .Q(
        \InstQueue[2][2] ) );
  DFFARX1 \InstQueue_reg[2][3]  ( .D(n1845), .CLK(CLOCK), .RSTB(n5283), .Q(
        \InstQueue[2][3] ) );
  DFFARX1 \InstQueue_reg[2][4]  ( .D(n1844), .CLK(CLOCK), .RSTB(n5283), .Q(
        \InstQueue[2][4] ) );
  DFFARX1 \InstQueue_reg[2][5]  ( .D(n1843), .CLK(CLOCK), .RSTB(n5284), .Q(
        \InstQueue[2][5] ) );
  DFFARX1 \InstQueue_reg[2][6]  ( .D(n1842), .CLK(CLOCK), .RSTB(n5284), .Q(
        \InstQueue[2][6] ) );
  DFFARX1 \InstQueue_reg[2][7]  ( .D(n1841), .CLK(CLOCK), .RSTB(n5284), .Q(
        \InstQueue[2][7] ) );
  DFFARX1 \InstQueue_reg[0][0]  ( .D(n1896), .CLK(CLOCK), .RSTB(n5280), .Q(
        \DP_OP_469J1_133_8416/n116 ) );
  DFFARX1 \InstQueue_reg[0][1]  ( .D(n1895), .CLK(CLOCK), .RSTB(n5283), .Q(
        \DP_OP_469J1_133_8416/n117 ) );
  DFFARX1 \InstQueue_reg[0][2]  ( .D(n1894), .CLK(CLOCK), .RSTB(n5279), .Q(
        \DP_OP_469J1_133_8416/n118 ) );
  DFFARX1 \InstQueue_reg[0][3]  ( .D(n1893), .CLK(CLOCK), .RSTB(n5277), .Q(
        \DP_OP_469J1_133_8416/n119 ) );
  DFFARX1 \InstQueue_reg[0][4]  ( .D(n1892), .CLK(CLOCK), .RSTB(n5278), .Q(
        \DP_OP_469J1_133_8416/n120 ) );
  DFFARX1 \InstQueue_reg[0][5]  ( .D(n1891), .CLK(CLOCK), .RSTB(n5286), .Q(
        \DP_OP_469J1_133_8416/n121 ) );
  DFFARX1 \InstQueue_reg[0][6]  ( .D(n1890), .CLK(CLOCK), .RSTB(n5288), .Q(
        \DP_OP_469J1_133_8416/n122 ) );
  DFFARX1 \InstQueue_reg[0][7]  ( .D(n1889), .CLK(CLOCK), .RSTB(n5280), .Q(
        \DP_OP_469J1_133_8416/n123 ) );
  DFFARX1 \InstQueue_reg[1][0]  ( .D(n1856), .CLK(CLOCK), .RSTB(n5284), .Q(
        \InstQueue[1][0] ) );
  DFFARX1 \InstQueue_reg[1][1]  ( .D(n1855), .CLK(CLOCK), .RSTB(n5284), .Q(
        \InstQueue[1][1] ) );
  DFFARX1 \InstQueue_reg[1][2]  ( .D(n1854), .CLK(CLOCK), .RSTB(n5284), .Q(
        \InstQueue[1][2] ) );
  DFFARX1 \InstQueue_reg[1][3]  ( .D(n1853), .CLK(CLOCK), .RSTB(n5284), .Q(
        \InstQueue[1][3] ) );
  DFFARX1 \InstQueue_reg[1][4]  ( .D(n1852), .CLK(CLOCK), .RSTB(n5284), .Q(
        \InstQueue[1][4] ) );
  DFFARX1 \InstQueue_reg[1][5]  ( .D(n1851), .CLK(CLOCK), .RSTB(n5284), .Q(
        \InstQueue[1][5] ) );
  DFFARX1 \InstQueue_reg[1][6]  ( .D(n1850), .CLK(CLOCK), .RSTB(n5284), .Q(
        \InstQueue[1][6] ) );
  DFFARX1 \InstQueue_reg[1][7]  ( .D(n1849), .CLK(CLOCK), .RSTB(n5284), .Q(
        \InstQueue[1][7] ) );
  DFFARX1 \InstQueue_reg[14][0]  ( .D(n1752), .CLK(CLOCK), .RSTB(n5284), .Q(
        \InstQueue[14][0] ), .QN(n5249) );
  DFFARX1 \InstQueue_reg[14][1]  ( .D(n1751), .CLK(CLOCK), .RSTB(n5285), .Q(
        \InstQueue[14][1] ) );
  DFFARX1 \InstQueue_reg[14][2]  ( .D(n1750), .CLK(CLOCK), .RSTB(n5285), .Q(
        \InstQueue[14][2] ) );
  DFFARX1 \InstQueue_reg[14][3]  ( .D(n1749), .CLK(CLOCK), .RSTB(n5285), .Q(
        \InstQueue[14][3] ) );
  DFFARX1 \InstQueue_reg[14][4]  ( .D(n1748), .CLK(CLOCK), .RSTB(n5285), .Q(
        \InstQueue[14][4] ) );
  DFFARX1 \InstQueue_reg[14][5]  ( .D(n1747), .CLK(CLOCK), .RSTB(n5285), .Q(
        \InstQueue[14][5] ) );
  DFFARX1 \InstQueue_reg[14][6]  ( .D(n1746), .CLK(CLOCK), .RSTB(n5285), .Q(
        \InstQueue[14][6] ) );
  DFFARX1 \InstQueue_reg[14][7]  ( .D(n1745), .CLK(CLOCK), .RSTB(n5285), .Q(
        \InstQueue[14][7] ) );
  DFFARX1 \InstQueue_reg[13][0]  ( .D(n1760), .CLK(CLOCK), .RSTB(n5285), .Q(
        \InstQueue[13][0] ) );
  DFFARX1 \InstQueue_reg[13][1]  ( .D(n1759), .CLK(CLOCK), .RSTB(n5285), .Q(
        \InstQueue[13][1] ) );
  DFFARX1 \InstQueue_reg[13][2]  ( .D(n1758), .CLK(CLOCK), .RSTB(n5285), .Q(
        \InstQueue[13][2] ) );
  DFFARX1 \InstQueue_reg[13][3]  ( .D(n1757), .CLK(CLOCK), .RSTB(n5285), .Q(
        \InstQueue[13][3] ) );
  DFFARX1 \InstQueue_reg[13][4]  ( .D(n1756), .CLK(CLOCK), .RSTB(n5285), .Q(
        \InstQueue[13][4] ) );
  DFFARX1 \InstQueue_reg[13][5]  ( .D(n1755), .CLK(CLOCK), .RSTB(n5286), .Q(
        \InstQueue[13][5] ) );
  DFFARX1 \InstQueue_reg[13][6]  ( .D(n1754), .CLK(CLOCK), .RSTB(n5286), .Q(
        \InstQueue[13][6] ) );
  DFFARX1 \InstQueue_reg[13][7]  ( .D(n1753), .CLK(CLOCK), .RSTB(n5286), .Q(
        \InstQueue[13][7] ) );
  DFFARX1 \InstQueue_reg[12][0]  ( .D(n1768), .CLK(CLOCK), .RSTB(n5286), .Q(
        \InstQueue[12][0] ) );
  DFFARX1 \InstQueue_reg[12][1]  ( .D(n1767), .CLK(CLOCK), .RSTB(n5286), .Q(
        \InstQueue[12][1] ) );
  DFFARX1 \InstQueue_reg[12][2]  ( .D(n1766), .CLK(CLOCK), .RSTB(n5286), .Q(
        \InstQueue[12][2] ) );
  DFFARX1 \InstQueue_reg[12][3]  ( .D(n1765), .CLK(CLOCK), .RSTB(n5286), .Q(
        \InstQueue[12][3] ) );
  DFFARX1 \InstQueue_reg[12][4]  ( .D(n1764), .CLK(CLOCK), .RSTB(n5286), .Q(
        \InstQueue[12][4] ) );
  DFFARX1 \InstQueue_reg[12][5]  ( .D(n1763), .CLK(CLOCK), .RSTB(n5286), .Q(
        \InstQueue[12][5] ) );
  DFFARX1 \InstQueue_reg[12][6]  ( .D(n1762), .CLK(CLOCK), .RSTB(n5286), .Q(
        \InstQueue[12][6] ) );
  DFFARX1 \InstQueue_reg[12][7]  ( .D(n1761), .CLK(CLOCK), .RSTB(n5286), .Q(
        \InstQueue[12][7] ) );
  DFFARX1 \InstQueue_reg[15][0]  ( .D(n1744), .CLK(CLOCK), .RSTB(n5286), .Q(
        \InstQueue[15][0] ), .QN(n5252) );
  DFFARX1 \InstQueue_reg[15][1]  ( .D(n1743), .CLK(CLOCK), .RSTB(n5287), .Q(
        \InstQueue[15][1] ) );
  DFFARX1 \InstQueue_reg[15][2]  ( .D(n1742), .CLK(CLOCK), .RSTB(n5287), .Q(
        \InstQueue[15][2] ) );
  DFFARX1 \InstQueue_reg[15][3]  ( .D(n1741), .CLK(CLOCK), .RSTB(n5287), .Q(
        \InstQueue[15][3] ) );
  DFFARX1 \InstQueue_reg[15][4]  ( .D(n1740), .CLK(CLOCK), .RSTB(n5287), .Q(
        \InstQueue[15][4] ) );
  DFFARX1 \InstQueue_reg[15][5]  ( .D(n1739), .CLK(CLOCK), .RSTB(n5287), .Q(
        \InstQueue[15][5] ) );
  DFFARX1 \InstQueue_reg[15][6]  ( .D(n1738), .CLK(CLOCK), .RSTB(n5287), .Q(
        \InstQueue[15][6] ) );
  DFFARX1 \InstQueue_reg[15][7]  ( .D(n1737), .CLK(CLOCK), .RSTB(n5287), .Q(
        \InstQueue[15][7] ) );
  DFFARX1 \DataWidth_reg[1]  ( .D(n1703), .CLK(CLOCK), .RSTB(n5287), .Q(
        DataWidth[1]) );
  DFFARX1 ADS_n_reg ( .D(n1669), .CLK(CLOCK), .RSTB(n5287), .Q(ADS_n) );
  DFFARX1 \BE_n_reg[3]  ( .D(n1668), .CLK(CLOCK), .RSTB(n5287), .Q(BE_n[3]) );
  DFFARX1 \BE_n_reg[2]  ( .D(n1667), .CLK(CLOCK), .RSTB(n5287), .Q(BE_n[2]) );
  DFFARX1 \BE_n_reg[1]  ( .D(n1666), .CLK(CLOCK), .RSTB(n5287), .Q(BE_n[1]) );
  DFFARX1 \BE_n_reg[0]  ( .D(n1664), .CLK(CLOCK), .RSTB(n5288), .Q(BE_n[0]) );
  DFFARX1 \ByteEnable_reg[3]  ( .D(n1663), .CLK(CLOCK), .RSTB(n5288), .Q(
        ByteEnable[3]) );
  DFFARX1 \ByteEnable_reg[2]  ( .D(n1662), .CLK(CLOCK), .RSTB(n5288), .Q(
        ByteEnable[2]) );
  DFFARX1 \ByteEnable_reg[1]  ( .D(n1661), .CLK(CLOCK), .RSTB(n5288), .Q(
        ByteEnable[1]) );
  DFFARX1 \ByteEnable_reg[0]  ( .D(n1660), .CLK(CLOCK), .RSTB(n5288), .Q(
        ByteEnable[0]) );
  HADDX1 \DP_OP_560J1_146_4463/U15  ( .A0(N1753), .B0(EAX[16]), .C1(
        \DP_OP_560J1_146_4463/n14 ), .SO(\C1/DATA1_16 ) );
  HADDX1 \DP_OP_560J1_146_4463/U14  ( .A0(\DP_OP_560J1_146_4463/n14 ), .B0(
        EAX[17]), .C1(\DP_OP_560J1_146_4463/n13 ), .SO(\C1/DATA1_17 ) );
  HADDX1 \DP_OP_560J1_146_4463/U13  ( .A0(\DP_OP_560J1_146_4463/n13 ), .B0(
        EAX[18]), .C1(\DP_OP_560J1_146_4463/n12 ), .SO(\C1/DATA1_18 ) );
  HADDX1 \DP_OP_560J1_146_4463/U12  ( .A0(\DP_OP_560J1_146_4463/n12 ), .B0(
        EAX[19]), .C1(\DP_OP_560J1_146_4463/n11 ), .SO(\C1/DATA1_19 ) );
  HADDX1 \DP_OP_560J1_146_4463/U11  ( .A0(\DP_OP_560J1_146_4463/n11 ), .B0(
        EAX[20]), .C1(\DP_OP_560J1_146_4463/n10 ), .SO(\C1/DATA1_20 ) );
  HADDX1 \DP_OP_560J1_146_4463/U10  ( .A0(\DP_OP_560J1_146_4463/n10 ), .B0(
        EAX[21]), .C1(\DP_OP_560J1_146_4463/n9 ), .SO(\C1/DATA1_21 ) );
  HADDX1 \DP_OP_560J1_146_4463/U9  ( .A0(\DP_OP_560J1_146_4463/n9 ), .B0(
        EAX[22]), .C1(\DP_OP_560J1_146_4463/n8 ), .SO(\C1/DATA1_22 ) );
  HADDX1 \DP_OP_560J1_146_4463/U8  ( .A0(\DP_OP_560J1_146_4463/n8 ), .B0(
        EAX[23]), .C1(\DP_OP_560J1_146_4463/n7 ), .SO(\C1/DATA1_23 ) );
  HADDX1 \DP_OP_560J1_146_4463/U7  ( .A0(\DP_OP_560J1_146_4463/n7 ), .B0(
        EAX[24]), .C1(\DP_OP_560J1_146_4463/n6 ), .SO(\C1/DATA1_24 ) );
  HADDX1 \DP_OP_560J1_146_4463/U6  ( .A0(\DP_OP_560J1_146_4463/n6 ), .B0(
        EAX[25]), .C1(\DP_OP_560J1_146_4463/n5 ), .SO(\C1/DATA1_25 ) );
  HADDX1 \DP_OP_560J1_146_4463/U5  ( .A0(\DP_OP_560J1_146_4463/n5 ), .B0(
        EAX[26]), .C1(\DP_OP_560J1_146_4463/n4 ), .SO(\C1/DATA1_26 ) );
  HADDX1 \DP_OP_560J1_146_4463/U4  ( .A0(\DP_OP_560J1_146_4463/n4 ), .B0(
        EAX[27]), .C1(\DP_OP_560J1_146_4463/n3 ), .SO(\C1/DATA1_27 ) );
  HADDX1 \DP_OP_560J1_146_4463/U3  ( .A0(\DP_OP_560J1_146_4463/n3 ), .B0(
        EAX[28]), .C1(\DP_OP_560J1_146_4463/n2 ), .SO(\C1/DATA1_28 ) );
  HADDX1 \DP_OP_560J1_146_4463/U2  ( .A0(\DP_OP_560J1_146_4463/n2 ), .B0(
        EAX[29]), .C1(\DP_OP_560J1_146_4463/n1 ), .SO(\C1/DATA1_29 ) );
  AND3X1 U2154 ( .IN1(n4280), .IN2(n4977), .IN3(n3314), .Q(n2090) );
  INVX0 U2155 ( .INP(RESET), .ZN(n5278) );
  INVX0 U2156 ( .INP(RESET), .ZN(n5277) );
  INVX0 U2157 ( .INP(RESET), .ZN(n5279) );
  INVX0 U2158 ( .INP(RESET), .ZN(n5280) );
  INVX0 U2159 ( .INP(RESET), .ZN(n5281) );
  INVX0 U2160 ( .INP(RESET), .ZN(n5289) );
  INVX0 U2161 ( .INP(RESET), .ZN(n5290) );
  INVX0 U2162 ( .INP(RESET), .ZN(n5291) );
  INVX0 U2163 ( .INP(RESET), .ZN(n5286) );
  INVX0 U2164 ( .INP(RESET), .ZN(n5284) );
  INVX0 U2165 ( .INP(RESET), .ZN(n5285) );
  INVX0 U2166 ( .INP(RESET), .ZN(n5283) );
  INVX0 U2167 ( .INP(RESET), .ZN(n5287) );
  INVX0 U2168 ( .INP(RESET), .ZN(n5288) );
  INVX0 U2169 ( .INP(RESET), .ZN(n5282) );
  NOR2X0 U2170 ( .IN1(N1351), .IN2(n5183), .QN(n2232) );
  INVX0 U2171 ( .INP(n2091), .ZN(n2304) );
  FADDX1 U2172 ( .A(InstQueueRd_Addr[1]), .B(n5182), .CI(n2232), .CO(n2092), 
        .S(n2091) );
  FADDX1 U2173 ( .A(InstQueueRd_Addr[2]), .B(n5198), .CI(n2092), .CO(n2094), 
        .S(n2235) );
  NOR2X0 U2174 ( .IN1(n2094), .IN2(n5200), .QN(n2093) );
  NAND2X0 U2175 ( .IN1(n2093), .IN2(n5206), .QN(n2236) );
  NAND2X0 U2176 ( .IN1(n2235), .IN2(n2236), .QN(n2306) );
  NAND2X0 U2177 ( .IN1(n5200), .IN2(InstQueueRd_Addr[3]), .QN(n2097) );
  NAND2X0 U2178 ( .IN1(N4186), .IN2(n5206), .QN(n2095) );
  NAND2X0 U2179 ( .IN1(n2095), .IN2(n2094), .QN(n2096) );
  NAND2X0 U2180 ( .IN1(n2097), .IN2(n2096), .QN(n2233) );
  INVX0 U2181 ( .INP(n2233), .ZN(n2303) );
  OA21X1 U2182 ( .IN1(n2304), .IN2(n2306), .IN3(n2303), .Q(n4515) );
  INVX0 U2183 ( .INP(n4515), .ZN(n2243) );
  NAND2X0 U2184 ( .IN1(n5177), .IN2(n5183), .QN(n2589) );
  NOR2X0 U2185 ( .IN1(InstQueueRd_Addr[2]), .IN2(InstQueueRd_Addr[3]), .QN(
        n2479) );
  INVX0 U2186 ( .INP(n2479), .ZN(n2323) );
  NOR2X0 U2187 ( .IN1(n2589), .IN2(n2323), .QN(n2547) );
  NAND2X0 U2188 ( .IN1(N2884), .IN2(n5177), .QN(n3020) );
  NOR2X0 U2189 ( .IN1(n2323), .IN2(n3020), .QN(n2168) );
  AO22X1 U2190 ( .IN1(n2547), .IN2(\DP_OP_469J1_133_8416/n117 ), .IN3(n2168), 
        .IN4(\InstQueue[1][1] ), .Q(n2101) );
  NAND2X0 U2191 ( .IN1(InstQueueRd_Addr[1]), .IN2(n5183), .QN(n3021) );
  NOR2X0 U2192 ( .IN1(n2323), .IN2(n3021), .QN(n2170) );
  NOR2X0 U2193 ( .IN1(n5180), .IN2(n5206), .QN(n2480) );
  INVX0 U2194 ( .INP(n2480), .ZN(n2262) );
  NOR2X0 U2195 ( .IN1(n5183), .IN2(n5177), .QN(n4306) );
  INVX0 U2196 ( .INP(n4306), .ZN(n4303) );
  NOR2X0 U2197 ( .IN1(n2262), .IN2(n4303), .QN(n2169) );
  AO22X1 U2198 ( .IN1(n2170), .IN2(\InstQueue[2][1] ), .IN3(n2169), .IN4(
        \InstQueue[15][1] ), .Q(n2100) );
  NOR2X0 U2199 ( .IN1(n2323), .IN2(n4303), .QN(n2592) );
  NOR2X0 U2200 ( .IN1(n5180), .IN2(InstQueueRd_Addr[3]), .QN(n2481) );
  INVX0 U2201 ( .INP(n2481), .ZN(n2260) );
  NOR2X0 U2202 ( .IN1(n2589), .IN2(n2260), .QN(n2498) );
  AO22X1 U2203 ( .IN1(n2592), .IN2(\InstQueue[3][1] ), .IN3(n2498), .IN4(
        \InstQueue[4][1] ), .Q(n2099) );
  NOR2X0 U2204 ( .IN1(n3020), .IN2(n2260), .QN(n2172) );
  NOR2X0 U2205 ( .IN1(n3021), .IN2(n2260), .QN(n2171) );
  AO22X1 U2206 ( .IN1(n2172), .IN2(\InstQueue[5][1] ), .IN3(n2171), .IN4(
        \InstQueue[6][1] ), .Q(n2098) );
  OR4X1 U2207 ( .IN1(n2101), .IN2(n2100), .IN3(n2099), .IN4(n2098), .Q(n2107)
         );
  NOR2X0 U2208 ( .IN1(n2260), .IN2(n4303), .QN(n2588) );
  NOR2X0 U2209 ( .IN1(n5206), .IN2(InstQueueRd_Addr[2]), .QN(n2478) );
  INVX0 U2210 ( .INP(n2478), .ZN(n2324) );
  NOR2X0 U2211 ( .IN1(n2324), .IN2(n2589), .QN(n2500) );
  AO22X1 U2212 ( .IN1(n2588), .IN2(\InstQueue[7][1] ), .IN3(n2500), .IN4(
        \InstQueue[8][1] ), .Q(n2105) );
  NOR2X0 U2213 ( .IN1(n3020), .IN2(n2324), .QN(n2178) );
  NOR2X0 U2214 ( .IN1(n3021), .IN2(n2324), .QN(n2177) );
  AO22X1 U2215 ( .IN1(n2178), .IN2(\InstQueue[9][1] ), .IN3(n2177), .IN4(
        \InstQueue[10][1] ), .Q(n2104) );
  NOR2X0 U2216 ( .IN1(n2324), .IN2(n4303), .QN(n2180) );
  NOR2X0 U2217 ( .IN1(n3021), .IN2(n2262), .QN(n2179) );
  AO22X1 U2218 ( .IN1(n2180), .IN2(\InstQueue[11][1] ), .IN3(n2179), .IN4(
        \InstQueue[14][1] ), .Q(n2103) );
  NOR2X0 U2219 ( .IN1(n2589), .IN2(n2262), .QN(n2546) );
  NOR2X0 U2220 ( .IN1(n2262), .IN2(n3020), .QN(n2181) );
  AO22X1 U2221 ( .IN1(n2546), .IN2(\InstQueue[12][1] ), .IN3(n2181), .IN4(
        \InstQueue[13][1] ), .Q(n2102) );
  OR4X1 U2222 ( .IN1(n2105), .IN2(n2104), .IN3(n2103), .IN4(n2102), .Q(n2106)
         );
  OR2X1 U2223 ( .IN1(n2107), .IN2(n2106), .Q(n2998) );
  NAND3X0 U2224 ( .IN1(State2[2]), .IN2(n5179), .IN3(n5242), .QN(n2239) );
  NOR2X0 U2225 ( .IN1(n5176), .IN2(n2239), .QN(n4445) );
  INVX0 U2226 ( .INP(n4445), .ZN(n4519) );
  AO22X1 U2227 ( .IN1(n2547), .IN2(\DP_OP_469J1_133_8416/n116 ), .IN3(n2168), 
        .IN4(\InstQueue[1][0] ), .Q(n2111) );
  AO22X1 U2228 ( .IN1(n2170), .IN2(\InstQueue[2][0] ), .IN3(n2169), .IN4(
        \InstQueue[15][0] ), .Q(n2110) );
  AO22X1 U2229 ( .IN1(n2592), .IN2(\InstQueue[3][0] ), .IN3(n2498), .IN4(
        \InstQueue[4][0] ), .Q(n2109) );
  AO22X1 U2230 ( .IN1(n2172), .IN2(\InstQueue[5][0] ), .IN3(n2171), .IN4(
        \InstQueue[6][0] ), .Q(n2108) );
  OR4X1 U2231 ( .IN1(n2111), .IN2(n2110), .IN3(n2109), .IN4(n2108), .Q(n2117)
         );
  AO22X1 U2232 ( .IN1(n2588), .IN2(\InstQueue[7][0] ), .IN3(n2500), .IN4(
        \InstQueue[8][0] ), .Q(n2115) );
  AO22X1 U2233 ( .IN1(n2178), .IN2(\InstQueue[9][0] ), .IN3(n2177), .IN4(
        \InstQueue[10][0] ), .Q(n2114) );
  AO22X1 U2234 ( .IN1(n2180), .IN2(\InstQueue[11][0] ), .IN3(n2179), .IN4(
        \InstQueue[14][0] ), .Q(n2113) );
  AO22X1 U2235 ( .IN1(n2546), .IN2(\InstQueue[12][0] ), .IN3(n2181), .IN4(
        \InstQueue[13][0] ), .Q(n2112) );
  OR4X1 U2236 ( .IN1(n2115), .IN2(n2114), .IN3(n2113), .IN4(n2112), .Q(n2116)
         );
  NOR2X0 U2237 ( .IN1(n2117), .IN2(n2116), .QN(n3026) );
  AO22X1 U2238 ( .IN1(\DP_OP_469J1_133_8416/n119 ), .IN2(n2547), .IN3(
        \InstQueue[1][3] ), .IN4(n2168), .Q(n2121) );
  AO22X1 U2239 ( .IN1(\InstQueue[2][3] ), .IN2(n2170), .IN3(\InstQueue[15][3] ), .IN4(n2169), .Q(n2120) );
  AO22X1 U2240 ( .IN1(\InstQueue[3][3] ), .IN2(n2592), .IN3(\InstQueue[4][3] ), 
        .IN4(n2498), .Q(n2119) );
  AO22X1 U2241 ( .IN1(\InstQueue[5][3] ), .IN2(n2172), .IN3(\InstQueue[6][3] ), 
        .IN4(n2171), .Q(n2118) );
  OR4X1 U2242 ( .IN1(n2121), .IN2(n2120), .IN3(n2119), .IN4(n2118), .Q(n2127)
         );
  AO22X1 U2243 ( .IN1(\InstQueue[7][3] ), .IN2(n2588), .IN3(\InstQueue[8][3] ), 
        .IN4(n2500), .Q(n2125) );
  AO22X1 U2244 ( .IN1(\InstQueue[9][3] ), .IN2(n2178), .IN3(\InstQueue[10][3] ), .IN4(n2177), .Q(n2124) );
  AO22X1 U2245 ( .IN1(\InstQueue[11][3] ), .IN2(n2180), .IN3(
        \InstQueue[14][3] ), .IN4(n2179), .Q(n2123) );
  AO22X1 U2246 ( .IN1(\InstQueue[12][3] ), .IN2(n2546), .IN3(
        \InstQueue[13][3] ), .IN4(n2181), .Q(n2122) );
  OR4X1 U2247 ( .IN1(n2125), .IN2(n2124), .IN3(n2123), .IN4(n2122), .Q(n2126)
         );
  OR2X1 U2248 ( .IN1(n2127), .IN2(n2126), .Q(n2979) );
  INVX0 U2249 ( .INP(n2979), .ZN(n2319) );
  AO22X1 U2250 ( .IN1(n2588), .IN2(\InstQueue[7][7] ), .IN3(n2500), .IN4(
        \InstQueue[8][7] ), .Q(n2131) );
  AO22X1 U2251 ( .IN1(n2178), .IN2(\InstQueue[9][7] ), .IN3(n2177), .IN4(
        \InstQueue[10][7] ), .Q(n2130) );
  AO22X1 U2252 ( .IN1(n2180), .IN2(\InstQueue[11][7] ), .IN3(n2179), .IN4(
        \InstQueue[14][7] ), .Q(n2129) );
  AO22X1 U2253 ( .IN1(n2546), .IN2(\InstQueue[12][7] ), .IN3(n2181), .IN4(
        \InstQueue[13][7] ), .Q(n2128) );
  OR4X1 U2254 ( .IN1(n2131), .IN2(n2130), .IN3(n2129), .IN4(n2128), .Q(n2137)
         );
  AO22X1 U2255 ( .IN1(n2547), .IN2(\DP_OP_469J1_133_8416/n123 ), .IN3(n2168), 
        .IN4(\InstQueue[1][7] ), .Q(n2135) );
  AO22X1 U2256 ( .IN1(n2170), .IN2(\InstQueue[2][7] ), .IN3(n2169), .IN4(
        \InstQueue[15][7] ), .Q(n2134) );
  AO22X1 U2257 ( .IN1(n2592), .IN2(\InstQueue[3][7] ), .IN3(n2498), .IN4(
        \InstQueue[4][7] ), .Q(n2133) );
  AO22X1 U2258 ( .IN1(n2172), .IN2(\InstQueue[5][7] ), .IN3(n2171), .IN4(
        \InstQueue[6][7] ), .Q(n2132) );
  OR4X1 U2259 ( .IN1(n2135), .IN2(n2134), .IN3(n2133), .IN4(n2132), .Q(n2136)
         );
  NOR2X0 U2260 ( .IN1(n2137), .IN2(n2136), .QN(n2941) );
  AO22X1 U2261 ( .IN1(n2547), .IN2(\DP_OP_469J1_133_8416/n118 ), .IN3(n2168), 
        .IN4(\InstQueue[1][2] ), .Q(n2141) );
  AO22X1 U2262 ( .IN1(n2170), .IN2(\InstQueue[2][2] ), .IN3(n2169), .IN4(
        \InstQueue[15][2] ), .Q(n2140) );
  AO22X1 U2263 ( .IN1(n2592), .IN2(\InstQueue[3][2] ), .IN3(n2498), .IN4(
        \InstQueue[4][2] ), .Q(n2139) );
  AO22X1 U2264 ( .IN1(n2172), .IN2(\InstQueue[5][2] ), .IN3(n2171), .IN4(
        \InstQueue[6][2] ), .Q(n2138) );
  NOR4X0 U2265 ( .IN1(n2141), .IN2(n2140), .IN3(n2139), .IN4(n2138), .QN(n2147) );
  AO22X1 U2266 ( .IN1(n2588), .IN2(\InstQueue[7][2] ), .IN3(n2500), .IN4(
        \InstQueue[8][2] ), .Q(n2145) );
  AO22X1 U2267 ( .IN1(n2178), .IN2(\InstQueue[9][2] ), .IN3(n2177), .IN4(
        \InstQueue[10][2] ), .Q(n2144) );
  AO22X1 U2268 ( .IN1(n2180), .IN2(\InstQueue[11][2] ), .IN3(n2179), .IN4(
        \InstQueue[14][2] ), .Q(n2143) );
  AO22X1 U2269 ( .IN1(n2546), .IN2(\InstQueue[12][2] ), .IN3(n2181), .IN4(
        \InstQueue[13][2] ), .Q(n2142) );
  NOR4X0 U2270 ( .IN1(n2145), .IN2(n2144), .IN3(n2143), .IN4(n2142), .QN(n2146) );
  NAND2X0 U2271 ( .IN1(n2147), .IN2(n2146), .QN(n2987) );
  OR2X1 U2272 ( .IN1(n2941), .IN2(n2987), .Q(n2237) );
  NOR3X0 U2273 ( .IN1(n3026), .IN2(n2319), .IN3(n2237), .QN(n2300) );
  INVX0 U2274 ( .INP(n2300), .ZN(n2302) );
  AO22X1 U2275 ( .IN1(n2588), .IN2(\InstQueue[7][6] ), .IN3(n2500), .IN4(
        \InstQueue[8][6] ), .Q(n2151) );
  AO22X1 U2276 ( .IN1(n2178), .IN2(\InstQueue[9][6] ), .IN3(n2177), .IN4(
        \InstQueue[10][6] ), .Q(n2150) );
  AO22X1 U2277 ( .IN1(n2180), .IN2(\InstQueue[11][6] ), .IN3(n2179), .IN4(
        \InstQueue[14][6] ), .Q(n2149) );
  AO22X1 U2278 ( .IN1(n2546), .IN2(\InstQueue[12][6] ), .IN3(n2181), .IN4(
        \InstQueue[13][6] ), .Q(n2148) );
  OR4X1 U2279 ( .IN1(n2151), .IN2(n2150), .IN3(n2149), .IN4(n2148), .Q(n2157)
         );
  AO22X1 U2280 ( .IN1(n2547), .IN2(\DP_OP_469J1_133_8416/n122 ), .IN3(n2168), 
        .IN4(\InstQueue[1][6] ), .Q(n2155) );
  AO22X1 U2281 ( .IN1(n2170), .IN2(\InstQueue[2][6] ), .IN3(n2169), .IN4(
        \InstQueue[15][6] ), .Q(n2154) );
  AO22X1 U2282 ( .IN1(n2592), .IN2(\InstQueue[3][6] ), .IN3(n2498), .IN4(
        \InstQueue[4][6] ), .Q(n2153) );
  AO22X1 U2283 ( .IN1(n2172), .IN2(\InstQueue[5][6] ), .IN3(n2171), .IN4(
        \InstQueue[6][6] ), .Q(n2152) );
  OR4X1 U2284 ( .IN1(n2155), .IN2(n2154), .IN3(n2153), .IN4(n2152), .Q(n2156)
         );
  NOR2X0 U2285 ( .IN1(n2157), .IN2(n2156), .QN(n2244) );
  INVX0 U2286 ( .INP(n2244), .ZN(n2955) );
  AO22X1 U2287 ( .IN1(n2588), .IN2(\InstQueue[7][5] ), .IN3(n2500), .IN4(
        \InstQueue[8][5] ), .Q(n2161) );
  AO22X1 U2288 ( .IN1(n2178), .IN2(\InstQueue[9][5] ), .IN3(n2177), .IN4(
        \InstQueue[10][5] ), .Q(n2160) );
  AO22X1 U2289 ( .IN1(n2180), .IN2(\InstQueue[11][5] ), .IN3(n2179), .IN4(
        \InstQueue[14][5] ), .Q(n2159) );
  AO22X1 U2290 ( .IN1(n2546), .IN2(\InstQueue[12][5] ), .IN3(n2181), .IN4(
        \InstQueue[13][5] ), .Q(n2158) );
  OR4X1 U2291 ( .IN1(n2161), .IN2(n2160), .IN3(n2159), .IN4(n2158), .Q(n2167)
         );
  AO22X1 U2292 ( .IN1(n2547), .IN2(\DP_OP_469J1_133_8416/n121 ), .IN3(n2168), 
        .IN4(\InstQueue[1][5] ), .Q(n2165) );
  AO22X1 U2293 ( .IN1(n2170), .IN2(\InstQueue[2][5] ), .IN3(n2169), .IN4(
        \InstQueue[15][5] ), .Q(n2164) );
  AO22X1 U2294 ( .IN1(n2592), .IN2(\InstQueue[3][5] ), .IN3(n2498), .IN4(
        \InstQueue[4][5] ), .Q(n2163) );
  AO22X1 U2295 ( .IN1(n2172), .IN2(\InstQueue[5][5] ), .IN3(n2171), .IN4(
        \InstQueue[6][5] ), .Q(n2162) );
  OR4X1 U2296 ( .IN1(n2165), .IN2(n2164), .IN3(n2163), .IN4(n2162), .Q(n2166)
         );
  NOR2X0 U2297 ( .IN1(n2167), .IN2(n2166), .QN(n2316) );
  INVX0 U2298 ( .INP(n2316), .ZN(n2966) );
  AO22X1 U2299 ( .IN1(n2547), .IN2(\DP_OP_469J1_133_8416/n120 ), .IN3(n2168), 
        .IN4(\InstQueue[1][4] ), .Q(n2176) );
  AO22X1 U2300 ( .IN1(n2170), .IN2(\InstQueue[2][4] ), .IN3(n2169), .IN4(
        \InstQueue[15][4] ), .Q(n2175) );
  AO22X1 U2301 ( .IN1(n2592), .IN2(\InstQueue[3][4] ), .IN3(n2498), .IN4(
        \InstQueue[4][4] ), .Q(n2174) );
  AO22X1 U2302 ( .IN1(n2172), .IN2(\InstQueue[5][4] ), .IN3(n2171), .IN4(
        \InstQueue[6][4] ), .Q(n2173) );
  OR4X1 U2303 ( .IN1(n2176), .IN2(n2175), .IN3(n2174), .IN4(n2173), .Q(n2187)
         );
  AO22X1 U2304 ( .IN1(n2588), .IN2(\InstQueue[7][4] ), .IN3(n2500), .IN4(
        \InstQueue[8][4] ), .Q(n2185) );
  AO22X1 U2305 ( .IN1(n2178), .IN2(\InstQueue[9][4] ), .IN3(n2177), .IN4(
        \InstQueue[10][4] ), .Q(n2184) );
  AO22X1 U2306 ( .IN1(n2180), .IN2(\InstQueue[11][4] ), .IN3(n2179), .IN4(
        \InstQueue[14][4] ), .Q(n2183) );
  AO22X1 U2307 ( .IN1(n2546), .IN2(\InstQueue[12][4] ), .IN3(n2181), .IN4(
        \InstQueue[13][4] ), .Q(n2182) );
  OR4X1 U2308 ( .IN1(n2185), .IN2(n2184), .IN3(n2183), .IN4(n2182), .Q(n2186)
         );
  NOR2X0 U2309 ( .IN1(n2187), .IN2(n2186), .QN(n2318) );
  INVX0 U2310 ( .INP(n2318), .ZN(n2971) );
  NOR4X0 U2311 ( .IN1(n2302), .IN2(n2955), .IN3(n2966), .IN4(n2971), .QN(n2246) );
  INVX0 U2312 ( .INP(n2246), .ZN(n2188) );
  NOR2X0 U2313 ( .IN1(n4519), .IN2(n2188), .QN(n4486) );
  INVX0 U2314 ( .INP(n4486), .ZN(n2189) );
  NOR2X0 U2315 ( .IN1(n2998), .IN2(n2189), .QN(n4443) );
  INVX0 U2316 ( .INP(n4443), .ZN(n4521) );
  INVX0 U2317 ( .INP(READY_n), .ZN(n4469) );
  NAND2X0 U2318 ( .IN1(n4515), .IN2(n4469), .QN(n2314) );
  NAND2X0 U2319 ( .IN1(n2246), .IN2(n2998), .QN(n2256) );
  INVX0 U2320 ( .INP(n2256), .ZN(n2599) );
  NAND2X0 U2321 ( .IN1(n2599), .IN2(n4445), .QN(n3284) );
  OA22X1 U2322 ( .IN1(n2243), .IN2(n4521), .IN3(n2314), .IN4(n3284), .Q(n4319)
         );
  NOR2X0 U2323 ( .IN1(n4319), .IN2(n2998), .QN(n4318) );
  AOI22X1 U2324 ( .IN1(n4319), .IN2(\C1/DATA2_29 ), .IN3(n4318), .IN4(
        \C1/DATA1_29 ), .QN(n2190) );
  NOR2X0 U2325 ( .IN1(n4319), .IN2(n2256), .QN(n4320) );
  NAND2X0 U2326 ( .IN1(Datai[13]), .IN2(n4320), .QN(n2223) );
  NAND2X0 U2327 ( .IN1(n2190), .IN2(n2223), .QN(n1945) );
  MUX21X1 U2328 ( .IN1(EAX[30]), .IN2(n5262), .S(\DP_OP_560J1_146_4463/n1 ), 
        .Q(n4524) );
  AOI22X1 U2329 ( .IN1(n4319), .IN2(\C1/DATA2_30 ), .IN3(n4318), .IN4(n4524), 
        .QN(n2191) );
  NAND2X0 U2330 ( .IN1(Datai[14]), .IN2(n4320), .QN(n2227) );
  NAND2X0 U2331 ( .IN1(n2191), .IN2(n2227), .QN(n1944) );
  AOI22X1 U2332 ( .IN1(n4319), .IN2(\C1/DATA2_27 ), .IN3(n4318), .IN4(
        \C1/DATA1_27 ), .QN(n2192) );
  NAND2X0 U2333 ( .IN1(Datai[11]), .IN2(n4320), .QN(n2218) );
  NAND2X0 U2334 ( .IN1(n2192), .IN2(n2218), .QN(n1947) );
  AOI22X1 U2335 ( .IN1(EAX[0]), .IN2(n4318), .IN3(n4319), .IN4(\C1/DATA2_0 ), 
        .QN(n2193) );
  NAND2X0 U2336 ( .IN1(Datai[0]), .IN2(n4320), .QN(n2297) );
  NAND2X0 U2337 ( .IN1(n2193), .IN2(n2297), .QN(n1943) );
  AOI22X1 U2338 ( .IN1(EAX[1]), .IN2(n4318), .IN3(n4319), .IN4(\C1/DATA2_1 ), 
        .QN(n2194) );
  NAND2X0 U2339 ( .IN1(Datai[1]), .IN2(n4320), .QN(n2229) );
  NAND2X0 U2340 ( .IN1(n2194), .IN2(n2229), .QN(n1942) );
  AOI22X1 U2341 ( .IN1(n4319), .IN2(\C1/DATA2_26 ), .IN3(n4318), .IN4(
        \C1/DATA1_26 ), .QN(n2195) );
  NAND2X0 U2342 ( .IN1(Datai[10]), .IN2(n4320), .QN(n2214) );
  NAND2X0 U2343 ( .IN1(n2195), .IN2(n2214), .QN(n1948) );
  AOI22X1 U2344 ( .IN1(EAX[2]), .IN2(n4318), .IN3(n4319), .IN4(\C1/DATA2_2 ), 
        .QN(n2196) );
  NAND2X0 U2345 ( .IN1(Datai[2]), .IN2(n4320), .QN(n2225) );
  NAND2X0 U2346 ( .IN1(n2196), .IN2(n2225), .QN(n1941) );
  AOI22X1 U2347 ( .IN1(n4319), .IN2(\C1/DATA2_25 ), .IN3(n4318), .IN4(
        \C1/DATA1_25 ), .QN(n2197) );
  NAND2X0 U2348 ( .IN1(Datai[9]), .IN2(n4320), .QN(n2212) );
  NAND2X0 U2349 ( .IN1(n2197), .IN2(n2212), .QN(n1949) );
  AOI22X1 U2350 ( .IN1(EAX[3]), .IN2(n4318), .IN3(n4319), .IN4(\C1/DATA2_3 ), 
        .QN(n2198) );
  NAND2X0 U2351 ( .IN1(Datai[3]), .IN2(n4320), .QN(n2220) );
  NAND2X0 U2352 ( .IN1(n2198), .IN2(n2220), .QN(n1940) );
  AOI22X1 U2353 ( .IN1(EAX[4]), .IN2(n4318), .IN3(n4319), .IN4(\C1/DATA2_4 ), 
        .QN(n2199) );
  NAND2X0 U2354 ( .IN1(Datai[4]), .IN2(n4320), .QN(n2216) );
  NAND2X0 U2355 ( .IN1(n2199), .IN2(n2216), .QN(n1939) );
  AOI22X1 U2356 ( .IN1(n4319), .IN2(\C1/DATA2_24 ), .IN3(n4318), .IN4(
        \C1/DATA1_24 ), .QN(n2200) );
  NAND2X0 U2357 ( .IN1(Datai[8]), .IN2(n4320), .QN(n2208) );
  NAND2X0 U2358 ( .IN1(n2200), .IN2(n2208), .QN(n1950) );
  AOI22X1 U2359 ( .IN1(EAX[5]), .IN2(n4318), .IN3(n4319), .IN4(\C1/DATA2_5 ), 
        .QN(n2201) );
  NAND2X0 U2360 ( .IN1(Datai[5]), .IN2(n4320), .QN(n2210) );
  NAND2X0 U2361 ( .IN1(n2201), .IN2(n2210), .QN(n1938) );
  AOI22X1 U2362 ( .IN1(n4319), .IN2(\C1/DATA2_23 ), .IN3(n4318), .IN4(
        \C1/DATA1_23 ), .QN(n2202) );
  NAND2X0 U2363 ( .IN1(Datai[7]), .IN2(n4320), .QN(n2204) );
  NAND2X0 U2364 ( .IN1(n2202), .IN2(n2204), .QN(n1951) );
  AOI22X1 U2365 ( .IN1(EAX[6]), .IN2(n4318), .IN3(n4319), .IN4(\C1/DATA2_6 ), 
        .QN(n2203) );
  NAND2X0 U2366 ( .IN1(Datai[6]), .IN2(n4320), .QN(n2206) );
  NAND2X0 U2367 ( .IN1(n2203), .IN2(n2206), .QN(n1937) );
  AOI22X1 U2368 ( .IN1(EAX[7]), .IN2(n4318), .IN3(n4319), .IN4(\C1/DATA2_7 ), 
        .QN(n2205) );
  NAND2X0 U2369 ( .IN1(n2205), .IN2(n2204), .QN(n1936) );
  AOI22X1 U2370 ( .IN1(n4319), .IN2(\C1/DATA2_22 ), .IN3(n4318), .IN4(
        \C1/DATA1_22 ), .QN(n2207) );
  NAND2X0 U2371 ( .IN1(n2207), .IN2(n2206), .QN(n1952) );
  AOI22X1 U2372 ( .IN1(EAX[8]), .IN2(n4318), .IN3(n4319), .IN4(\C1/DATA2_8 ), 
        .QN(n2209) );
  NAND2X0 U2373 ( .IN1(n2209), .IN2(n2208), .QN(n1935) );
  AOI22X1 U2374 ( .IN1(n4319), .IN2(\C1/DATA2_21 ), .IN3(n4318), .IN4(
        \C1/DATA1_21 ), .QN(n2211) );
  NAND2X0 U2375 ( .IN1(n2211), .IN2(n2210), .QN(n1953) );
  AOI22X1 U2376 ( .IN1(EAX[9]), .IN2(n4318), .IN3(n4319), .IN4(\C1/DATA2_9 ), 
        .QN(n2213) );
  NAND2X0 U2377 ( .IN1(n2213), .IN2(n2212), .QN(n1934) );
  AOI22X1 U2378 ( .IN1(EAX[10]), .IN2(n4318), .IN3(n4319), .IN4(\C1/DATA2_10 ), 
        .QN(n2215) );
  NAND2X0 U2379 ( .IN1(n2215), .IN2(n2214), .QN(n1933) );
  AOI22X1 U2380 ( .IN1(n4319), .IN2(\C1/DATA2_20 ), .IN3(n4318), .IN4(
        \C1/DATA1_20 ), .QN(n2217) );
  NAND2X0 U2381 ( .IN1(n2217), .IN2(n2216), .QN(n1954) );
  AOI22X1 U2382 ( .IN1(EAX[11]), .IN2(n4318), .IN3(n4319), .IN4(\C1/DATA2_11 ), 
        .QN(n2219) );
  NAND2X0 U2383 ( .IN1(n2219), .IN2(n2218), .QN(n1932) );
  AOI22X1 U2384 ( .IN1(n4319), .IN2(\C1/DATA2_19 ), .IN3(n4318), .IN4(
        \C1/DATA1_19 ), .QN(n2221) );
  NAND2X0 U2385 ( .IN1(n2221), .IN2(n2220), .QN(n1955) );
  AOI22X1 U2386 ( .IN1(EAX[12]), .IN2(n4318), .IN3(n4319), .IN4(\C1/DATA2_12 ), 
        .QN(n2222) );
  NAND2X0 U2387 ( .IN1(Datai[12]), .IN2(n4320), .QN(n2664) );
  NAND2X0 U2388 ( .IN1(n2222), .IN2(n2664), .QN(n1931) );
  AOI22X1 U2389 ( .IN1(EAX[13]), .IN2(n4318), .IN3(n4319), .IN4(\C1/DATA2_13 ), 
        .QN(n2224) );
  NAND2X0 U2390 ( .IN1(n2224), .IN2(n2223), .QN(n1930) );
  AOI22X1 U2391 ( .IN1(n4319), .IN2(\C1/DATA2_18 ), .IN3(n4318), .IN4(
        \C1/DATA1_18 ), .QN(n2226) );
  NAND2X0 U2392 ( .IN1(n2226), .IN2(n2225), .QN(n1956) );
  AOI22X1 U2393 ( .IN1(EAX[14]), .IN2(n4318), .IN3(n4319), .IN4(\C1/DATA2_14 ), 
        .QN(n2228) );
  NAND2X0 U2394 ( .IN1(n2228), .IN2(n2227), .QN(n1929) );
  AOI22X1 U2395 ( .IN1(n4319), .IN2(\C1/DATA2_17 ), .IN3(n4318), .IN4(
        \C1/DATA1_17 ), .QN(n2230) );
  NAND2X0 U2396 ( .IN1(n2230), .IN2(n2229), .QN(n1957) );
  NAND2X0 U2397 ( .IN1(n2589), .IN2(n5208), .QN(n2231) );
  NOR2X0 U2398 ( .IN1(n2262), .IN2(n2231), .QN(n4493) );
  NAND3X0 U2399 ( .IN1(State2[0]), .IN2(State2[2]), .IN3(State2[1]), .QN(n4466) );
  NAND3X0 U2400 ( .IN1(State2[0]), .IN2(n5179), .IN3(n5236), .QN(n4468) );
  OA22X1 U2401 ( .IN1(n4493), .IN2(n4466), .IN3(n4469), .IN4(n4468), .Q(n2296)
         );
  NAND4X0 U2402 ( .IN1(State2[2]), .IN2(State2[1]), .IN3(n5176), .IN4(n5179), 
        .QN(n4516) );
  AO21X1 U2403 ( .IN1(N1351), .IN2(n5183), .IN3(n2232), .Q(n2305) );
  NOR2X0 U2404 ( .IN1(n2305), .IN2(n2304), .QN(n2234) );
  AO221X1 U2405 ( .IN1(n2236), .IN2(n2235), .IN3(n2236), .IN4(n2234), .IN5(
        n2233), .Q(n2785) );
  INVX0 U2406 ( .INP(n2785), .ZN(n3052) );
  NOR2X0 U2407 ( .IN1(n2318), .IN2(n2955), .QN(n2238) );
  AND4X1 U2408 ( .IN1(n2300), .IN2(n2238), .IN3(n2998), .IN4(n2966), .Q(n3053)
         );
  INVX0 U2409 ( .INP(n2998), .ZN(n3027) );
  NAND2X0 U2410 ( .IN1(n3027), .IN2(n3026), .QN(n2320) );
  NOR2X0 U2411 ( .IN1(n2237), .IN2(n2320), .QN(n2247) );
  NAND4X0 U2412 ( .IN1(n2247), .IN2(n2238), .IN3(n2979), .IN4(n2966), .QN(
        n2313) );
  INVX0 U2413 ( .INP(n2313), .ZN(n2600) );
  NOR2X0 U2414 ( .IN1(n3053), .IN2(n2600), .QN(n2266) );
  NOR3X0 U2415 ( .IN1(n4519), .IN2(n3052), .IN3(n2266), .QN(n2310) );
  NAND2X0 U2416 ( .IN1(n5236), .IN2(n5242), .QN(n2940) );
  NOR2X0 U2417 ( .IN1(State2[3]), .IN2(n2940), .QN(n4487) );
  INVX0 U2418 ( .INP(n4487), .ZN(n4447) );
  NOR2X0 U2419 ( .IN1(n4447), .IN2(State2[0]), .QN(n4104) );
  NOR4X0 U2420 ( .IN1(State2[3]), .IN2(State2[0]), .IN3(State2[2]), .IN4(n5242), .QN(n4977) );
  INVX0 U2421 ( .INP(n4977), .ZN(n5101) );
  OR2X1 U2422 ( .IN1(State2[0]), .IN2(n2239), .Q(n4479) );
  NAND2X0 U2423 ( .IN1(n5101), .IN2(n4479), .QN(n5096) );
  NOR2X0 U2424 ( .IN1(n4104), .IN2(n5096), .QN(n4450) );
  NOR2X0 U2425 ( .IN1(n5179), .IN2(n2940), .QN(n2240) );
  NAND2X0 U2426 ( .IN1(State2[0]), .IN2(n2240), .QN(n3288) );
  INVX0 U2427 ( .INP(n2987), .ZN(n2317) );
  INVX0 U2428 ( .INP(n3026), .ZN(n2241) );
  NOR4X0 U2429 ( .IN1(n2941), .IN2(n2317), .IN3(n2241), .IN4(n2979), .QN(n2249) );
  INVX0 U2430 ( .INP(n2249), .ZN(n2245) );
  NAND4X0 U2431 ( .IN1(n2318), .IN2(n4445), .IN3(n2955), .IN4(n2966), .QN(
        n2242) );
  NOR2X0 U2432 ( .IN1(n2245), .IN2(n2242), .QN(n4277) );
  OR2X1 U2433 ( .IN1(n4486), .IN2(n4277), .Q(n3178) );
  NAND2X0 U2434 ( .IN1(n2243), .IN2(n3178), .QN(n2311) );
  NOR4X0 U2435 ( .IN1(n2244), .IN2(n2316), .IN3(n2971), .IN4(n2302), .QN(n2286) );
  NAND3X0 U2436 ( .IN1(n2318), .IN2(n2955), .IN3(n2966), .QN(n2248) );
  OR2X1 U2437 ( .IN1(n3027), .IN2(n2248), .Q(n2301) );
  NOR2X0 U2438 ( .IN1(n2301), .IN2(n2245), .QN(n4444) );
  NOR2X0 U2439 ( .IN1(n2246), .IN2(n4444), .QN(n2257) );
  NAND4X0 U2440 ( .IN1(n2319), .IN2(n2316), .IN3(n2247), .IN4(n2955), .QN(
        n2258) );
  INVX0 U2441 ( .INP(n2258), .ZN(n2926) );
  NOR2X0 U2442 ( .IN1(n2926), .IN2(n2286), .QN(n2269) );
  NOR2X0 U2443 ( .IN1(n2998), .IN2(n2248), .QN(n2299) );
  NAND2X0 U2444 ( .IN1(n2299), .IN2(n2249), .QN(n2322) );
  NAND4X0 U2445 ( .IN1(n2257), .IN2(n2266), .IN3(n2269), .IN4(n2322), .QN(
        n2783) );
  NAND3X0 U2446 ( .IN1(n2257), .IN2(n2322), .IN3(n2258), .QN(n2276) );
  NAND2X0 U2447 ( .IN1(n5177), .IN2(n2276), .QN(n2271) );
  OAI221X1 U2448 ( .IN1(n4303), .IN2(n2266), .IN3(n4306), .IN4(n2783), .IN5(
        n2271), .QN(n2254) );
  INVX0 U2449 ( .INP(n2783), .ZN(n2263) );
  INVX0 U2450 ( .INP(n2266), .ZN(n2923) );
  AND2X1 U2451 ( .IN1(n2257), .IN2(n2258), .Q(n2250) );
  NOR2X0 U2452 ( .IN1(n2250), .IN2(n5177), .QN(n2251) );
  AO221X1 U2453 ( .IN1(n4306), .IN2(n2263), .IN3(n4303), .IN4(n2923), .IN5(
        n2251), .Q(n2253) );
  NOR3X0 U2454 ( .IN1(n5177), .IN2(n2322), .IN3(InstQueueRd_Addr[2]), .QN(
        n2252) );
  AO221X1 U2455 ( .IN1(InstQueueRd_Addr[2]), .IN2(n2254), .IN3(n5180), .IN4(
        n2253), .IN5(n2252), .Q(n4304) );
  NAND2X0 U2456 ( .IN1(n5178), .IN2(n5207), .QN(n4465) );
  NAND2X0 U2457 ( .IN1(State[1]), .IN2(State[2]), .QN(n2255) );
  NAND3X0 U2458 ( .IN1(n5202), .IN2(n4465), .IN3(n2255), .QN(n4518) );
  NAND2X0 U2459 ( .IN1(n2256), .IN2(n2322), .QN(n4489) );
  INVX0 U2460 ( .INP(n4489), .ZN(n2315) );
  OA21X1 U2461 ( .IN1(n4518), .IN2(n2257), .IN3(n2315), .Q(n2267) );
  OA22X1 U2462 ( .IN1(n2267), .IN2(n2314), .IN3(n2266), .IN4(n2785), .Q(n2259)
         );
  NAND3X0 U2463 ( .IN1(n2259), .IN2(n2258), .IN3(n2783), .QN(n3016) );
  MUX21X1 U2464 ( .IN1(InstQueueRd_Addr[2]), .IN2(n4304), .S(n3016), .Q(n2281)
         );
  NAND3X0 U2465 ( .IN1(n4303), .IN2(n2260), .IN3(n2324), .QN(n2265) );
  NAND2X0 U2466 ( .IN1(InstQueueRd_Addr[2]), .IN2(InstQueueRd_Addr[1]), .QN(
        n2261) );
  NOR2X0 U2467 ( .IN1(InstQueueRd_Addr[3]), .IN2(n2261), .QN(n2399) );
  AO21X1 U2468 ( .IN1(InstQueueRd_Addr[3]), .IN2(n2261), .IN3(n2399), .Q(n2264) );
  OA221X1 U2469 ( .IN1(n4306), .IN2(InstQueueRd_Addr[3]), .IN3(n4303), .IN4(
        n2262), .IN5(n2323), .Q(n4271) );
  AO222X1 U2470 ( .IN1(n2923), .IN2(n2265), .IN3(n2276), .IN4(n2264), .IN5(
        n2263), .IN6(n4271), .Q(n4272) );
  MUX21X1 U2471 ( .IN1(InstQueueRd_Addr[3]), .IN2(n4272), .S(n3016), .Q(n2279)
         );
  OA21X1 U2472 ( .IN1(n2281), .IN2(n5200), .IN3(n2279), .Q(n2285) );
  NAND2X0 U2473 ( .IN1(n2783), .IN2(n2266), .QN(n2275) );
  INVX0 U2474 ( .INP(n2275), .ZN(n2270) );
  OA21X1 U2475 ( .IN1(READY_n), .IN2(n2267), .IN3(n2270), .Q(n2268) );
  AND3X1 U2476 ( .IN1(n4515), .IN2(n2269), .IN3(n2268), .Q(n2307) );
  OA21X1 U2477 ( .IN1(Flush), .IN2(More), .IN3(n2307), .Q(n2284) );
  NOR2X0 U2478 ( .IN1(N4186), .IN2(N4187), .QN(n4605) );
  INVX0 U2479 ( .INP(n3016), .ZN(n2274) );
  NOR2X0 U2480 ( .IN1(n3021), .IN2(n2270), .QN(n2273) );
  NAND2X0 U2481 ( .IN1(n2271), .IN2(n3020), .QN(n2272) );
  NOR2X0 U2482 ( .IN1(n2273), .IN2(n2272), .QN(n3018) );
  NOR2X0 U2483 ( .IN1(n2274), .IN2(n3018), .QN(n2278) );
  MUX21X1 U2484 ( .IN1(n2276), .IN2(n2275), .S(n5183), .Q(n4299) );
  OA22X1 U2485 ( .IN1(n2278), .IN2(n5182), .IN3(n5199), .IN4(n4299), .Q(n2277)
         );
  AO21X1 U2486 ( .IN1(n5182), .IN2(n2278), .IN3(n2277), .Q(n2282) );
  NAND2X0 U2487 ( .IN1(N4186), .IN2(N4187), .QN(n4426) );
  AO22X1 U2488 ( .IN1(n2279), .IN2(n4426), .IN3(n2281), .IN4(n5200), .Q(n2280)
         );
  AO222X1 U2489 ( .IN1(n4605), .IN2(n2282), .IN3(n4605), .IN4(n2281), .IN5(
        n2282), .IN6(n2280), .Q(n2283) );
  OR4X1 U2490 ( .IN1(n2286), .IN2(n2285), .IN3(n2284), .IN4(n2283), .Q(n2287)
         );
  NAND2X0 U2491 ( .IN1(n4445), .IN2(n2287), .QN(n2288) );
  NAND4X0 U2492 ( .IN1(n4450), .IN2(n3288), .IN3(n2311), .IN4(n2288), .QN(
        n2289) );
  NOR2X0 U2493 ( .IN1(n2310), .IN2(n2289), .QN(n2292) );
  AND2X1 U2494 ( .IN1(n4516), .IN2(n2292), .Q(n2294) );
  NAND2X0 U2495 ( .IN1(State2[1]), .IN2(n5179), .QN(n2290) );
  OA221X1 U2496 ( .IN1(n2290), .IN2(READY_n), .IN3(n2290), .IN4(n5176), .IN5(
        n4468), .Q(n2293) );
  NAND2X0 U2497 ( .IN1(n5203), .IN2(n4469), .QN(n3286) );
  NOR2X0 U2498 ( .IN1(n4518), .IN2(n3286), .QN(n2291) );
  NAND3X0 U2499 ( .IN1(n3027), .IN2(n2291), .IN3(n4486), .QN(n4446) );
  NAND3X0 U2500 ( .IN1(n2293), .IN2(n4446), .IN3(n2292), .QN(n4473) );
  INVX0 U2501 ( .INP(n4473), .ZN(n4474) );
  MUX21X1 U2502 ( .IN1(n2294), .IN2(n5176), .S(n4474), .Q(n2295) );
  NAND2X0 U2503 ( .IN1(n2296), .IN2(n2295), .QN(n2068) );
  AOI22X1 U2504 ( .IN1(n4319), .IN2(\C1/DATA2_16 ), .IN3(\C1/DATA1_16 ), .IN4(
        n4318), .QN(n2298) );
  NAND2X0 U2505 ( .IN1(n2298), .IN2(n2297), .QN(n1958) );
  NAND2X0 U2506 ( .IN1(n2300), .IN2(n2299), .QN(n2786) );
  INVX0 U2507 ( .INP(n2786), .ZN(n3301) );
  NOR2X0 U2508 ( .IN1(n2302), .IN2(n2301), .QN(n2828) );
  OAI221X1 U2509 ( .IN1(n2306), .IN2(n2305), .IN3(n2306), .IN4(n2304), .IN5(
        n2303), .QN(n2784) );
  AO22X1 U2510 ( .IN1(n3301), .IN2(n2785), .IN3(n2828), .IN4(n2784), .Q(n2308)
         );
  NOR2X0 U2511 ( .IN1(n2307), .IN2(n4519), .QN(n4491) );
  MUX21X1 U2512 ( .IN1(More), .IN2(n2308), .S(n4491), .Q(n2309) );
  NOR2X0 U2513 ( .IN1(n2310), .IN2(n2309), .QN(n2312) );
  NAND2X0 U2514 ( .IN1(n2312), .IN2(n2311), .QN(n2029) );
  OA22X1 U2515 ( .IN1(n2315), .IN2(n2314), .IN3(n2785), .IN4(n2313), .Q(n2321)
         );
  NAND2X0 U2516 ( .IN1(n2316), .IN2(n2941), .QN(n3025) );
  NAND4X0 U2517 ( .IN1(n2319), .IN2(n2318), .IN3(n2317), .IN4(n2955), .QN(
        n3024) );
  OR3X1 U2518 ( .IN1(n2320), .IN2(n3025), .IN3(n3024), .Q(n2335) );
  AO21X1 U2519 ( .IN1(n2321), .IN2(n2335), .IN3(n4519), .Q(n4321) );
  NOR2X0 U2520 ( .IN1(n2322), .IN2(n4321), .QN(n4322) );
  AOI22X1 U2521 ( .IN1(n4322), .IN2(Datai[30]), .IN3(EAX[30]), .IN4(n4321), 
        .QN(n2603) );
  NAND2X0 U2522 ( .IN1(\InstQueue[11][1] ), .IN2(n2588), .QN(n2334) );
  NOR2X0 U2523 ( .IN1(n2323), .IN2(n5177), .QN(n2397) );
  NOR2X0 U2524 ( .IN1(n5177), .IN2(n2324), .QN(n2398) );
  AO22X1 U2525 ( .IN1(\InstQueue[6][1] ), .IN2(n2397), .IN3(\InstQueue[14][1] ), .IN4(n2398), .Q(n2326) );
  AND2X1 U2526 ( .IN1(n2399), .IN2(\InstQueue[10][1] ), .Q(n2325) );
  NOR2X0 U2527 ( .IN1(n2326), .IN2(n2325), .QN(n2412) );
  AO22X1 U2528 ( .IN1(n2479), .IN2(\InstQueue[4][1] ), .IN3(n2478), .IN4(
        \InstQueue[12][1] ), .Q(n2328) );
  AO22X1 U2529 ( .IN1(n2480), .IN2(\DP_OP_469J1_133_8416/n117 ), .IN3(n2481), 
        .IN4(\InstQueue[8][1] ), .Q(n2327) );
  NOR2X0 U2530 ( .IN1(n2328), .IN2(n2327), .QN(n2472) );
  OA22X1 U2531 ( .IN1(N2884), .IN2(n2412), .IN3(n2472), .IN4(n2589), .Q(n2333)
         );
  NAND2X0 U2532 ( .IN1(\InstQueue[7][1] ), .IN2(n2592), .QN(n2332) );
  INVX0 U2533 ( .INP(n3020), .ZN(n2594) );
  AO22X1 U2534 ( .IN1(n2480), .IN2(\InstQueue[1][1] ), .IN3(n2481), .IN4(
        \InstQueue[9][1] ), .Q(n2330) );
  AO22X1 U2535 ( .IN1(n2479), .IN2(\InstQueue[5][1] ), .IN3(n2478), .IN4(
        \InstQueue[13][1] ), .Q(n2329) );
  OR2X1 U2536 ( .IN1(n2330), .IN2(n2329), .Q(n2413) );
  NAND2X0 U2537 ( .IN1(n2594), .IN2(n2413), .QN(n2331) );
  NAND4X0 U2538 ( .IN1(n2334), .IN2(n2333), .IN3(n2332), .IN4(n2331), .QN(
        n3028) );
  INVX0 U2539 ( .INP(n2335), .ZN(n4328) );
  AO222X1 U2540 ( .IN1(n3028), .IN2(n2600), .IN3(n4328), .IN4(EAX[24]), .IN5(
        n2599), .IN6(Datai[8]), .Q(n2629) );
  NAND2X0 U2541 ( .IN1(\InstQueue[11][0] ), .IN2(n2588), .QN(n2345) );
  AO22X1 U2542 ( .IN1(\InstQueue[6][0] ), .IN2(n2397), .IN3(\InstQueue[14][0] ), .IN4(n2398), .Q(n2337) );
  AND2X1 U2543 ( .IN1(n2399), .IN2(\InstQueue[10][0] ), .Q(n2336) );
  NOR2X0 U2544 ( .IN1(n2337), .IN2(n2336), .QN(n2418) );
  AO22X1 U2545 ( .IN1(n2479), .IN2(\InstQueue[4][0] ), .IN3(n2478), .IN4(
        \InstQueue[12][0] ), .Q(n2339) );
  AO22X1 U2546 ( .IN1(n2480), .IN2(\DP_OP_469J1_133_8416/n116 ), .IN3(n2481), 
        .IN4(\InstQueue[8][0] ), .Q(n2338) );
  NOR2X0 U2547 ( .IN1(n2339), .IN2(n2338), .QN(n2485) );
  OA22X1 U2548 ( .IN1(N2884), .IN2(n2418), .IN3(n2485), .IN4(n2589), .Q(n2344)
         );
  NAND2X0 U2549 ( .IN1(\InstQueue[7][0] ), .IN2(n2592), .QN(n2343) );
  AO22X1 U2550 ( .IN1(n2480), .IN2(\InstQueue[1][0] ), .IN3(n2481), .IN4(
        \InstQueue[9][0] ), .Q(n2341) );
  AO22X1 U2551 ( .IN1(n2479), .IN2(\InstQueue[5][0] ), .IN3(n2478), .IN4(
        \InstQueue[13][0] ), .Q(n2340) );
  OR2X1 U2552 ( .IN1(n2341), .IN2(n2340), .Q(n2419) );
  NAND2X0 U2553 ( .IN1(n2594), .IN2(n2419), .QN(n2342) );
  NAND4X0 U2554 ( .IN1(n2345), .IN2(n2344), .IN3(n2343), .IN4(n2342), .QN(
        n3029) );
  AO222X1 U2555 ( .IN1(n3029), .IN2(n2600), .IN3(n4328), .IN4(EAX[23]), .IN5(
        n2599), .IN6(Datai[7]), .Q(n2636) );
  AO22X1 U2556 ( .IN1(n2480), .IN2(\InstQueue[15][7] ), .IN3(n2481), .IN4(
        \InstQueue[7][7] ), .Q(n2347) );
  AO22X1 U2557 ( .IN1(n2479), .IN2(\InstQueue[3][7] ), .IN3(n2478), .IN4(
        \InstQueue[11][7] ), .Q(n2346) );
  OR2X1 U2558 ( .IN1(n2347), .IN2(n2346), .Q(n2492) );
  INVX0 U2559 ( .INP(n2492), .ZN(n2350) );
  AO22X1 U2560 ( .IN1(\InstQueue[6][7] ), .IN2(n2397), .IN3(\InstQueue[14][7] ), .IN4(n2398), .Q(n2349) );
  AND2X1 U2561 ( .IN1(n2399), .IN2(\InstQueue[10][7] ), .Q(n2348) );
  NOR2X0 U2562 ( .IN1(n2349), .IN2(n2348), .QN(n2591) );
  OA22X1 U2563 ( .IN1(n2350), .IN2(n2589), .IN3(n2591), .IN4(n5183), .Q(n2356)
         );
  INVX0 U2564 ( .INP(n3021), .ZN(n2493) );
  AO22X1 U2565 ( .IN1(n2480), .IN2(\InstQueue[1][7] ), .IN3(n2481), .IN4(
        \InstQueue[9][7] ), .Q(n2352) );
  AO22X1 U2566 ( .IN1(n2479), .IN2(\InstQueue[5][7] ), .IN3(n2478), .IN4(
        \InstQueue[13][7] ), .Q(n2351) );
  OR2X1 U2567 ( .IN1(n2352), .IN2(n2351), .Q(n2593) );
  AO22X1 U2568 ( .IN1(n2479), .IN2(\InstQueue[4][7] ), .IN3(n2478), .IN4(
        \InstQueue[12][7] ), .Q(n2354) );
  AO22X1 U2569 ( .IN1(n2480), .IN2(\DP_OP_469J1_133_8416/n123 ), .IN3(n2481), 
        .IN4(\InstQueue[8][7] ), .Q(n2353) );
  NOR2X0 U2570 ( .IN1(n2354), .IN2(n2353), .QN(n2590) );
  INVX0 U2571 ( .INP(n2590), .ZN(n2426) );
  AOI22X1 U2572 ( .IN1(n2493), .IN2(n2593), .IN3(n2594), .IN4(n2426), .QN(
        n2355) );
  NAND2X0 U2573 ( .IN1(n2356), .IN2(n2355), .QN(n3030) );
  AND2X1 U2574 ( .IN1(n3030), .IN2(n2600), .Q(n2635) );
  AO22X1 U2575 ( .IN1(n2599), .IN2(Datai[6]), .IN3(n4328), .IN4(EAX[22]), .Q(
        n2642) );
  AO22X1 U2576 ( .IN1(n2480), .IN2(\InstQueue[15][6] ), .IN3(n2481), .IN4(
        \InstQueue[7][6] ), .Q(n2358) );
  AO22X1 U2577 ( .IN1(n2479), .IN2(\InstQueue[3][6] ), .IN3(n2478), .IN4(
        \InstQueue[11][6] ), .Q(n2357) );
  NOR2X0 U2578 ( .IN1(n2358), .IN2(n2357), .QN(n2499) );
  AO22X1 U2579 ( .IN1(\InstQueue[14][6] ), .IN2(n2398), .IN3(\InstQueue[6][6] ), .IN4(n2397), .Q(n2360) );
  AND2X1 U2580 ( .IN1(n2399), .IN2(\InstQueue[10][6] ), .Q(n2359) );
  NOR2X0 U2581 ( .IN1(n2360), .IN2(n2359), .QN(n2582) );
  OA22X1 U2582 ( .IN1(n2499), .IN2(n2589), .IN3(n2582), .IN4(n5183), .Q(n2366)
         );
  AO22X1 U2583 ( .IN1(n2479), .IN2(\InstQueue[4][6] ), .IN3(n2478), .IN4(
        \InstQueue[12][6] ), .Q(n2362) );
  AO22X1 U2584 ( .IN1(n2480), .IN2(\DP_OP_469J1_133_8416/n122 ), .IN3(n2481), 
        .IN4(\InstQueue[8][6] ), .Q(n2361) );
  NOR2X0 U2585 ( .IN1(n2362), .IN2(n2361), .QN(n2581) );
  AO22X1 U2586 ( .IN1(n2480), .IN2(\InstQueue[1][6] ), .IN3(n2481), .IN4(
        \InstQueue[9][6] ), .Q(n2364) );
  AO22X1 U2587 ( .IN1(n2479), .IN2(\InstQueue[5][6] ), .IN3(n2478), .IN4(
        \InstQueue[13][6] ), .Q(n2363) );
  OR2X1 U2588 ( .IN1(n2364), .IN2(n2363), .Q(n2583) );
  INVX0 U2589 ( .INP(n2583), .ZN(n2434) );
  OA22X1 U2590 ( .IN1(n2581), .IN2(n3020), .IN3(n2434), .IN4(n3021), .Q(n2365)
         );
  NAND2X0 U2591 ( .IN1(n2366), .IN2(n2365), .QN(n3031) );
  AND2X1 U2592 ( .IN1(n3031), .IN2(n2600), .Q(n2641) );
  AO22X1 U2593 ( .IN1(n2599), .IN2(Datai[5]), .IN3(n4328), .IN4(EAX[21]), .Q(
        n2648) );
  AO22X1 U2594 ( .IN1(n2480), .IN2(\InstQueue[15][5] ), .IN3(n2481), .IN4(
        \InstQueue[7][5] ), .Q(n2368) );
  AO22X1 U2595 ( .IN1(n2479), .IN2(\InstQueue[3][5] ), .IN3(n2478), .IN4(
        \InstQueue[11][5] ), .Q(n2367) );
  NOR2X0 U2596 ( .IN1(n2368), .IN2(n2367), .QN(n2507) );
  AO22X1 U2597 ( .IN1(\InstQueue[14][5] ), .IN2(n2398), .IN3(\InstQueue[6][5] ), .IN4(n2397), .Q(n2370) );
  AND2X1 U2598 ( .IN1(n2399), .IN2(\InstQueue[10][5] ), .Q(n2369) );
  NOR2X0 U2599 ( .IN1(n2370), .IN2(n2369), .QN(n2575) );
  OA22X1 U2600 ( .IN1(n2507), .IN2(n2589), .IN3(n2575), .IN4(n5183), .Q(n2376)
         );
  AO22X1 U2601 ( .IN1(n2479), .IN2(\InstQueue[4][5] ), .IN3(n2478), .IN4(
        \InstQueue[12][5] ), .Q(n2372) );
  AO22X1 U2602 ( .IN1(n2480), .IN2(\DP_OP_469J1_133_8416/n121 ), .IN3(n2481), 
        .IN4(\InstQueue[8][5] ), .Q(n2371) );
  NOR2X0 U2603 ( .IN1(n2372), .IN2(n2371), .QN(n2574) );
  AO22X1 U2604 ( .IN1(n2480), .IN2(\InstQueue[1][5] ), .IN3(n2481), .IN4(
        \InstQueue[9][5] ), .Q(n2374) );
  AO22X1 U2605 ( .IN1(n2479), .IN2(\InstQueue[5][5] ), .IN3(n2478), .IN4(
        \InstQueue[13][5] ), .Q(n2373) );
  OR2X1 U2606 ( .IN1(n2374), .IN2(n2373), .Q(n2576) );
  INVX0 U2607 ( .INP(n2576), .ZN(n2442) );
  OA22X1 U2608 ( .IN1(n2574), .IN2(n3020), .IN3(n2442), .IN4(n3021), .Q(n2375)
         );
  NAND2X0 U2609 ( .IN1(n2376), .IN2(n2375), .QN(n3032) );
  AND2X1 U2610 ( .IN1(n3032), .IN2(n2600), .Q(n2647) );
  AO22X1 U2611 ( .IN1(n2599), .IN2(Datai[4]), .IN3(n4328), .IN4(EAX[20]), .Q(
        n2654) );
  AO22X1 U2612 ( .IN1(n2480), .IN2(\InstQueue[15][4] ), .IN3(n2481), .IN4(
        \InstQueue[7][4] ), .Q(n2378) );
  AO22X1 U2613 ( .IN1(n2479), .IN2(\InstQueue[3][4] ), .IN3(n2478), .IN4(
        \InstQueue[11][4] ), .Q(n2377) );
  NOR2X0 U2614 ( .IN1(n2378), .IN2(n2377), .QN(n2514) );
  AO22X1 U2615 ( .IN1(\InstQueue[6][4] ), .IN2(n2397), .IN3(\InstQueue[14][4] ), .IN4(n2398), .Q(n2380) );
  AND2X1 U2616 ( .IN1(n2399), .IN2(\InstQueue[10][4] ), .Q(n2379) );
  NOR2X0 U2617 ( .IN1(n2380), .IN2(n2379), .QN(n2568) );
  OA22X1 U2618 ( .IN1(n2514), .IN2(n2589), .IN3(n2568), .IN4(n5183), .Q(n2386)
         );
  AO22X1 U2619 ( .IN1(n2479), .IN2(\InstQueue[4][4] ), .IN3(n2478), .IN4(
        \InstQueue[12][4] ), .Q(n2382) );
  AO22X1 U2620 ( .IN1(n2480), .IN2(\DP_OP_469J1_133_8416/n120 ), .IN3(n2481), 
        .IN4(\InstQueue[8][4] ), .Q(n2381) );
  NOR2X0 U2621 ( .IN1(n2382), .IN2(n2381), .QN(n2567) );
  AO22X1 U2622 ( .IN1(n2480), .IN2(\InstQueue[1][4] ), .IN3(n2481), .IN4(
        \InstQueue[9][4] ), .Q(n2384) );
  AO22X1 U2623 ( .IN1(n2479), .IN2(\InstQueue[5][4] ), .IN3(n2478), .IN4(
        \InstQueue[13][4] ), .Q(n2383) );
  OR2X1 U2624 ( .IN1(n2384), .IN2(n2383), .Q(n2569) );
  INVX0 U2625 ( .INP(n2569), .ZN(n2450) );
  OA22X1 U2626 ( .IN1(n2567), .IN2(n3020), .IN3(n2450), .IN4(n3021), .Q(n2385)
         );
  NAND2X0 U2627 ( .IN1(n2386), .IN2(n2385), .QN(n3033) );
  AND2X1 U2628 ( .IN1(n3033), .IN2(n2600), .Q(n2653) );
  AO22X1 U2629 ( .IN1(n2599), .IN2(Datai[3]), .IN3(n4328), .IN4(EAX[19]), .Q(
        n2660) );
  AO22X1 U2630 ( .IN1(\InstQueue[15][3] ), .IN2(n2480), .IN3(n2481), .IN4(
        \InstQueue[7][3] ), .Q(n2388) );
  AO22X1 U2631 ( .IN1(n2479), .IN2(\InstQueue[3][3] ), .IN3(n2478), .IN4(
        \InstQueue[11][3] ), .Q(n2387) );
  NOR2X0 U2632 ( .IN1(n2388), .IN2(n2387), .QN(n2521) );
  AO22X1 U2633 ( .IN1(\InstQueue[6][3] ), .IN2(n2397), .IN3(\InstQueue[14][3] ), .IN4(n2398), .Q(n2390) );
  AND2X1 U2634 ( .IN1(n2399), .IN2(\InstQueue[10][3] ), .Q(n2389) );
  NOR2X0 U2635 ( .IN1(n2390), .IN2(n2389), .QN(n2561) );
  OA22X1 U2636 ( .IN1(n2521), .IN2(n2589), .IN3(n2561), .IN4(n5183), .Q(n2396)
         );
  AO22X1 U2637 ( .IN1(n2479), .IN2(\InstQueue[4][3] ), .IN3(n2478), .IN4(
        \InstQueue[12][3] ), .Q(n2392) );
  AO22X1 U2638 ( .IN1(n2480), .IN2(\DP_OP_469J1_133_8416/n119 ), .IN3(n2481), 
        .IN4(\InstQueue[8][3] ), .Q(n2391) );
  NOR2X0 U2639 ( .IN1(n2392), .IN2(n2391), .QN(n2560) );
  AO22X1 U2640 ( .IN1(n2480), .IN2(\InstQueue[1][3] ), .IN3(n2481), .IN4(
        \InstQueue[9][3] ), .Q(n2394) );
  AO22X1 U2641 ( .IN1(n2479), .IN2(\InstQueue[5][3] ), .IN3(n2478), .IN4(
        \InstQueue[13][3] ), .Q(n2393) );
  OR2X1 U2642 ( .IN1(n2394), .IN2(n2393), .Q(n2562) );
  INVX0 U2643 ( .INP(n2562), .ZN(n2458) );
  OA22X1 U2644 ( .IN1(n2560), .IN2(n3020), .IN3(n2458), .IN4(n3021), .Q(n2395)
         );
  NAND2X0 U2645 ( .IN1(n2396), .IN2(n2395), .QN(n3034) );
  AND2X1 U2646 ( .IN1(n3034), .IN2(n2600), .Q(n2659) );
  AO22X1 U2647 ( .IN1(n2599), .IN2(Datai[2]), .IN3(n4328), .IN4(EAX[18]), .Q(
        n2668) );
  AO22X1 U2648 ( .IN1(\InstQueue[14][2] ), .IN2(n2398), .IN3(\InstQueue[6][2] ), .IN4(n2397), .Q(n2401) );
  AND2X1 U2649 ( .IN1(n2399), .IN2(\InstQueue[10][2] ), .Q(n2400) );
  NOR2X0 U2650 ( .IN1(n2401), .IN2(n2400), .QN(n2554) );
  AO22X1 U2651 ( .IN1(n2480), .IN2(\InstQueue[15][2] ), .IN3(n2481), .IN4(
        \InstQueue[7][2] ), .Q(n2403) );
  AO22X1 U2652 ( .IN1(n2479), .IN2(\InstQueue[3][2] ), .IN3(n2478), .IN4(
        \InstQueue[11][2] ), .Q(n2402) );
  NOR2X0 U2653 ( .IN1(n2403), .IN2(n2402), .QN(n2528) );
  OA22X1 U2654 ( .IN1(n2554), .IN2(n5183), .IN3(n2528), .IN4(n2589), .Q(n2409)
         );
  AO22X1 U2655 ( .IN1(n2480), .IN2(\InstQueue[1][2] ), .IN3(n2481), .IN4(
        \InstQueue[9][2] ), .Q(n2405) );
  AO22X1 U2656 ( .IN1(n2479), .IN2(\InstQueue[5][2] ), .IN3(n2478), .IN4(
        \InstQueue[13][2] ), .Q(n2404) );
  OR2X1 U2657 ( .IN1(n2405), .IN2(n2404), .Q(n2555) );
  INVX0 U2658 ( .INP(n2555), .ZN(n2466) );
  AO22X1 U2659 ( .IN1(n2479), .IN2(\InstQueue[4][2] ), .IN3(n2478), .IN4(
        \InstQueue[12][2] ), .Q(n2407) );
  AO22X1 U2660 ( .IN1(n2480), .IN2(\DP_OP_469J1_133_8416/n118 ), .IN3(n2481), 
        .IN4(\InstQueue[8][2] ), .Q(n2406) );
  NOR2X0 U2661 ( .IN1(n2407), .IN2(n2406), .QN(n2553) );
  OA22X1 U2662 ( .IN1(n2466), .IN2(n3021), .IN3(n2553), .IN4(n3020), .Q(n2408)
         );
  NAND2X0 U2663 ( .IN1(n2409), .IN2(n2408), .QN(n3035) );
  AND2X1 U2664 ( .IN1(n3035), .IN2(n2600), .Q(n2667) );
  AO22X1 U2665 ( .IN1(n2599), .IN2(Datai[1]), .IN3(n4328), .IN4(EAX[17]), .Q(
        n2674) );
  AO22X1 U2666 ( .IN1(n2480), .IN2(\InstQueue[15][1] ), .IN3(n2481), .IN4(
        \InstQueue[7][1] ), .Q(n2411) );
  AO22X1 U2667 ( .IN1(n2479), .IN2(\InstQueue[3][1] ), .IN3(n2478), .IN4(
        \InstQueue[11][1] ), .Q(n2410) );
  NOR2X0 U2668 ( .IN1(n2411), .IN2(n2410), .QN(n2543) );
  OA22X1 U2669 ( .IN1(n2543), .IN2(n2589), .IN3(n2412), .IN4(n5183), .Q(n2415)
         );
  INVX0 U2670 ( .INP(n2413), .ZN(n2475) );
  OA22X1 U2671 ( .IN1(n2472), .IN2(n3020), .IN3(n2475), .IN4(n3021), .Q(n2414)
         );
  NAND2X0 U2672 ( .IN1(n2415), .IN2(n2414), .QN(n3036) );
  AND2X1 U2673 ( .IN1(n3036), .IN2(n2600), .Q(n2673) );
  AO22X1 U2674 ( .IN1(n2599), .IN2(Datai[0]), .IN3(n4328), .IN4(EAX[16]), .Q(
        n2680) );
  AO22X1 U2675 ( .IN1(n2480), .IN2(\InstQueue[15][0] ), .IN3(n2481), .IN4(
        \InstQueue[7][0] ), .Q(n2417) );
  AO22X1 U2676 ( .IN1(n2479), .IN2(\InstQueue[3][0] ), .IN3(n2478), .IN4(
        \InstQueue[11][0] ), .Q(n2416) );
  NOR2X0 U2677 ( .IN1(n2417), .IN2(n2416), .QN(n2535) );
  OA22X1 U2678 ( .IN1(n2418), .IN2(n5183), .IN3(n2535), .IN4(n2589), .Q(n2421)
         );
  INVX0 U2679 ( .INP(n2419), .ZN(n2488) );
  OA22X1 U2680 ( .IN1(n2488), .IN2(n3021), .IN3(n2485), .IN4(n3020), .Q(n2420)
         );
  NAND2X0 U2681 ( .IN1(n2421), .IN2(n2420), .QN(n3037) );
  AND2X1 U2682 ( .IN1(n3037), .IN2(n2600), .Q(n2679) );
  AND2X1 U2683 ( .IN1(n4328), .IN2(EAX[15]), .Q(n2686) );
  AOI22X1 U2684 ( .IN1(n2479), .IN2(\InstQueue[2][7] ), .IN3(n2478), .IN4(
        \InstQueue[10][7] ), .QN(n2424) );
  NAND2X0 U2685 ( .IN1(n2480), .IN2(\InstQueue[14][7] ), .QN(n2423) );
  NAND2X0 U2686 ( .IN1(n2481), .IN2(\InstQueue[6][7] ), .QN(n2422) );
  NAND4X0 U2687 ( .IN1(n2424), .IN2(n2423), .IN3(n2422), .IN4(n5177), .QN(
        n2425) );
  OA21X1 U2688 ( .IN1(n5177), .IN2(n2426), .IN3(n2425), .Q(n2491) );
  AO22X1 U2689 ( .IN1(n4306), .IN2(n2593), .IN3(n2594), .IN4(n2492), .Q(n2427)
         );
  AO21X1 U2690 ( .IN1(n2491), .IN2(n5183), .IN3(n2427), .Q(n3038) );
  AND2X1 U2691 ( .IN1(n2599), .IN2(Datai[15]), .Q(n2428) );
  AO21X1 U2692 ( .IN1(n3038), .IN2(n2600), .IN3(n2428), .Q(n2685) );
  AND2X1 U2693 ( .IN1(n4328), .IN2(EAX[14]), .Q(n2692) );
  AOI22X1 U2694 ( .IN1(n2479), .IN2(\InstQueue[2][6] ), .IN3(n2478), .IN4(
        \InstQueue[10][6] ), .QN(n2431) );
  NAND2X0 U2695 ( .IN1(n2480), .IN2(\InstQueue[14][6] ), .QN(n2430) );
  NAND2X0 U2696 ( .IN1(n2481), .IN2(\InstQueue[6][6] ), .QN(n2429) );
  NAND4X0 U2697 ( .IN1(n2431), .IN2(n2430), .IN3(n2429), .IN4(n5177), .QN(
        n2433) );
  NAND2X0 U2698 ( .IN1(InstQueueRd_Addr[1]), .IN2(n2581), .QN(n2432) );
  NAND2X0 U2699 ( .IN1(n2433), .IN2(n2432), .QN(n2501) );
  OA22X1 U2700 ( .IN1(n2499), .IN2(n3020), .IN3(n2434), .IN4(n4303), .Q(n2435)
         );
  OAI21X1 U2701 ( .IN1(N2884), .IN2(n2501), .IN3(n2435), .QN(n3039) );
  AND2X1 U2702 ( .IN1(n2599), .IN2(Datai[14]), .Q(n2436) );
  AO21X1 U2703 ( .IN1(n3039), .IN2(n2600), .IN3(n2436), .Q(n2691) );
  AND2X1 U2704 ( .IN1(n4328), .IN2(EAX[13]), .Q(n2698) );
  AOI22X1 U2705 ( .IN1(n2479), .IN2(\InstQueue[2][5] ), .IN3(n2478), .IN4(
        \InstQueue[10][5] ), .QN(n2439) );
  NAND2X0 U2706 ( .IN1(n2480), .IN2(\InstQueue[14][5] ), .QN(n2438) );
  NAND2X0 U2707 ( .IN1(n2481), .IN2(\InstQueue[6][5] ), .QN(n2437) );
  NAND4X0 U2708 ( .IN1(n2439), .IN2(n2438), .IN3(n2437), .IN4(n5177), .QN(
        n2441) );
  NAND2X0 U2709 ( .IN1(InstQueueRd_Addr[1]), .IN2(n2574), .QN(n2440) );
  NAND2X0 U2710 ( .IN1(n2441), .IN2(n2440), .QN(n2508) );
  OA22X1 U2711 ( .IN1(n2507), .IN2(n3020), .IN3(n2442), .IN4(n4303), .Q(n2443)
         );
  OAI21X1 U2712 ( .IN1(N2884), .IN2(n2508), .IN3(n2443), .QN(n3040) );
  AND2X1 U2713 ( .IN1(n2599), .IN2(Datai[13]), .Q(n2444) );
  AO21X1 U2714 ( .IN1(n3040), .IN2(n2600), .IN3(n2444), .Q(n2697) );
  AND2X1 U2715 ( .IN1(n4328), .IN2(EAX[12]), .Q(n2704) );
  AOI22X1 U2716 ( .IN1(n2479), .IN2(\InstQueue[2][4] ), .IN3(n2478), .IN4(
        \InstQueue[10][4] ), .QN(n2447) );
  NAND2X0 U2717 ( .IN1(n2480), .IN2(\InstQueue[14][4] ), .QN(n2446) );
  NAND2X0 U2718 ( .IN1(n2481), .IN2(\InstQueue[6][4] ), .QN(n2445) );
  NAND4X0 U2719 ( .IN1(n2447), .IN2(n2446), .IN3(n2445), .IN4(n5177), .QN(
        n2449) );
  NAND2X0 U2720 ( .IN1(InstQueueRd_Addr[1]), .IN2(n2567), .QN(n2448) );
  NAND2X0 U2721 ( .IN1(n2449), .IN2(n2448), .QN(n2515) );
  OA22X1 U2722 ( .IN1(n2514), .IN2(n3020), .IN3(n2450), .IN4(n4303), .Q(n2451)
         );
  OAI21X1 U2723 ( .IN1(N2884), .IN2(n2515), .IN3(n2451), .QN(n3041) );
  AND2X1 U2724 ( .IN1(n2599), .IN2(Datai[12]), .Q(n2452) );
  AO21X1 U2725 ( .IN1(n3041), .IN2(n2600), .IN3(n2452), .Q(n2703) );
  AND2X1 U2726 ( .IN1(n4328), .IN2(EAX[11]), .Q(n2710) );
  AOI22X1 U2727 ( .IN1(\InstQueue[2][3] ), .IN2(n2479), .IN3(n2478), .IN4(
        \InstQueue[10][3] ), .QN(n2455) );
  NAND2X0 U2728 ( .IN1(n2480), .IN2(\InstQueue[14][3] ), .QN(n2454) );
  NAND2X0 U2729 ( .IN1(n2481), .IN2(\InstQueue[6][3] ), .QN(n2453) );
  NAND4X0 U2730 ( .IN1(n2455), .IN2(n2454), .IN3(n2453), .IN4(n5177), .QN(
        n2457) );
  NAND2X0 U2731 ( .IN1(InstQueueRd_Addr[1]), .IN2(n2560), .QN(n2456) );
  NAND2X0 U2732 ( .IN1(n2457), .IN2(n2456), .QN(n2522) );
  OA22X1 U2733 ( .IN1(n2521), .IN2(n3020), .IN3(n2458), .IN4(n4303), .Q(n2459)
         );
  OAI21X1 U2734 ( .IN1(N2884), .IN2(n2522), .IN3(n2459), .QN(n3042) );
  AND2X1 U2735 ( .IN1(n2599), .IN2(Datai[11]), .Q(n2460) );
  AO21X1 U2736 ( .IN1(n3042), .IN2(n2600), .IN3(n2460), .Q(n2709) );
  AND2X1 U2737 ( .IN1(n4328), .IN2(EAX[10]), .Q(n2716) );
  AOI22X1 U2738 ( .IN1(n2479), .IN2(\InstQueue[2][2] ), .IN3(n2478), .IN4(
        \InstQueue[10][2] ), .QN(n2463) );
  NAND2X0 U2739 ( .IN1(n2480), .IN2(\InstQueue[14][2] ), .QN(n2462) );
  NAND2X0 U2740 ( .IN1(n2481), .IN2(\InstQueue[6][2] ), .QN(n2461) );
  NAND4X0 U2741 ( .IN1(n2463), .IN2(n2462), .IN3(n2461), .IN4(n5177), .QN(
        n2465) );
  NAND2X0 U2742 ( .IN1(InstQueueRd_Addr[1]), .IN2(n2553), .QN(n2464) );
  NAND2X0 U2743 ( .IN1(n2465), .IN2(n2464), .QN(n2529) );
  OA22X1 U2744 ( .IN1(n2466), .IN2(n4303), .IN3(n2528), .IN4(n3020), .Q(n2467)
         );
  OAI21X1 U2745 ( .IN1(N2884), .IN2(n2529), .IN3(n2467), .QN(n3043) );
  AND2X1 U2746 ( .IN1(n2599), .IN2(Datai[10]), .Q(n2468) );
  AO21X1 U2747 ( .IN1(n3043), .IN2(n2600), .IN3(n2468), .Q(n2715) );
  AND2X1 U2748 ( .IN1(n4328), .IN2(EAX[9]), .Q(n2722) );
  AOI22X1 U2749 ( .IN1(n2479), .IN2(\InstQueue[2][1] ), .IN3(n2478), .IN4(
        \InstQueue[10][1] ), .QN(n2471) );
  NAND2X0 U2750 ( .IN1(n2480), .IN2(\InstQueue[14][1] ), .QN(n2470) );
  NAND2X0 U2751 ( .IN1(n2481), .IN2(\InstQueue[6][1] ), .QN(n2469) );
  NAND4X0 U2752 ( .IN1(n2471), .IN2(n2470), .IN3(n2469), .IN4(n5177), .QN(
        n2474) );
  NAND2X0 U2753 ( .IN1(InstQueueRd_Addr[1]), .IN2(n2472), .QN(n2473) );
  NAND2X0 U2754 ( .IN1(n2474), .IN2(n2473), .QN(n2544) );
  OA22X1 U2755 ( .IN1(n2543), .IN2(n3020), .IN3(n2475), .IN4(n4303), .Q(n2476)
         );
  OAI21X1 U2756 ( .IN1(N2884), .IN2(n2544), .IN3(n2476), .QN(n3044) );
  AND2X1 U2757 ( .IN1(n2599), .IN2(Datai[9]), .Q(n2477) );
  AO21X1 U2758 ( .IN1(n3044), .IN2(n2600), .IN3(n2477), .Q(n2721) );
  AND2X1 U2759 ( .IN1(n4328), .IN2(EAX[8]), .Q(n2728) );
  AOI22X1 U2760 ( .IN1(n2479), .IN2(\InstQueue[2][0] ), .IN3(n2478), .IN4(
        \InstQueue[10][0] ), .QN(n2484) );
  NAND2X0 U2761 ( .IN1(n2480), .IN2(\InstQueue[14][0] ), .QN(n2483) );
  NAND2X0 U2762 ( .IN1(n2481), .IN2(\InstQueue[6][0] ), .QN(n2482) );
  NAND4X0 U2763 ( .IN1(n2484), .IN2(n2483), .IN3(n2482), .IN4(n5177), .QN(
        n2487) );
  NAND2X0 U2764 ( .IN1(InstQueueRd_Addr[1]), .IN2(n2485), .QN(n2486) );
  NAND2X0 U2765 ( .IN1(n2487), .IN2(n2486), .QN(n2536) );
  OA22X1 U2766 ( .IN1(n2488), .IN2(n4303), .IN3(n2535), .IN4(n3020), .Q(n2489)
         );
  OAI21X1 U2767 ( .IN1(N2884), .IN2(n2536), .IN3(n2489), .QN(n3045) );
  AND2X1 U2768 ( .IN1(n2599), .IN2(Datai[8]), .Q(n2490) );
  AO21X1 U2769 ( .IN1(n3045), .IN2(n2600), .IN3(n2490), .Q(n2727) );
  AND2X1 U2770 ( .IN1(n4328), .IN2(EAX[7]), .Q(n2734) );
  AO22X1 U2771 ( .IN1(n2500), .IN2(\InstQueue[9][7] ), .IN3(N2884), .IN4(n2491), .Q(n2496) );
  AO22X1 U2772 ( .IN1(n2498), .IN2(\InstQueue[5][7] ), .IN3(n2493), .IN4(n2492), .Q(n2495) );
  AO22X1 U2773 ( .IN1(n2546), .IN2(\InstQueue[13][7] ), .IN3(n2547), .IN4(
        \InstQueue[1][7] ), .Q(n2494) );
  NOR3X0 U2774 ( .IN1(n2496), .IN2(n2495), .IN3(n2494), .QN(n4132) );
  INVX0 U2775 ( .INP(n4132), .ZN(n3947) );
  AND2X1 U2776 ( .IN1(n2599), .IN2(Datai[7]), .Q(n2497) );
  AO21X1 U2777 ( .IN1(n3947), .IN2(n2600), .IN3(n2497), .Q(n2733) );
  AND2X1 U2778 ( .IN1(n4328), .IN2(EAX[6]), .Q(n2740) );
  INVX0 U2779 ( .INP(n2498), .ZN(n2542) );
  OA22X1 U2780 ( .IN1(n2499), .IN2(n3021), .IN3(n2542), .IN4(n5271), .Q(n2505)
         );
  INVX0 U2781 ( .INP(n2500), .ZN(n2545) );
  OA22X1 U2782 ( .IN1(n2545), .IN2(n5264), .IN3(n5183), .IN4(n2501), .Q(n2504)
         );
  NAND2X0 U2783 ( .IN1(n2546), .IN2(\InstQueue[13][6] ), .QN(n2503) );
  NAND2X0 U2784 ( .IN1(n2547), .IN2(\InstQueue[1][6] ), .QN(n2502) );
  NAND4X0 U2785 ( .IN1(n2505), .IN2(n2504), .IN3(n2503), .IN4(n2502), .QN(
        n2895) );
  AND2X1 U2786 ( .IN1(n2599), .IN2(Datai[6]), .Q(n2506) );
  AO21X1 U2787 ( .IN1(n2895), .IN2(n2600), .IN3(n2506), .Q(n2739) );
  AND2X1 U2788 ( .IN1(n4328), .IN2(EAX[5]), .Q(n2746) );
  OA22X1 U2789 ( .IN1(n2507), .IN2(n3021), .IN3(n2542), .IN4(n5272), .Q(n2512)
         );
  OA22X1 U2790 ( .IN1(n2545), .IN2(n5265), .IN3(n5183), .IN4(n2508), .Q(n2511)
         );
  NAND2X0 U2791 ( .IN1(n2546), .IN2(\InstQueue[13][5] ), .QN(n2510) );
  NAND2X0 U2792 ( .IN1(n2547), .IN2(\InstQueue[1][5] ), .QN(n2509) );
  NAND4X0 U2793 ( .IN1(n2512), .IN2(n2511), .IN3(n2510), .IN4(n2509), .QN(
        n2899) );
  AND2X1 U2794 ( .IN1(n2599), .IN2(Datai[5]), .Q(n2513) );
  AO21X1 U2795 ( .IN1(n2899), .IN2(n2600), .IN3(n2513), .Q(n2745) );
  AND2X1 U2796 ( .IN1(n4328), .IN2(EAX[4]), .Q(n2752) );
  OA22X1 U2797 ( .IN1(n2514), .IN2(n3021), .IN3(n2542), .IN4(n5273), .Q(n2519)
         );
  OA22X1 U2798 ( .IN1(n2545), .IN2(n5266), .IN3(n5183), .IN4(n2515), .Q(n2518)
         );
  NAND2X0 U2799 ( .IN1(n2546), .IN2(\InstQueue[13][4] ), .QN(n2517) );
  NAND2X0 U2800 ( .IN1(n2547), .IN2(\InstQueue[1][4] ), .QN(n2516) );
  NAND4X0 U2801 ( .IN1(n2519), .IN2(n2518), .IN3(n2517), .IN4(n2516), .QN(
        n4078) );
  AND2X1 U2802 ( .IN1(n2599), .IN2(Datai[4]), .Q(n2520) );
  AO21X1 U2803 ( .IN1(n4078), .IN2(n2600), .IN3(n2520), .Q(n2751) );
  AND2X1 U2804 ( .IN1(n4328), .IN2(EAX[3]), .Q(n2758) );
  OA22X1 U2805 ( .IN1(n2521), .IN2(n3021), .IN3(n2542), .IN4(n5270), .Q(n2526)
         );
  OA22X1 U2806 ( .IN1(n2545), .IN2(n5263), .IN3(n5183), .IN4(n2522), .Q(n2525)
         );
  NAND2X0 U2807 ( .IN1(n2546), .IN2(\InstQueue[13][3] ), .QN(n2524) );
  NAND2X0 U2808 ( .IN1(n2547), .IN2(\InstQueue[1][3] ), .QN(n2523) );
  NAND4X0 U2809 ( .IN1(n2526), .IN2(n2525), .IN3(n2524), .IN4(n2523), .QN(
        n2907) );
  AND2X1 U2810 ( .IN1(n2599), .IN2(Datai[3]), .Q(n2527) );
  AO21X1 U2811 ( .IN1(n2907), .IN2(n2600), .IN3(n2527), .Q(n2757) );
  AND2X1 U2812 ( .IN1(n4328), .IN2(EAX[2]), .Q(n2764) );
  OA22X1 U2813 ( .IN1(n2528), .IN2(n3021), .IN3(n2542), .IN4(n5274), .Q(n2533)
         );
  OA22X1 U2814 ( .IN1(n2545), .IN2(n5267), .IN3(n5183), .IN4(n2529), .Q(n2532)
         );
  NAND2X0 U2815 ( .IN1(n2546), .IN2(\InstQueue[13][2] ), .QN(n2531) );
  NAND2X0 U2816 ( .IN1(n2547), .IN2(\InstQueue[1][2] ), .QN(n2530) );
  NAND4X0 U2817 ( .IN1(n2533), .IN2(n2532), .IN3(n2531), .IN4(n2530), .QN(
        n2910) );
  AND2X1 U2818 ( .IN1(n2599), .IN2(Datai[2]), .Q(n2534) );
  AO21X1 U2819 ( .IN1(n2910), .IN2(n2600), .IN3(n2534), .Q(n2763) );
  AND2X1 U2820 ( .IN1(n4328), .IN2(EAX[1]), .Q(n2770) );
  OA22X1 U2821 ( .IN1(n2535), .IN2(n3021), .IN3(n2542), .IN4(n5276), .Q(n2540)
         );
  OA22X1 U2822 ( .IN1(n2545), .IN2(n5269), .IN3(n5183), .IN4(n2536), .Q(n2539)
         );
  NAND2X0 U2823 ( .IN1(n2546), .IN2(\InstQueue[13][0] ), .QN(n2538) );
  NAND2X0 U2824 ( .IN1(n2547), .IN2(\InstQueue[1][0] ), .QN(n2537) );
  NAND4X0 U2825 ( .IN1(n2540), .IN2(n2539), .IN3(n2538), .IN4(n2537), .QN(
        n4261) );
  AO21X1 U2826 ( .IN1(n2599), .IN2(Datai[0]), .IN3(n4328), .Q(n2541) );
  AO21X1 U2827 ( .IN1(n4261), .IN2(n2600), .IN3(n2541), .Q(n2775) );
  AND2X1 U2828 ( .IN1(n4328), .IN2(EAX[0]), .Q(n2774) );
  OA22X1 U2829 ( .IN1(n2543), .IN2(n3021), .IN3(n2542), .IN4(n5275), .Q(n2551)
         );
  OA22X1 U2830 ( .IN1(n2545), .IN2(n5268), .IN3(n5183), .IN4(n2544), .Q(n2550)
         );
  NAND2X0 U2831 ( .IN1(n2546), .IN2(\InstQueue[13][1] ), .QN(n2549) );
  NAND2X0 U2832 ( .IN1(n2547), .IN2(\InstQueue[1][1] ), .QN(n2548) );
  NAND4X0 U2833 ( .IN1(n2551), .IN2(n2550), .IN3(n2549), .IN4(n2548), .QN(
        n4223) );
  AND2X1 U2834 ( .IN1(n2599), .IN2(Datai[1]), .Q(n2552) );
  AO21X1 U2835 ( .IN1(n4223), .IN2(n2600), .IN3(n2552), .Q(n2768) );
  AND2X1 U2836 ( .IN1(n2629), .IN2(n2630), .Q(n2625) );
  NAND2X0 U2837 ( .IN1(\InstQueue[11][2] ), .IN2(n2588), .QN(n2559) );
  OA22X1 U2838 ( .IN1(N2884), .IN2(n2554), .IN3(n2553), .IN4(n2589), .Q(n2558)
         );
  NAND2X0 U2839 ( .IN1(\InstQueue[7][2] ), .IN2(n2592), .QN(n2557) );
  NAND2X0 U2840 ( .IN1(n2594), .IN2(n2555), .QN(n2556) );
  NAND4X0 U2841 ( .IN1(n2559), .IN2(n2558), .IN3(n2557), .IN4(n2556), .QN(
        n3046) );
  AO222X1 U2842 ( .IN1(n3046), .IN2(n2600), .IN3(n4328), .IN4(EAX[25]), .IN5(
        n2599), .IN6(Datai[9]), .Q(n2624) );
  NAND2X0 U2843 ( .IN1(\InstQueue[11][3] ), .IN2(n2588), .QN(n2566) );
  OA22X1 U2844 ( .IN1(N2884), .IN2(n2561), .IN3(n2560), .IN4(n2589), .Q(n2565)
         );
  NAND2X0 U2845 ( .IN1(\InstQueue[7][3] ), .IN2(n2592), .QN(n2564) );
  NAND2X0 U2846 ( .IN1(n2594), .IN2(n2562), .QN(n2563) );
  NAND4X0 U2847 ( .IN1(n2566), .IN2(n2565), .IN3(n2564), .IN4(n2563), .QN(
        n3047) );
  AO222X1 U2848 ( .IN1(n3047), .IN2(n2600), .IN3(n4328), .IN4(EAX[26]), .IN5(
        n2599), .IN6(Datai[10]), .Q(n2619) );
  NAND2X0 U2849 ( .IN1(\InstQueue[11][4] ), .IN2(n2588), .QN(n2573) );
  OA22X1 U2850 ( .IN1(N2884), .IN2(n2568), .IN3(n2567), .IN4(n2589), .Q(n2572)
         );
  NAND2X0 U2851 ( .IN1(\InstQueue[7][4] ), .IN2(n2592), .QN(n2571) );
  NAND2X0 U2852 ( .IN1(n2594), .IN2(n2569), .QN(n2570) );
  NAND4X0 U2853 ( .IN1(n2573), .IN2(n2572), .IN3(n2571), .IN4(n2570), .QN(
        n3048) );
  AO222X1 U2854 ( .IN1(n3048), .IN2(n2600), .IN3(n4328), .IN4(EAX[27]), .IN5(
        n2599), .IN6(Datai[11]), .Q(n2614) );
  NAND2X0 U2855 ( .IN1(\InstQueue[11][5] ), .IN2(n2588), .QN(n2580) );
  OA22X1 U2856 ( .IN1(N2884), .IN2(n2575), .IN3(n2574), .IN4(n2589), .Q(n2579)
         );
  NAND2X0 U2857 ( .IN1(\InstQueue[7][5] ), .IN2(n2592), .QN(n2578) );
  NAND2X0 U2858 ( .IN1(n2594), .IN2(n2576), .QN(n2577) );
  NAND4X0 U2859 ( .IN1(n2580), .IN2(n2579), .IN3(n2578), .IN4(n2577), .QN(
        n3049) );
  AO222X1 U2860 ( .IN1(n3049), .IN2(n2600), .IN3(n4328), .IN4(EAX[28]), .IN5(
        n2599), .IN6(Datai[12]), .Q(n2609) );
  NAND2X0 U2861 ( .IN1(\InstQueue[11][6] ), .IN2(n2588), .QN(n2587) );
  OA22X1 U2862 ( .IN1(N2884), .IN2(n2582), .IN3(n2581), .IN4(n2589), .Q(n2586)
         );
  NAND2X0 U2863 ( .IN1(\InstQueue[7][6] ), .IN2(n2592), .QN(n2585) );
  NAND2X0 U2864 ( .IN1(n2594), .IN2(n2583), .QN(n2584) );
  NAND4X0 U2865 ( .IN1(n2587), .IN2(n2586), .IN3(n2585), .IN4(n2584), .QN(
        n3050) );
  AO222X1 U2866 ( .IN1(n3050), .IN2(n2600), .IN3(n4328), .IN4(EAX[29]), .IN5(
        n2599), .IN6(Datai[13]), .Q(n2604) );
  NAND2X0 U2867 ( .IN1(\InstQueue[11][7] ), .IN2(n2588), .QN(n2598) );
  OA22X1 U2868 ( .IN1(N2884), .IN2(n2591), .IN3(n2590), .IN4(n2589), .Q(n2597)
         );
  NAND2X0 U2869 ( .IN1(\InstQueue[7][7] ), .IN2(n2592), .QN(n2596) );
  NAND2X0 U2870 ( .IN1(n2594), .IN2(n2593), .QN(n2595) );
  NAND4X0 U2871 ( .IN1(n2598), .IN2(n2597), .IN3(n2596), .IN4(n2595), .QN(
        n3051) );
  AO222X1 U2872 ( .IN1(n3051), .IN2(n2600), .IN3(n4328), .IN4(EAX[30]), .IN5(
        n2599), .IN6(Datai[14]), .Q(n4323) );
  INVX0 U2873 ( .INP(n4321), .ZN(n4327) );
  NAND2X0 U2874 ( .IN1(n2601), .IN2(n4327), .QN(n2602) );
  NAND2X0 U2875 ( .IN1(n2603), .IN2(n2602), .QN(n1960) );
  AOI22X1 U2876 ( .IN1(n4322), .IN2(Datai[29]), .IN3(EAX[29]), .IN4(n4321), 
        .QN(n2608) );
  HADDX1 U2877 ( .A0(n2605), .B0(n2604), .C1(n4324), .SO(n2606) );
  NAND2X0 U2878 ( .IN1(n2606), .IN2(n4327), .QN(n2607) );
  NAND2X0 U2879 ( .IN1(n2608), .IN2(n2607), .QN(n1961) );
  AOI22X1 U2880 ( .IN1(n4322), .IN2(Datai[28]), .IN3(EAX[28]), .IN4(n4321), 
        .QN(n2613) );
  HADDX1 U2881 ( .A0(n2610), .B0(n2609), .C1(n2605), .SO(n2611) );
  NAND2X0 U2882 ( .IN1(n2611), .IN2(n4327), .QN(n2612) );
  NAND2X0 U2883 ( .IN1(n2613), .IN2(n2612), .QN(n1962) );
  AOI22X1 U2884 ( .IN1(n4322), .IN2(Datai[27]), .IN3(EAX[27]), .IN4(n4321), 
        .QN(n2618) );
  HADDX1 U2885 ( .A0(n2615), .B0(n2614), .C1(n2610), .SO(n2616) );
  NAND2X0 U2886 ( .IN1(n2616), .IN2(n4327), .QN(n2617) );
  NAND2X0 U2887 ( .IN1(n2618), .IN2(n2617), .QN(n1963) );
  AOI22X1 U2888 ( .IN1(n4322), .IN2(Datai[26]), .IN3(EAX[26]), .IN4(n4321), 
        .QN(n2623) );
  HADDX1 U2889 ( .A0(n2620), .B0(n2619), .C1(n2615), .SO(n2621) );
  NAND2X0 U2890 ( .IN1(n2621), .IN2(n4327), .QN(n2622) );
  NAND2X0 U2891 ( .IN1(n2623), .IN2(n2622), .QN(n1964) );
  AOI22X1 U2892 ( .IN1(n4322), .IN2(Datai[25]), .IN3(EAX[25]), .IN4(n4321), 
        .QN(n2628) );
  HADDX1 U2893 ( .A0(n2625), .B0(n2624), .C1(n2620), .SO(n2626) );
  NAND2X0 U2894 ( .IN1(n2626), .IN2(n4327), .QN(n2627) );
  NAND2X0 U2895 ( .IN1(n2628), .IN2(n2627), .QN(n1965) );
  AOI22X1 U2896 ( .IN1(n4322), .IN2(Datai[24]), .IN3(EAX[24]), .IN4(n4321), 
        .QN(n2633) );
  XOR2X1 U2897 ( .IN1(n2630), .IN2(n2629), .Q(n2631) );
  NAND2X0 U2898 ( .IN1(n2631), .IN2(n4327), .QN(n2632) );
  NAND2X0 U2899 ( .IN1(n2633), .IN2(n2632), .QN(n1966) );
  AOI22X1 U2900 ( .IN1(n4322), .IN2(Datai[23]), .IN3(EAX[23]), .IN4(n4321), 
        .QN(n2639) );
  FADDX1 U2901 ( .A(n2636), .B(n2635), .CI(n2634), .CO(n2630), .S(n2637) );
  NAND2X0 U2902 ( .IN1(n2637), .IN2(n4327), .QN(n2638) );
  NAND2X0 U2903 ( .IN1(n2639), .IN2(n2638), .QN(n1967) );
  AOI22X1 U2904 ( .IN1(n4322), .IN2(Datai[22]), .IN3(EAX[22]), .IN4(n4321), 
        .QN(n2645) );
  FADDX1 U2905 ( .A(n2642), .B(n2641), .CI(n2640), .CO(n2634), .S(n2643) );
  NAND2X0 U2906 ( .IN1(n2643), .IN2(n4327), .QN(n2644) );
  NAND2X0 U2907 ( .IN1(n2645), .IN2(n2644), .QN(n1968) );
  AOI22X1 U2908 ( .IN1(n4322), .IN2(Datai[21]), .IN3(EAX[21]), .IN4(n4321), 
        .QN(n2651) );
  FADDX1 U2909 ( .A(n2648), .B(n2647), .CI(n2646), .CO(n2640), .S(n2649) );
  NAND2X0 U2910 ( .IN1(n2649), .IN2(n4327), .QN(n2650) );
  NAND2X0 U2911 ( .IN1(n2651), .IN2(n2650), .QN(n1969) );
  AOI22X1 U2912 ( .IN1(n4322), .IN2(Datai[20]), .IN3(EAX[20]), .IN4(n4321), 
        .QN(n2657) );
  FADDX1 U2913 ( .A(n2654), .B(n2653), .CI(n2652), .CO(n2646), .S(n2655) );
  NAND2X0 U2914 ( .IN1(n2655), .IN2(n4327), .QN(n2656) );
  NAND2X0 U2915 ( .IN1(n2657), .IN2(n2656), .QN(n1970) );
  AOI22X1 U2916 ( .IN1(n4322), .IN2(Datai[19]), .IN3(EAX[19]), .IN4(n4321), 
        .QN(n2663) );
  FADDX1 U2917 ( .A(n2660), .B(n2659), .CI(n2658), .CO(n2652), .S(n2661) );
  NAND2X0 U2918 ( .IN1(n2661), .IN2(n4327), .QN(n2662) );
  NAND2X0 U2919 ( .IN1(n2663), .IN2(n2662), .QN(n1971) );
  AOI22X1 U2920 ( .IN1(n4319), .IN2(\C1/DATA2_28 ), .IN3(n4318), .IN4(
        \C1/DATA1_28 ), .QN(n2665) );
  NAND2X0 U2921 ( .IN1(n2665), .IN2(n2664), .QN(n1946) );
  AOI22X1 U2922 ( .IN1(n4322), .IN2(Datai[18]), .IN3(EAX[18]), .IN4(n4321), 
        .QN(n2671) );
  FADDX1 U2923 ( .A(n2668), .B(n2667), .CI(n2666), .CO(n2658), .S(n2669) );
  NAND2X0 U2924 ( .IN1(n2669), .IN2(n4327), .QN(n2670) );
  NAND2X0 U2925 ( .IN1(n2671), .IN2(n2670), .QN(n1972) );
  AOI22X1 U2926 ( .IN1(n4322), .IN2(Datai[17]), .IN3(EAX[17]), .IN4(n4321), 
        .QN(n2677) );
  FADDX1 U2927 ( .A(n2674), .B(n2673), .CI(n2672), .CO(n2666), .S(n2675) );
  NAND2X0 U2928 ( .IN1(n2675), .IN2(n4327), .QN(n2676) );
  NAND2X0 U2929 ( .IN1(n2677), .IN2(n2676), .QN(n1973) );
  AOI22X1 U2930 ( .IN1(n4322), .IN2(Datai[16]), .IN3(EAX[16]), .IN4(n4321), 
        .QN(n2683) );
  FADDX1 U2931 ( .A(n2680), .B(n2679), .CI(n2678), .CO(n2672), .S(n2681) );
  NAND2X0 U2932 ( .IN1(n2681), .IN2(n4327), .QN(n2682) );
  NAND2X0 U2933 ( .IN1(n2683), .IN2(n2682), .QN(n1974) );
  AOI22X1 U2934 ( .IN1(n4322), .IN2(Datai[15]), .IN3(EAX[15]), .IN4(n4321), 
        .QN(n2689) );
  FADDX1 U2935 ( .A(n2686), .B(n2685), .CI(n2684), .CO(n2678), .S(n2687) );
  NAND2X0 U2936 ( .IN1(n2687), .IN2(n4327), .QN(n2688) );
  NAND2X0 U2937 ( .IN1(n2689), .IN2(n2688), .QN(n1975) );
  AOI22X1 U2938 ( .IN1(n4322), .IN2(Datai[14]), .IN3(EAX[14]), .IN4(n4321), 
        .QN(n2695) );
  FADDX1 U2939 ( .A(n2692), .B(n2691), .CI(n2690), .CO(n2684), .S(n2693) );
  NAND2X0 U2940 ( .IN1(n2693), .IN2(n4327), .QN(n2694) );
  NAND2X0 U2941 ( .IN1(n2695), .IN2(n2694), .QN(n1976) );
  AOI22X1 U2942 ( .IN1(n4322), .IN2(Datai[13]), .IN3(EAX[13]), .IN4(n4321), 
        .QN(n2701) );
  FADDX1 U2943 ( .A(n2698), .B(n2697), .CI(n2696), .CO(n2690), .S(n2699) );
  NAND2X0 U2944 ( .IN1(n2699), .IN2(n4327), .QN(n2700) );
  NAND2X0 U2945 ( .IN1(n2701), .IN2(n2700), .QN(n1977) );
  AOI22X1 U2946 ( .IN1(n4322), .IN2(Datai[12]), .IN3(EAX[12]), .IN4(n4321), 
        .QN(n2707) );
  FADDX1 U2947 ( .A(n2704), .B(n2703), .CI(n2702), .CO(n2696), .S(n2705) );
  NAND2X0 U2948 ( .IN1(n2705), .IN2(n4327), .QN(n2706) );
  NAND2X0 U2949 ( .IN1(n2707), .IN2(n2706), .QN(n1978) );
  AOI22X1 U2950 ( .IN1(n4322), .IN2(Datai[11]), .IN3(EAX[11]), .IN4(n4321), 
        .QN(n2713) );
  FADDX1 U2951 ( .A(n2710), .B(n2709), .CI(n2708), .CO(n2702), .S(n2711) );
  NAND2X0 U2952 ( .IN1(n2711), .IN2(n4327), .QN(n2712) );
  NAND2X0 U2953 ( .IN1(n2713), .IN2(n2712), .QN(n1979) );
  AOI22X1 U2954 ( .IN1(n4322), .IN2(Datai[10]), .IN3(EAX[10]), .IN4(n4321), 
        .QN(n2719) );
  FADDX1 U2955 ( .A(n2716), .B(n2715), .CI(n2714), .CO(n2708), .S(n2717) );
  NAND2X0 U2956 ( .IN1(n2717), .IN2(n4327), .QN(n2718) );
  NAND2X0 U2957 ( .IN1(n2719), .IN2(n2718), .QN(n1980) );
  AOI22X1 U2958 ( .IN1(n4322), .IN2(Datai[9]), .IN3(EAX[9]), .IN4(n4321), .QN(
        n2725) );
  FADDX1 U2959 ( .A(n2722), .B(n2721), .CI(n2720), .CO(n2714), .S(n2723) );
  NAND2X0 U2960 ( .IN1(n2723), .IN2(n4327), .QN(n2724) );
  NAND2X0 U2961 ( .IN1(n2725), .IN2(n2724), .QN(n1981) );
  AOI22X1 U2962 ( .IN1(n4322), .IN2(Datai[8]), .IN3(EAX[8]), .IN4(n4321), .QN(
        n2731) );
  FADDX1 U2963 ( .A(n2728), .B(n2727), .CI(n2726), .CO(n2720), .S(n2729) );
  NAND2X0 U2964 ( .IN1(n2729), .IN2(n4327), .QN(n2730) );
  NAND2X0 U2965 ( .IN1(n2731), .IN2(n2730), .QN(n1982) );
  AOI22X1 U2966 ( .IN1(n4322), .IN2(Datai[7]), .IN3(EAX[7]), .IN4(n4321), .QN(
        n2737) );
  FADDX1 U2967 ( .A(n2734), .B(n2733), .CI(n2732), .CO(n2726), .S(n2735) );
  NAND2X0 U2968 ( .IN1(n2735), .IN2(n4327), .QN(n2736) );
  NAND2X0 U2969 ( .IN1(n2737), .IN2(n2736), .QN(n1983) );
  AOI22X1 U2970 ( .IN1(n4322), .IN2(Datai[6]), .IN3(EAX[6]), .IN4(n4321), .QN(
        n2743) );
  FADDX1 U2971 ( .A(n2740), .B(n2739), .CI(n2738), .CO(n2732), .S(n2741) );
  NAND2X0 U2972 ( .IN1(n2741), .IN2(n4327), .QN(n2742) );
  NAND2X0 U2973 ( .IN1(n2743), .IN2(n2742), .QN(n1984) );
  AOI22X1 U2974 ( .IN1(n4322), .IN2(Datai[5]), .IN3(EAX[5]), .IN4(n4321), .QN(
        n2749) );
  FADDX1 U2975 ( .A(n2746), .B(n2745), .CI(n2744), .CO(n2738), .S(n2747) );
  NAND2X0 U2976 ( .IN1(n2747), .IN2(n4327), .QN(n2748) );
  NAND2X0 U2977 ( .IN1(n2749), .IN2(n2748), .QN(n1985) );
  AOI22X1 U2978 ( .IN1(n4322), .IN2(Datai[4]), .IN3(EAX[4]), .IN4(n4321), .QN(
        n2755) );
  FADDX1 U2979 ( .A(n2752), .B(n2751), .CI(n2750), .CO(n2744), .S(n2753) );
  NAND2X0 U2980 ( .IN1(n2753), .IN2(n4327), .QN(n2754) );
  NAND2X0 U2981 ( .IN1(n2755), .IN2(n2754), .QN(n1986) );
  AOI22X1 U2982 ( .IN1(n4322), .IN2(Datai[3]), .IN3(EAX[3]), .IN4(n4321), .QN(
        n2761) );
  FADDX1 U2983 ( .A(n2758), .B(n2757), .CI(n2756), .CO(n2750), .S(n2759) );
  NAND2X0 U2984 ( .IN1(n2759), .IN2(n4327), .QN(n2760) );
  NAND2X0 U2985 ( .IN1(n2761), .IN2(n2760), .QN(n1987) );
  AOI22X1 U2986 ( .IN1(n4322), .IN2(Datai[2]), .IN3(EAX[2]), .IN4(n4321), .QN(
        n2767) );
  FADDX1 U2987 ( .A(n2764), .B(n2763), .CI(n2762), .CO(n2756), .S(n2765) );
  NAND2X0 U2988 ( .IN1(n2765), .IN2(n4327), .QN(n2766) );
  NAND2X0 U2989 ( .IN1(n2767), .IN2(n2766), .QN(n1988) );
  AOI22X1 U2990 ( .IN1(n4322), .IN2(Datai[1]), .IN3(EAX[1]), .IN4(n4321), .QN(
        n2773) );
  FADDX1 U2991 ( .A(n2770), .B(n2769), .CI(n2768), .CO(n2762), .S(n2771) );
  NAND2X0 U2992 ( .IN1(n2771), .IN2(n4327), .QN(n2772) );
  NAND2X0 U2993 ( .IN1(n2773), .IN2(n2772), .QN(n1989) );
  AOI22X1 U2994 ( .IN1(n4322), .IN2(Datai[0]), .IN3(EAX[0]), .IN4(n4321), .QN(
        n2778) );
  HADDX1 U2995 ( .A0(n2775), .B0(n2774), .C1(n2769), .SO(n2776) );
  NAND2X0 U2996 ( .IN1(n2776), .IN2(n4327), .QN(n2777) );
  NAND2X0 U2997 ( .IN1(n2778), .IN2(n2777), .QN(n1990) );
  NOR2X0 U2998 ( .IN1(n5203), .IN2(n5101), .QN(n5098) );
  NOR3X0 U2999 ( .IN1(READY_n), .IN2(n5242), .IN3(n4468), .QN(n2779) );
  NOR2X0 U3000 ( .IN1(n5098), .IN2(n2779), .QN(n2782) );
  NAND3X0 U3001 ( .IN1(State2[1]), .IN2(State2[0]), .IN3(n4473), .QN(n2780) );
  NAND2X0 U3002 ( .IN1(State2[2]), .IN2(n2780), .QN(n2781) );
  NAND2X0 U3003 ( .IN1(n2782), .IN2(n2781), .QN(n2066) );
  NOR2X0 U3004 ( .IN1(n4519), .IN2(n2783), .QN(n4236) );
  INVX0 U3005 ( .INP(n4236), .ZN(n4205) );
  NAND3X0 U3006 ( .IN1(InstAddrPointer[2]), .IN2(N1868), .IN3(
        InstAddrPointer[1]), .QN(n4061) );
  INVX0 U3007 ( .INP(n4061), .ZN(n4189) );
  NAND3X0 U3008 ( .IN1(InstAddrPointer[3]), .IN2(InstAddrPointer[4]), .IN3(
        n4189), .QN(n4180) );
  NOR2X0 U3009 ( .IN1(n5205), .IN2(n4180), .QN(n4174) );
  NAND2X0 U3010 ( .IN1(InstAddrPointer[6]), .IN2(n4174), .QN(n4154) );
  NOR2X0 U3011 ( .IN1(n5209), .IN2(n4154), .QN(n4017) );
  NAND2X0 U3012 ( .IN1(InstAddrPointer[8]), .IN2(n4017), .QN(n3976) );
  NOR2X0 U3013 ( .IN1(n5218), .IN2(n3976), .QN(n3966) );
  NAND2X0 U3014 ( .IN1(InstAddrPointer[10]), .IN2(n3966), .QN(n3913) );
  NOR2X0 U3015 ( .IN1(n5219), .IN2(n3913), .QN(n3903) );
  NAND2X0 U3016 ( .IN1(InstAddrPointer[12]), .IN2(n3903), .QN(n3851) );
  NOR2X0 U3017 ( .IN1(n5220), .IN2(n3851), .QN(n3841) );
  NAND2X0 U3018 ( .IN1(InstAddrPointer[14]), .IN2(n3841), .QN(n3789) );
  NOR2X0 U3019 ( .IN1(n5221), .IN2(n3789), .QN(n3779) );
  NAND2X0 U3020 ( .IN1(InstAddrPointer[16]), .IN2(n3779), .QN(n3730) );
  NOR2X0 U3021 ( .IN1(n5234), .IN2(n3730), .QN(n3723) );
  NAND2X0 U3022 ( .IN1(InstAddrPointer[18]), .IN2(n3723), .QN(n3665) );
  NOR2X0 U3023 ( .IN1(n5235), .IN2(n3665), .QN(n3560) );
  NAND2X0 U3024 ( .IN1(InstAddrPointer[20]), .IN2(n3560), .QN(n3566) );
  NOR2X0 U3025 ( .IN1(n5210), .IN2(n3566), .QN(n3583) );
  NAND2X0 U3026 ( .IN1(InstAddrPointer[22]), .IN2(n3583), .QN(n3591) );
  NOR2X0 U3027 ( .IN1(n5211), .IN2(n3591), .QN(n3608) );
  NAND2X0 U3028 ( .IN1(InstAddrPointer[24]), .IN2(n3608), .QN(n3616) );
  NOR2X0 U3029 ( .IN1(n5212), .IN2(n3616), .QN(n3633) );
  NAND2X0 U3030 ( .IN1(InstAddrPointer[26]), .IN2(n3633), .QN(n3641) );
  NOR2X0 U3031 ( .IN1(n5213), .IN2(n3641), .QN(n3658) );
  NAND2X0 U3032 ( .IN1(InstAddrPointer[28]), .IN2(n3658), .QN(n2922) );
  NOR2X0 U3033 ( .IN1(n4205), .IN2(n2922), .QN(n3327) );
  INVX0 U3034 ( .INP(n3327), .ZN(n2827) );
  INVX0 U3035 ( .INP(n2828), .ZN(n3295) );
  OA22X1 U3036 ( .IN1(n2786), .IN2(n2785), .IN3(n3295), .IN4(n2784), .Q(n3293)
         );
  INVX0 U3037 ( .INP(n3293), .ZN(n4492) );
  OA21X1 U3038 ( .IN1(n4492), .IN2(n3016), .IN3(n4445), .Q(n2924) );
  NAND2X0 U3039 ( .IN1(n3301), .IN2(n2924), .QN(n4208) );
  NOR2X0 U3040 ( .IN1(n5204), .IN2(n5185), .QN(n2800) );
  NOR2X0 U3041 ( .IN1(InstAddrPointer[2]), .IN2(n2800), .QN(n2802) );
  NOR2X0 U3042 ( .IN1(n2802), .IN2(n5222), .QN(n2806) );
  NAND2X0 U3043 ( .IN1(n2806), .IN2(InstAddrPointer[4]), .QN(n2805) );
  NOR2X0 U3044 ( .IN1(n2805), .IN2(n5205), .QN(n2797) );
  NAND2X0 U3045 ( .IN1(n2797), .IN2(InstAddrPointer[6]), .QN(n2796) );
  NOR2X0 U3046 ( .IN1(n2796), .IN2(n5209), .QN(n2815) );
  NAND2X0 U3047 ( .IN1(n2815), .IN2(InstAddrPointer[8]), .QN(n2816) );
  NOR2X0 U3048 ( .IN1(n2816), .IN2(n5218), .QN(n2795) );
  NAND2X0 U3049 ( .IN1(n2795), .IN2(InstAddrPointer[10]), .QN(n2817) );
  NOR2X0 U3050 ( .IN1(n2817), .IN2(n5219), .QN(n2794) );
  NAND2X0 U3051 ( .IN1(n2794), .IN2(InstAddrPointer[12]), .QN(n2818) );
  NOR2X0 U3052 ( .IN1(n2818), .IN2(n5220), .QN(n2793) );
  NAND2X0 U3053 ( .IN1(n2793), .IN2(InstAddrPointer[14]), .QN(n2819) );
  NOR2X0 U3054 ( .IN1(n2819), .IN2(n5221), .QN(n2792) );
  NAND2X0 U3055 ( .IN1(n2792), .IN2(InstAddrPointer[16]), .QN(n2820) );
  NOR2X0 U3056 ( .IN1(n2820), .IN2(n5234), .QN(n2791) );
  NAND2X0 U3057 ( .IN1(n2791), .IN2(InstAddrPointer[18]), .QN(n2821) );
  NOR2X0 U3058 ( .IN1(n2821), .IN2(n5235), .QN(n2790) );
  NAND2X0 U3059 ( .IN1(n2790), .IN2(InstAddrPointer[20]), .QN(n2822) );
  NOR2X0 U3060 ( .IN1(n2822), .IN2(n5210), .QN(n2789) );
  NAND2X0 U3061 ( .IN1(n2789), .IN2(InstAddrPointer[22]), .QN(n2823) );
  NOR2X0 U3062 ( .IN1(n2823), .IN2(n5211), .QN(n2788) );
  NAND2X0 U3063 ( .IN1(n2788), .IN2(InstAddrPointer[24]), .QN(n2824) );
  NOR2X0 U3064 ( .IN1(n2824), .IN2(n5212), .QN(n2787) );
  NAND2X0 U3065 ( .IN1(n2787), .IN2(InstAddrPointer[26]), .QN(n2825) );
  NOR2X0 U3066 ( .IN1(n2825), .IN2(n5213), .QN(n2826) );
  MUX21X1 U3067 ( .IN1(n5237), .IN2(InstAddrPointer[28]), .S(n2826), .Q(n3652)
         );
  MUX21X1 U3068 ( .IN1(n5233), .IN2(InstAddrPointer[26]), .S(n2787), .Q(n3627)
         );
  MUX21X1 U3069 ( .IN1(n5232), .IN2(InstAddrPointer[24]), .S(n2788), .Q(n3602)
         );
  MUX21X1 U3070 ( .IN1(n5231), .IN2(InstAddrPointer[22]), .S(n2789), .Q(n3577)
         );
  MUX21X1 U3071 ( .IN1(n5215), .IN2(InstAddrPointer[20]), .S(n2790), .Q(n3557)
         );
  XNOR2X1 U3072 ( .IN1(n2791), .IN2(InstAddrPointer[18]), .Q(n3722) );
  MUX21X1 U3073 ( .IN1(n5226), .IN2(InstAddrPointer[16]), .S(n2792), .Q(n3778)
         );
  MUX21X1 U3074 ( .IN1(n5227), .IN2(InstAddrPointer[14]), .S(n2793), .Q(n3840)
         );
  MUX21X1 U3075 ( .IN1(n5228), .IN2(InstAddrPointer[12]), .S(n2794), .Q(n3902)
         );
  MUX21X1 U3076 ( .IN1(n5229), .IN2(InstAddrPointer[10]), .S(n2795), .Q(n3965)
         );
  AO21X1 U3077 ( .IN1(n2796), .IN2(n5209), .IN3(n2815), .Q(n4155) );
  INVX0 U3078 ( .INP(n2895), .ZN(n4117) );
  OAI21X1 U3079 ( .IN1(n2797), .IN2(InstAddrPointer[6]), .IN3(n2796), .QN(
        n4179) );
  INVX0 U3080 ( .INP(n2899), .ZN(n4099) );
  AO21X1 U3081 ( .IN1(n2805), .IN2(n5205), .IN3(n2797), .Q(n4166) );
  INVX0 U3082 ( .INP(n2802), .ZN(n2799) );
  INVX0 U3083 ( .INP(n2806), .ZN(n2798) );
  OA21X1 U3084 ( .IN1(InstAddrPointer[3]), .IN2(n2799), .IN3(n2798), .Q(n4070)
         );
  INVX0 U3085 ( .INP(n2910), .ZN(n4030) );
  NAND2X0 U3086 ( .IN1(n5204), .IN2(n4261), .QN(n4260) );
  AO21X1 U3087 ( .IN1(n5204), .IN2(n5185), .IN3(n2800), .Q(n4238) );
  INVX0 U3088 ( .INP(n4223), .ZN(n2912) );
  OA21X1 U3089 ( .IN1(n4238), .IN2(n4260), .IN3(n2912), .Q(n2801) );
  AO21X1 U3090 ( .IN1(n4260), .IN2(n4238), .IN3(n2801), .Q(n4029) );
  NOR2X0 U3091 ( .IN1(n2802), .IN2(n4189), .QN(n4204) );
  INVX0 U3092 ( .INP(n2907), .ZN(n4044) );
  NOR2X0 U3093 ( .IN1(n4045), .IN2(n4044), .QN(n2804) );
  INVX0 U3094 ( .INP(n4045), .ZN(n2803) );
  OA22X1 U3095 ( .IN1(n4070), .IN2(n2804), .IN3(n2907), .IN4(n2803), .Q(n4079)
         );
  OAI21X1 U3096 ( .IN1(n2806), .IN2(InstAddrPointer[4]), .IN3(n2805), .QN(
        n4198) );
  INVX0 U3097 ( .INP(n4078), .ZN(n2901) );
  NOR2X0 U3098 ( .IN1(n4198), .IN2(n2901), .QN(n2808) );
  INVX0 U3099 ( .INP(n4198), .ZN(n2807) );
  OAI22X1 U3100 ( .IN1(n4079), .IN2(n2808), .IN3(n4078), .IN4(n2807), .QN(
        n4098) );
  INVX0 U3101 ( .INP(n4166), .ZN(n2809) );
  NAND2X0 U3102 ( .IN1(n2809), .IN2(n2899), .QN(n2810) );
  AO22X1 U3103 ( .IN1(n4099), .IN2(n4166), .IN3(n4098), .IN4(n2810), .Q(n4116)
         );
  INVX0 U3104 ( .INP(n4179), .ZN(n2811) );
  NAND2X0 U3105 ( .IN1(n2811), .IN2(n2895), .QN(n2812) );
  AO22X1 U3106 ( .IN1(n4117), .IN2(n4179), .IN3(n4116), .IN4(n2812), .Q(n4131)
         );
  INVX0 U3107 ( .INP(n4155), .ZN(n2813) );
  NAND2X0 U3108 ( .IN1(n3947), .IN2(n2813), .QN(n2814) );
  AO22X1 U3109 ( .IN1(n4155), .IN2(n4132), .IN3(n4131), .IN4(n2814), .Q(n3990)
         );
  MUX21X1 U3110 ( .IN1(n5225), .IN2(InstAddrPointer[8]), .S(n2815), .Q(n4010)
         );
  NOR2X0 U3111 ( .IN1(n3990), .IN2(n4010), .QN(n3989) );
  MUX21X1 U3112 ( .IN1(n5218), .IN2(InstAddrPointer[9]), .S(n2816), .Q(n3979)
         );
  NAND2X0 U3113 ( .IN1(n3989), .IN2(n3979), .QN(n3944) );
  NOR2X0 U3114 ( .IN1(n3965), .IN2(n3944), .QN(n3943) );
  MUX21X1 U3115 ( .IN1(n5219), .IN2(InstAddrPointer[11]), .S(n2817), .Q(n3916)
         );
  NAND2X0 U3116 ( .IN1(n3943), .IN2(n3916), .QN(n3882) );
  NOR2X0 U3117 ( .IN1(n3902), .IN2(n3882), .QN(n3881) );
  MUX21X1 U3118 ( .IN1(n5220), .IN2(InstAddrPointer[13]), .S(n2818), .Q(n3854)
         );
  NAND2X0 U3119 ( .IN1(n3881), .IN2(n3854), .QN(n3820) );
  NOR2X0 U3120 ( .IN1(n3840), .IN2(n3820), .QN(n3819) );
  MUX21X1 U3121 ( .IN1(n5221), .IN2(InstAddrPointer[15]), .S(n2819), .Q(n3792)
         );
  NAND2X0 U3122 ( .IN1(n3819), .IN2(n3792), .QN(n3760) );
  NOR2X0 U3123 ( .IN1(n3778), .IN2(n3760), .QN(n3759) );
  XNOR2X1 U3124 ( .IN1(n2820), .IN2(InstAddrPointer[17]), .Q(n3736) );
  NAND2X0 U3125 ( .IN1(n3759), .IN2(n3736), .QN(n3697) );
  NOR2X0 U3126 ( .IN1(n3722), .IN2(n3697), .QN(n3696) );
  XNOR2X1 U3127 ( .IN1(n2821), .IN2(InstAddrPointer[19]), .Q(n3677) );
  NAND2X0 U3128 ( .IN1(n3696), .IN2(n3677), .QN(n3535) );
  NOR2X0 U3129 ( .IN1(n3557), .IN2(n3535), .QN(n3534) );
  MUX21X1 U3130 ( .IN1(n5210), .IN2(InstAddrPointer[21]), .S(n2822), .Q(n3567)
         );
  NAND2X0 U3131 ( .IN1(n3534), .IN2(n3567), .QN(n3500) );
  NOR2X0 U3132 ( .IN1(n3577), .IN2(n3500), .QN(n3499) );
  MUX21X1 U3133 ( .IN1(n5211), .IN2(InstAddrPointer[23]), .S(n2823), .Q(n3592)
         );
  NAND2X0 U3134 ( .IN1(n3499), .IN2(n3592), .QN(n3464) );
  NOR2X0 U3135 ( .IN1(n3602), .IN2(n3464), .QN(n3463) );
  MUX21X1 U3136 ( .IN1(n5212), .IN2(InstAddrPointer[25]), .S(n2824), .Q(n3617)
         );
  NAND2X0 U3137 ( .IN1(n3463), .IN2(n3617), .QN(n3428) );
  NOR2X0 U3138 ( .IN1(n3627), .IN2(n3428), .QN(n3427) );
  MUX21X1 U3139 ( .IN1(n5213), .IN2(InstAddrPointer[27]), .S(n2825), .Q(n3642)
         );
  NAND2X0 U3140 ( .IN1(n3427), .IN2(n3642), .QN(n3392) );
  NOR2X0 U3141 ( .IN1(n3652), .IN2(n3392), .QN(n3391) );
  NAND2X0 U3142 ( .IN1(n2826), .IN2(InstAddrPointer[28]), .QN(n3302) );
  MUX21X1 U3143 ( .IN1(n5223), .IN2(InstAddrPointer[29]), .S(n3302), .Q(n2925)
         );
  NAND2X0 U3144 ( .IN1(n3391), .IN2(n2925), .QN(n3303) );
  OAI21X1 U3145 ( .IN1(n3391), .IN2(n2925), .IN3(n3303), .QN(n3357) );
  OA22X1 U3146 ( .IN1(InstAddrPointer[29]), .IN2(n2827), .IN3(n4208), .IN4(
        n3357), .Q(n2932) );
  NAND2X0 U3147 ( .IN1(n2828), .IN2(n2924), .QN(n4060) );
  INVX1 U3148 ( .INP(n4132), .ZN(n3993) );
  AO22X1 U3149 ( .IN1(n4132), .IN2(n2927), .IN3(n2829), .IN4(n2916), .Q(n3300)
         );
  HADDX1 U3150 ( .A0(n2830), .B0(InstAddrPointer[28]), .C1(n3296), .SO(n3654)
         );
  HADDX1 U3151 ( .A0(n2831), .B0(InstAddrPointer[28]), .C1(n3297), .SO(n2832)
         );
  AO22X1 U3152 ( .IN1(n4132), .IN2(n3654), .IN3(n2832), .IN4(n2916), .Q(n3394)
         );
  HADDX1 U3153 ( .A0(n2833), .B0(InstAddrPointer[27]), .C1(n2830), .SO(n3646)
         );
  HADDX1 U3154 ( .A0(n2834), .B0(InstAddrPointer[27]), .C1(n2831), .SO(n2835)
         );
  AO22X1 U3155 ( .IN1(n4132), .IN2(n3646), .IN3(n2835), .IN4(n2916), .Q(n3381)
         );
  HADDX1 U3156 ( .A0(n2836), .B0(InstAddrPointer[26]), .C1(n2833), .SO(n3629)
         );
  HADDX1 U3157 ( .A0(n2837), .B0(InstAddrPointer[26]), .C1(n2834), .SO(n2838)
         );
  AO22X1 U3158 ( .IN1(n4132), .IN2(n3629), .IN3(n2838), .IN4(n2916), .Q(n3430)
         );
  HADDX1 U3159 ( .A0(n2839), .B0(InstAddrPointer[25]), .C1(n2836), .SO(n3621)
         );
  HADDX1 U3160 ( .A0(n2840), .B0(InstAddrPointer[25]), .C1(n2837), .SO(n2841)
         );
  AO22X1 U3161 ( .IN1(n4132), .IN2(n3621), .IN3(n2841), .IN4(n2916), .Q(n3417)
         );
  HADDX1 U3162 ( .A0(n2842), .B0(InstAddrPointer[24]), .C1(n2839), .SO(n3604)
         );
  HADDX1 U3163 ( .A0(n2843), .B0(InstAddrPointer[24]), .C1(n2840), .SO(n2844)
         );
  AO22X1 U3164 ( .IN1(n4132), .IN2(n3604), .IN3(n2844), .IN4(n2916), .Q(n3466)
         );
  HADDX1 U3165 ( .A0(n2845), .B0(InstAddrPointer[23]), .C1(n2842), .SO(n3596)
         );
  HADDX1 U3166 ( .A0(n2846), .B0(InstAddrPointer[23]), .C1(n2843), .SO(n2847)
         );
  INVX0 U3167 ( .INP(n4132), .ZN(n2916) );
  AO22X1 U3168 ( .IN1(n4132), .IN2(n3596), .IN3(n2847), .IN4(n2916), .Q(n3453)
         );
  HADDX1 U3169 ( .A0(n2848), .B0(InstAddrPointer[22]), .C1(n2845), .SO(n3579)
         );
  HADDX1 U3170 ( .A0(n2849), .B0(InstAddrPointer[22]), .C1(n2846), .SO(n2850)
         );
  AO22X1 U3171 ( .IN1(n4132), .IN2(n3579), .IN3(n2850), .IN4(n2916), .Q(n3502)
         );
  HADDX1 U3172 ( .A0(n2851), .B0(InstAddrPointer[21]), .C1(n2848), .SO(n3571)
         );
  HADDX1 U3173 ( .A0(n2852), .B0(InstAddrPointer[21]), .C1(n2849), .SO(n2853)
         );
  AO22X1 U3174 ( .IN1(n4132), .IN2(n3571), .IN3(n2853), .IN4(n2916), .Q(n3489)
         );
  HADDX1 U3175 ( .A0(n2854), .B0(InstAddrPointer[20]), .C1(n2851), .SO(n3559)
         );
  HADDX1 U3176 ( .A0(n2855), .B0(InstAddrPointer[20]), .C1(n2852), .SO(n2856)
         );
  AO22X1 U3177 ( .IN1(n4132), .IN2(n3559), .IN3(n2856), .IN4(n2916), .Q(n3537)
         );
  HADDX1 U3178 ( .A0(n2857), .B0(InstAddrPointer[19]), .C1(n2854), .SO(n3668)
         );
  HADDX1 U3179 ( .A0(n2858), .B0(InstAddrPointer[19]), .C1(n2855), .SO(n2859)
         );
  AO22X1 U3180 ( .IN1(n4132), .IN2(n3668), .IN3(n2859), .IN4(n2916), .Q(n3527)
         );
  HADDX1 U3181 ( .A0(n2860), .B0(InstAddrPointer[18]), .C1(n2857), .SO(n3715)
         );
  HADDX1 U3182 ( .A0(n2861), .B0(InstAddrPointer[18]), .C1(n2858), .SO(n2862)
         );
  AO22X1 U3183 ( .IN1(n4132), .IN2(n3715), .IN3(n2862), .IN4(n2916), .Q(n3699)
         );
  HADDX1 U3184 ( .A0(n2863), .B0(InstAddrPointer[17]), .C1(n2860), .SO(n3735)
         );
  HADDX1 U3185 ( .A0(n2864), .B0(InstAddrPointer[17]), .C1(n2861), .SO(n2865)
         );
  AO22X1 U3186 ( .IN1(n4132), .IN2(n3735), .IN3(n2865), .IN4(n2916), .Q(n3688)
         );
  HADDX1 U3187 ( .A0(n2866), .B0(InstAddrPointer[16]), .C1(n2863), .SO(n3780)
         );
  HADDX1 U3188 ( .A0(n2867), .B0(InstAddrPointer[16]), .C1(n2864), .SO(n2868)
         );
  AO22X1 U3189 ( .IN1(n4132), .IN2(n3780), .IN3(n2868), .IN4(n2916), .Q(n3762)
         );
  HADDX1 U3190 ( .A0(n2869), .B0(InstAddrPointer[15]), .C1(n2866), .SO(n3794)
         );
  HADDX1 U3191 ( .A0(n2870), .B0(InstAddrPointer[15]), .C1(n2867), .SO(n2871)
         );
  AO22X1 U3192 ( .IN1(n4132), .IN2(n3794), .IN3(n2871), .IN4(n2916), .Q(n3751)
         );
  HADDX1 U3193 ( .A0(n2872), .B0(InstAddrPointer[14]), .C1(n2869), .SO(n3842)
         );
  HADDX1 U3194 ( .A0(n2873), .B0(InstAddrPointer[14]), .C1(n2870), .SO(n2874)
         );
  AO22X1 U3195 ( .IN1(n4132), .IN2(n3842), .IN3(n2874), .IN4(n2916), .Q(n3822)
         );
  HADDX1 U3196 ( .A0(n2875), .B0(InstAddrPointer[13]), .C1(n2872), .SO(n3856)
         );
  HADDX1 U3197 ( .A0(n2876), .B0(InstAddrPointer[13]), .C1(n2873), .SO(n2877)
         );
  AO22X1 U3198 ( .IN1(n4132), .IN2(n3856), .IN3(n2877), .IN4(n2916), .Q(n3812)
         );
  HADDX1 U3199 ( .A0(n2878), .B0(InstAddrPointer[12]), .C1(n2875), .SO(n3904)
         );
  HADDX1 U3200 ( .A0(n2879), .B0(InstAddrPointer[12]), .C1(n2876), .SO(n2880)
         );
  AO22X1 U3201 ( .IN1(n4132), .IN2(n3904), .IN3(n2880), .IN4(n2916), .Q(n3884)
         );
  HADDX1 U3202 ( .A0(n2881), .B0(InstAddrPointer[11]), .C1(n2878), .SO(n3918)
         );
  HADDX1 U3203 ( .A0(n2882), .B0(InstAddrPointer[11]), .C1(n2879), .SO(n2883)
         );
  AO22X1 U3204 ( .IN1(n4132), .IN2(n3918), .IN3(n2883), .IN4(n2916), .Q(n3874)
         );
  HADDX1 U3205 ( .A0(n2884), .B0(InstAddrPointer[10]), .C1(n2881), .SO(n3967)
         );
  HADDX1 U3206 ( .A0(n2885), .B0(InstAddrPointer[10]), .C1(n2882), .SO(n2886)
         );
  AO22X1 U3207 ( .IN1(n4132), .IN2(n3967), .IN3(n2886), .IN4(n2916), .Q(n3946)
         );
  HADDX1 U3208 ( .A0(n2887), .B0(InstAddrPointer[9]), .C1(n2884), .SO(n3981)
         );
  HADDX1 U3209 ( .A0(n2888), .B0(InstAddrPointer[9]), .C1(n2885), .SO(n2889)
         );
  AO22X1 U3210 ( .IN1(n4132), .IN2(n3981), .IN3(n2889), .IN4(n2916), .Q(n3936)
         );
  HADDX1 U3211 ( .A0(n2890), .B0(InstAddrPointer[8]), .C1(n2887), .SO(n4012)
         );
  HADDX1 U3212 ( .A0(n2891), .B0(InstAddrPointer[8]), .C1(n2888), .SO(n2892)
         );
  AO22X1 U3213 ( .IN1(n4132), .IN2(n4012), .IN3(n2892), .IN4(n2916), .Q(n3992)
         );
  NOR2X0 U3214 ( .IN1(n4117), .IN2(n3947), .QN(n4120) );
  HADDX1 U3215 ( .A0(n2893), .B0(InstAddrPointer[6]), .C1(n2918), .SO(n4175)
         );
  FADDX1 U3216 ( .A(InstAddrPointer[6]), .B(n2895), .CI(n2894), .CO(n2919), 
        .S(n2896) );
  AO22X1 U3217 ( .IN1(n4132), .IN2(n4175), .IN3(n2896), .IN4(n2916), .Q(n4119)
         );
  NOR2X0 U3218 ( .IN1(n4099), .IN2(n3947), .QN(n4102) );
  HADDX1 U3219 ( .A0(n2897), .B0(InstAddrPointer[5]), .C1(n2893), .SO(n4167)
         );
  FADDX1 U3220 ( .A(InstAddrPointer[5]), .B(n2899), .CI(n2898), .CO(n2894), 
        .S(n2900) );
  AO22X1 U3221 ( .IN1(n4132), .IN2(n4167), .IN3(n2900), .IN4(n2916), .Q(n4101)
         );
  NOR2X0 U3222 ( .IN1(n2901), .IN2(n3947), .QN(n4082) );
  HADDX1 U3223 ( .A0(n2902), .B0(InstAddrPointer[4]), .C1(n2897), .SO(n4190)
         );
  FADDX1 U3224 ( .A(InstAddrPointer[4]), .B(n4078), .CI(n2903), .CO(n2898), 
        .S(n2904) );
  AO22X1 U3225 ( .IN1(n4132), .IN2(n4190), .IN3(n2904), .IN4(n2916), .Q(n4081)
         );
  NOR2X0 U3226 ( .IN1(n4044), .IN2(n3947), .QN(n4041) );
  HADDX1 U3227 ( .A0(n2905), .B0(InstAddrPointer[3]), .C1(n2902), .SO(n4064)
         );
  FADDX1 U3228 ( .A(InstAddrPointer[3]), .B(n2907), .CI(n2906), .CO(n2903), 
        .S(n2908) );
  AO22X1 U3229 ( .IN1(n4132), .IN2(n4064), .IN3(n2908), .IN4(n2916), .Q(n4040)
         );
  NOR2X0 U3230 ( .IN1(n4030), .IN2(n3947), .QN(n4033) );
  HADDX1 U3231 ( .A0(InstAddrPointer[1]), .B0(InstAddrPointer[2]), .C1(n2905), 
        .SO(n4211) );
  FADDX1 U3232 ( .A(InstAddrPointer[2]), .B(n2910), .CI(n2909), .CO(n2906), 
        .S(n2911) );
  AO22X1 U3233 ( .IN1(n4132), .IN2(n4211), .IN3(n2911), .IN4(n2916), .Q(n4032)
         );
  NAND2X0 U3234 ( .IN1(n4132), .IN2(n2912), .QN(n4220) );
  HADDX1 U3235 ( .A0(n4261), .B0(N1868), .C1(n2915), .SO(n2913) );
  AO22X1 U3236 ( .IN1(N1868), .IN2(n4132), .IN3(n2913), .IN4(n2916), .Q(n4265)
         );
  INVX0 U3237 ( .INP(n4261), .ZN(n2914) );
  NOR2X0 U3238 ( .IN1(n2914), .IN2(n3947), .QN(n4264) );
  FADDX1 U3239 ( .A(InstAddrPointer[1]), .B(n4223), .CI(n2915), .CO(n2909), 
        .S(n2917) );
  AO22X1 U3240 ( .IN1(n4132), .IN2(n5185), .IN3(n2917), .IN4(n2916), .Q(n4218)
         );
  HADDX1 U3241 ( .A0(n2918), .B0(InstAddrPointer[7]), .C1(n2890), .SO(n4156)
         );
  FADDX1 U3242 ( .A(InstAddrPointer[7]), .B(n3993), .CI(n2919), .CO(n2891), 
        .S(n2920) );
  AO22X1 U3243 ( .IN1(n4132), .IN2(n4156), .IN3(n2920), .IN4(n2916), .Q(n4134)
         );
  AND2X1 U3244 ( .IN1(n4133), .IN2(n4134), .Q(n3991) );
  INVX0 U3245 ( .INP(n2921), .ZN(n3356) );
  NOR2X0 U3246 ( .IN1(n2924), .IN2(n4104), .QN(n4217) );
  AOI21X1 U3247 ( .IN1(n2922), .IN2(n4236), .IN3(n4217), .QN(n3328) );
  OA22X1 U3248 ( .IN1(n4060), .IN2(n3356), .IN3(n3328), .IN4(n5223), .Q(n2930)
         );
  NAND2X0 U3249 ( .IN1(n2924), .IN2(n2923), .QN(n4206) );
  INVX0 U3250 ( .INP(n4206), .ZN(n4237) );
  NAND2X0 U3251 ( .IN1(n2925), .IN2(n4237), .QN(n2929) );
  INVX0 U3252 ( .INP(n4217), .ZN(n4294) );
  AO22X1 U3253 ( .IN1(n4445), .IN2(n2926), .IN3(n4294), .IN4(n3178), .Q(n4290)
         );
  NAND2X0 U3254 ( .IN1(n4290), .IN2(n2927), .QN(n2928) );
  NAND2X0 U3255 ( .IN1(n4104), .IN2(rEIP[29]), .QN(n3363) );
  AND4X1 U3256 ( .IN1(n2930), .IN2(n2929), .IN3(n2928), .IN4(n3363), .Q(n2931)
         );
  NAND2X0 U3257 ( .IN1(n2932), .IN2(n2931), .QN(n1992) );
  NOR3X0 U3258 ( .IN1(rEIP[0]), .IN2(DataWidth[1]), .IN3(DataWidth[0]), .QN(
        n2935) );
  NAND2X0 U3259 ( .IN1(DataWidth[1]), .IN2(DataWidth[0]), .QN(n5174) );
  INVX0 U3260 ( .INP(n5174), .ZN(n5175) );
  NOR2X0 U3261 ( .IN1(n5175), .IN2(n5190), .QN(n5173) );
  NOR2X0 U3262 ( .IN1(n2935), .IN2(n5173), .QN(n2934) );
  NAND2X0 U3263 ( .IN1(n5175), .IN2(ByteEnable[1]), .QN(n2933) );
  NAND2X0 U3264 ( .IN1(n2934), .IN2(n2933), .QN(n1661) );
  NOR2X0 U3265 ( .IN1(N4154), .IN2(DataWidth[1]), .QN(n5171) );
  NOR2X0 U3266 ( .IN1(n2935), .IN2(n5171), .QN(n2937) );
  NAND2X0 U3267 ( .IN1(n5175), .IN2(ByteEnable[3]), .QN(n2936) );
  NAND2X0 U3268 ( .IN1(n2937), .IN2(n2936), .QN(n1663) );
  NOR2X0 U3269 ( .IN1(n5198), .IN2(n5182), .QN(n4504) );
  NAND2X0 U3270 ( .IN1(N4186), .IN2(n4504), .QN(n4480) );
  NOR2X0 U3271 ( .IN1(N1351), .IN2(n4480), .QN(n5097) );
  NOR2X0 U3272 ( .IN1(n5199), .IN2(N4188), .QN(n4848) );
  INVX0 U3273 ( .INP(n4848), .ZN(n2938) );
  NOR2X0 U3274 ( .IN1(n4426), .IN2(n2938), .QN(n5106) );
  NOR2X0 U3275 ( .IN1(n5097), .IN2(n5106), .QN(n4430) );
  INVX0 U3276 ( .INP(n5098), .ZN(n5020) );
  NOR2X0 U3277 ( .IN1(n5199), .IN2(n5182), .QN(n4604) );
  INVX0 U3278 ( .INP(n4604), .ZN(n2939) );
  NOR2X0 U3279 ( .IN1(n2939), .IN2(n4426), .QN(n5095) );
  INVX0 U3280 ( .INP(n5095), .ZN(n4566) );
  INVX0 U3281 ( .INP(n5096), .ZN(n4973) );
  NOR2X0 U3282 ( .IN1(N1351), .IN2(N4188), .QN(n4807) );
  NAND2X0 U3283 ( .IN1(n4605), .IN2(n4807), .QN(n4608) );
  NOR3X0 U3284 ( .IN1(State2[0]), .IN2(n5179), .IN3(n2940), .QN(n5016) );
  INVX0 U3285 ( .INP(n5016), .ZN(n4485) );
  NAND2X0 U3286 ( .IN1(n4485), .IN2(n4973), .QN(n5094) );
  INVX0 U3287 ( .INP(n5094), .ZN(n4972) );
  OA222X1 U3288 ( .IN1(n5020), .IN2(n4430), .IN3(n4566), .IN4(n4973), .IN5(
        n4608), .IN6(n4972), .Q(n3011) );
  INVX0 U3289 ( .INP(n3011), .ZN(n2999) );
  AND3X1 U3290 ( .IN1(n4430), .IN2(n4977), .IN3(n2999), .Q(n3010) );
  NAND2X0 U3291 ( .IN1(Datai[7]), .IN2(n3010), .QN(n2954) );
  NAND2X0 U3292 ( .IN1(n4977), .IN2(n5203), .QN(n4470) );
  AND2X1 U3293 ( .IN1(n4479), .IN2(n4470), .Q(n4431) );
  INVX0 U3294 ( .INP(n2941), .ZN(n2942) );
  AOI22X1 U3295 ( .IN1(n4255), .IN2(Datai[7]), .IN3(n2942), .IN4(n5016), .QN(
        n5156) );
  INVX0 U3296 ( .INP(Datai[29]), .ZN(n2965) );
  INVX0 U3297 ( .INP(Datai[27]), .ZN(n2981) );
  INVX0 U3298 ( .INP(Datai[25]), .ZN(n2997) );
  OR4X1 U3299 ( .IN1(Datai[19]), .IN2(Datai[20]), .IN3(Datai[21]), .IN4(
        Datai[22]), .Q(n2949) );
  OR4X1 U3300 ( .IN1(Datai[16]), .IN2(Datai[17]), .IN3(Datai[18]), .IN4(
        Datai[23]), .Q(n2948) );
  NOR4X0 U3301 ( .IN1(Datai[0]), .IN2(Datai[1]), .IN3(Datai[2]), .IN4(Datai[3]), .QN(n2946) );
  NOR4X0 U3302 ( .IN1(Datai[4]), .IN2(Datai[5]), .IN3(Datai[6]), .IN4(Datai[7]), .QN(n2945) );
  NOR4X0 U3303 ( .IN1(Datai[8]), .IN2(Datai[9]), .IN3(Datai[10]), .IN4(
        Datai[11]), .QN(n2944) );
  NOR4X0 U3304 ( .IN1(Datai[12]), .IN2(Datai[13]), .IN3(Datai[14]), .IN4(
        Datai[15]), .QN(n2943) );
  NAND4X0 U3305 ( .IN1(n2946), .IN2(n2945), .IN3(n2944), .IN4(n2943), .QN(
        n2947) );
  AND2X1 U3306 ( .IN1(Datai[31]), .IN2(n2947), .Q(n3005) );
  AO221X1 U3307 ( .IN1(Datai[31]), .IN2(n2949), .IN3(Datai[31]), .IN4(n2948), 
        .IN5(n3005), .Q(n3008) );
  NAND2X0 U3308 ( .IN1(Datai[24]), .IN2(n3008), .QN(n3007) );
  NOR2X0 U3309 ( .IN1(n2997), .IN2(n3007), .QN(n2996) );
  NAND2X0 U3310 ( .IN1(Datai[26]), .IN2(n2996), .QN(n2988) );
  NOR2X0 U3311 ( .IN1(n2981), .IN2(n2988), .QN(n2980) );
  NAND2X0 U3312 ( .IN1(Datai[28]), .IN2(n2980), .QN(n2972) );
  NOR2X0 U3313 ( .IN1(n2965), .IN2(n2972), .QN(n2964) );
  NAND2X0 U3314 ( .IN1(Datai[30]), .IN2(n2964), .QN(n2956) );
  NAND2X0 U3315 ( .IN1(Datai[31]), .IN2(n2956), .QN(n5155) );
  NAND2X0 U3316 ( .IN1(n5106), .IN2(n2999), .QN(n3009) );
  OA22X1 U3317 ( .IN1(n5156), .IN2(n3011), .IN3(n5155), .IN4(n3009), .Q(n2953)
         );
  INVX0 U3318 ( .INP(Datai[23]), .ZN(n2950) );
  INVX0 U3319 ( .INP(Datai[21]), .ZN(n2963) );
  INVX0 U3320 ( .INP(Datai[19]), .ZN(n2982) );
  INVX0 U3321 ( .INP(Datai[17]), .ZN(n2995) );
  NAND2X0 U3322 ( .IN1(Datai[16]), .IN2(n3005), .QN(n3004) );
  NOR2X0 U3323 ( .IN1(n2995), .IN2(n3004), .QN(n2994) );
  NAND2X0 U3324 ( .IN1(Datai[18]), .IN2(n2994), .QN(n2989) );
  NOR2X0 U3325 ( .IN1(n2982), .IN2(n2989), .QN(n2974) );
  NAND2X0 U3326 ( .IN1(Datai[20]), .IN2(n2974), .QN(n2973) );
  NOR2X0 U3327 ( .IN1(n2963), .IN2(n2973), .QN(n2962) );
  NAND2X0 U3328 ( .IN1(Datai[22]), .IN2(n2962), .QN(n2957) );
  MUX21X1 U3329 ( .IN1(n2950), .IN2(Datai[23]), .S(n2957), .Q(n5158) );
  NAND2X0 U3330 ( .IN1(n5098), .IN2(n5097), .QN(n4556) );
  INVX0 U3331 ( .INP(n4556), .ZN(n3006) );
  NAND2X0 U3332 ( .IN1(n5158), .IN2(n3006), .QN(n2952) );
  NAND2X0 U3333 ( .IN1(n3011), .IN2(\DP_OP_469J1_133_8416/n123 ), .QN(n2951)
         );
  NAND4X0 U3334 ( .IN1(n2954), .IN2(n2953), .IN3(n2952), .IN4(n2951), .QN(
        n1889) );
  NAND2X0 U3335 ( .IN1(Datai[6]), .IN2(n3010), .QN(n2961) );
  AOI22X1 U3336 ( .IN1(n4255), .IN2(Datai[6]), .IN3(n2955), .IN4(n5016), .QN(
        n5148) );
  OAI21X1 U3337 ( .IN1(Datai[30]), .IN2(n2964), .IN3(n2956), .QN(n5147) );
  OA22X1 U3338 ( .IN1(n3011), .IN2(n5148), .IN3(n5147), .IN4(n3009), .Q(n2960)
         );
  OA21X1 U3339 ( .IN1(Datai[22]), .IN2(n2962), .IN3(n2957), .Q(n5149) );
  NAND2X0 U3340 ( .IN1(n3006), .IN2(n5149), .QN(n2959) );
  NAND2X0 U3341 ( .IN1(n3011), .IN2(\DP_OP_469J1_133_8416/n122 ), .QN(n2958)
         );
  NAND4X0 U3342 ( .IN1(n2961), .IN2(n2960), .IN3(n2959), .IN4(n2958), .QN(
        n1890) );
  NAND2X0 U3343 ( .IN1(Datai[5]), .IN2(n3010), .QN(n2970) );
  AO21X1 U3344 ( .IN1(n2963), .IN2(n2973), .IN3(n2962), .Q(n5042) );
  AO21X1 U3345 ( .IN1(n2965), .IN2(n2972), .IN3(n2964), .Q(n5140) );
  OA22X1 U3346 ( .IN1(n4556), .IN2(n5042), .IN3(n3009), .IN4(n5140), .Q(n2969)
         );
  AO22X1 U3347 ( .IN1(Datai[5]), .IN2(n4255), .IN3(n5016), .IN4(n2966), .Q(
        n5041) );
  NAND2X0 U3348 ( .IN1(n2999), .IN2(n5041), .QN(n2968) );
  NAND2X0 U3349 ( .IN1(n3011), .IN2(\DP_OP_469J1_133_8416/n121 ), .QN(n2967)
         );
  NAND4X0 U3350 ( .IN1(n2970), .IN2(n2969), .IN3(n2968), .IN4(n2967), .QN(
        n1891) );
  NAND2X0 U3351 ( .IN1(Datai[4]), .IN2(n3010), .QN(n2978) );
  AOI22X1 U3352 ( .IN1(n4255), .IN2(Datai[4]), .IN3(n2971), .IN4(n5016), .QN(
        n5134) );
  OAI21X1 U3353 ( .IN1(Datai[28]), .IN2(n2980), .IN3(n2972), .QN(n5133) );
  OA22X1 U3354 ( .IN1(n3011), .IN2(n5134), .IN3(n5133), .IN4(n3009), .Q(n2977)
         );
  OA21X1 U3355 ( .IN1(Datai[20]), .IN2(n2974), .IN3(n2973), .Q(n5135) );
  NAND2X0 U3356 ( .IN1(n3006), .IN2(n5135), .QN(n2976) );
  NAND2X0 U3357 ( .IN1(n3011), .IN2(\DP_OP_469J1_133_8416/n120 ), .QN(n2975)
         );
  NAND4X0 U3358 ( .IN1(n2978), .IN2(n2977), .IN3(n2976), .IN4(n2975), .QN(
        n1892) );
  NAND2X0 U3359 ( .IN1(Datai[3]), .IN2(n3010), .QN(n2986) );
  AOI22X1 U3360 ( .IN1(n4255), .IN2(Datai[3]), .IN3(n2979), .IN4(n5016), .QN(
        n5127) );
  AO21X1 U3361 ( .IN1(n2981), .IN2(n2988), .IN3(n2980), .Q(n5126) );
  OA22X1 U3362 ( .IN1(n3011), .IN2(n5127), .IN3(n5126), .IN4(n3009), .Q(n2985)
         );
  MUX21X1 U3363 ( .IN1(n2982), .IN2(Datai[19]), .S(n2989), .Q(n5128) );
  NAND2X0 U3364 ( .IN1(n3006), .IN2(n5128), .QN(n2984) );
  NAND2X0 U3365 ( .IN1(n3011), .IN2(\DP_OP_469J1_133_8416/n119 ), .QN(n2983)
         );
  NAND4X0 U3366 ( .IN1(n2986), .IN2(n2985), .IN3(n2984), .IN4(n2983), .QN(
        n1893) );
  NAND2X0 U3367 ( .IN1(Datai[2]), .IN2(n3010), .QN(n2993) );
  AOI22X1 U3368 ( .IN1(n4255), .IN2(Datai[2]), .IN3(n2987), .IN4(n5016), .QN(
        n5120) );
  OAI21X1 U3369 ( .IN1(Datai[26]), .IN2(n2996), .IN3(n2988), .QN(n5119) );
  OA22X1 U3370 ( .IN1(n3011), .IN2(n5120), .IN3(n5119), .IN4(n3009), .Q(n2992)
         );
  OA21X1 U3371 ( .IN1(Datai[18]), .IN2(n2994), .IN3(n2989), .Q(n5121) );
  NAND2X0 U3372 ( .IN1(n3006), .IN2(n5121), .QN(n2991) );
  NAND2X0 U3373 ( .IN1(n3011), .IN2(\DP_OP_469J1_133_8416/n118 ), .QN(n2990)
         );
  NAND4X0 U3374 ( .IN1(n2993), .IN2(n2992), .IN3(n2991), .IN4(n2990), .QN(
        n1894) );
  NAND2X0 U3375 ( .IN1(Datai[1]), .IN2(n3010), .QN(n3003) );
  AO21X1 U3376 ( .IN1(n2995), .IN2(n3004), .IN3(n2994), .Q(n5063) );
  AO21X1 U3377 ( .IN1(n2997), .IN2(n3007), .IN3(n2996), .Q(n5112) );
  OA22X1 U3378 ( .IN1(n4556), .IN2(n5063), .IN3(n3009), .IN4(n5112), .Q(n3002)
         );
  AO22X1 U3379 ( .IN1(Datai[1]), .IN2(n4255), .IN3(n5016), .IN4(n2998), .Q(
        n5068) );
  NAND2X0 U3380 ( .IN1(n2999), .IN2(n5068), .QN(n3001) );
  NAND2X0 U3381 ( .IN1(n3011), .IN2(\DP_OP_469J1_133_8416/n117 ), .QN(n3000)
         );
  NAND4X0 U3382 ( .IN1(n3003), .IN2(n3002), .IN3(n3001), .IN4(n3000), .QN(
        n1895) );
  OA21X1 U3383 ( .IN1(Datai[16]), .IN2(n3005), .IN3(n3004), .Q(n5108) );
  NAND2X0 U3384 ( .IN1(n3006), .IN2(n5108), .QN(n3015) );
  INVX0 U3385 ( .INP(Datai[0]), .ZN(n5104) );
  OA22X1 U3386 ( .IN1(n4431), .IN2(n5104), .IN3(n3026), .IN4(n4485), .Q(n5105)
         );
  OAI21X1 U3387 ( .IN1(Datai[24]), .IN2(n3008), .IN3(n3007), .QN(n5100) );
  OA22X1 U3388 ( .IN1(n3011), .IN2(n5105), .IN3(n5100), .IN4(n3009), .Q(n3014)
         );
  NAND2X0 U3389 ( .IN1(Datai[0]), .IN2(n3010), .QN(n3013) );
  NAND2X0 U3390 ( .IN1(n3011), .IN2(\DP_OP_469J1_133_8416/n116 ), .QN(n3012)
         );
  NAND4X0 U3391 ( .IN1(n3015), .IN2(n3014), .IN3(n3013), .IN4(n3012), .QN(
        n1896) );
  NOR2X0 U3392 ( .IN1(State2[3]), .IN2(n4466), .QN(n4495) );
  AO22X1 U3393 ( .IN1(n4445), .IN2(n3016), .IN3(Flush), .IN4(n4495), .Q(n3017)
         );
  NOR2X0 U3394 ( .IN1(n5016), .IN2(n3017), .QN(n4302) );
  MUX21X1 U3395 ( .IN1(n5185), .IN2(InstAddrPointer[1]), .S(n5224), .Q(n4305)
         );
  NAND2X0 U3396 ( .IN1(N1868), .IN2(n4495), .QN(n3019) );
  OA222X1 U3397 ( .IN1(n3020), .IN2(n4485), .IN3(n4305), .IN4(n3019), .IN5(
        n4519), .IN6(n3018), .Q(n3023) );
  INVX0 U3398 ( .INP(n4302), .ZN(n4310) );
  OA22X1 U3399 ( .IN1(n5177), .IN2(n4310), .IN3(n3021), .IN4(n4485), .Q(n3022)
         );
  OAI21X1 U3400 ( .IN1(n4302), .IN2(n3023), .IN3(n3022), .QN(n2027) );
  NOR4X0 U3401 ( .IN1(n3027), .IN2(n3026), .IN3(n3025), .IN4(n3024), .QN(n3175) );
  AO22X1 U3402 ( .IN1(EBX[24]), .IN2(n3175), .IN3(n3053), .IN4(n3028), .Q(
        n3071) );
  AO22X1 U3403 ( .IN1(EBX[23]), .IN2(n3175), .IN3(n3053), .IN4(n3029), .Q(
        n3076) );
  AND2X1 U3404 ( .IN1(n3030), .IN2(n3053), .Q(n3075) );
  AND2X1 U3405 ( .IN1(EBX[22]), .IN2(n3175), .Q(n3080) );
  AND2X1 U3406 ( .IN1(n3031), .IN2(n3053), .Q(n3079) );
  AND2X1 U3407 ( .IN1(EBX[21]), .IN2(n3175), .Q(n3085) );
  AND2X1 U3408 ( .IN1(n3032), .IN2(n3053), .Q(n3084) );
  AND2X1 U3409 ( .IN1(EBX[20]), .IN2(n3175), .Q(n3089) );
  AND2X1 U3410 ( .IN1(n3033), .IN2(n3053), .Q(n3088) );
  AND2X1 U3411 ( .IN1(EBX[19]), .IN2(n3175), .Q(n3093) );
  AND2X1 U3412 ( .IN1(n3034), .IN2(n3053), .Q(n3092) );
  AND2X1 U3413 ( .IN1(EBX[18]), .IN2(n3175), .Q(n3097) );
  AND2X1 U3414 ( .IN1(n3035), .IN2(n3053), .Q(n3096) );
  AND2X1 U3415 ( .IN1(EBX[17]), .IN2(n3175), .Q(n3101) );
  AND2X1 U3416 ( .IN1(n3036), .IN2(n3053), .Q(n3100) );
  AND2X1 U3417 ( .IN1(EBX[16]), .IN2(n3175), .Q(n3105) );
  AND2X1 U3418 ( .IN1(n3037), .IN2(n3053), .Q(n3104) );
  AND2X1 U3419 ( .IN1(EBX[15]), .IN2(n3175), .Q(n3109) );
  AND2X1 U3420 ( .IN1(n3038), .IN2(n3053), .Q(n3108) );
  AND2X1 U3421 ( .IN1(EBX[14]), .IN2(n3175), .Q(n3113) );
  AND2X1 U3422 ( .IN1(n3039), .IN2(n3053), .Q(n3112) );
  AND2X1 U3423 ( .IN1(EBX[13]), .IN2(n3175), .Q(n3117) );
  AND2X1 U3424 ( .IN1(n3040), .IN2(n3053), .Q(n3116) );
  AND2X1 U3425 ( .IN1(EBX[12]), .IN2(n3175), .Q(n3121) );
  AND2X1 U3426 ( .IN1(n3041), .IN2(n3053), .Q(n3120) );
  AND2X1 U3427 ( .IN1(EBX[11]), .IN2(n3175), .Q(n3125) );
  AND2X1 U3428 ( .IN1(n3042), .IN2(n3053), .Q(n3124) );
  AND2X1 U3429 ( .IN1(EBX[10]), .IN2(n3175), .Q(n3129) );
  AND2X1 U3430 ( .IN1(n3043), .IN2(n3053), .Q(n3128) );
  AND2X1 U3431 ( .IN1(EBX[9]), .IN2(n3175), .Q(n3133) );
  AND2X1 U3432 ( .IN1(n3044), .IN2(n3053), .Q(n3132) );
  AND2X1 U3433 ( .IN1(EBX[8]), .IN2(n3175), .Q(n3137) );
  AND2X1 U3434 ( .IN1(n3045), .IN2(n3053), .Q(n3136) );
  AND2X1 U3435 ( .IN1(EBX[7]), .IN2(n3175), .Q(n3141) );
  AND2X1 U3436 ( .IN1(\DP_OP_469J1_133_8416/n123 ), .IN2(n3053), .Q(n3140) );
  AND2X1 U3437 ( .IN1(EBX[6]), .IN2(n3175), .Q(n3145) );
  AND2X1 U3438 ( .IN1(\DP_OP_469J1_133_8416/n122 ), .IN2(n3053), .Q(n3144) );
  AND2X1 U3439 ( .IN1(EBX[5]), .IN2(n3175), .Q(n3149) );
  AND2X1 U3440 ( .IN1(\DP_OP_469J1_133_8416/n121 ), .IN2(n3053), .Q(n3148) );
  AND2X1 U3441 ( .IN1(EBX[4]), .IN2(n3175), .Q(n3153) );
  AND2X1 U3442 ( .IN1(\DP_OP_469J1_133_8416/n120 ), .IN2(n3053), .Q(n3152) );
  AND2X1 U3443 ( .IN1(EBX[3]), .IN2(n3175), .Q(n3157) );
  AND2X1 U3444 ( .IN1(\DP_OP_469J1_133_8416/n119 ), .IN2(n3053), .Q(n3156) );
  AND2X1 U3445 ( .IN1(EBX[2]), .IN2(n3175), .Q(n3161) );
  AND2X1 U3446 ( .IN1(\DP_OP_469J1_133_8416/n118 ), .IN2(n3053), .Q(n3160) );
  AND2X1 U3447 ( .IN1(EBX[1]), .IN2(n3175), .Q(n3165) );
  OR2X1 U3448 ( .IN1(n3175), .IN2(\DP_OP_469J1_133_8416/n116 ), .Q(n3168) );
  AND2X1 U3449 ( .IN1(EBX[0]), .IN2(n3175), .Q(n3167) );
  AND2X1 U3450 ( .IN1(\DP_OP_469J1_133_8416/n117 ), .IN2(n3053), .Q(n3163) );
  AND2X1 U3451 ( .IN1(n3071), .IN2(n3072), .Q(n3069) );
  AO22X1 U3452 ( .IN1(EBX[25]), .IN2(n3175), .IN3(n3053), .IN4(n3046), .Q(
        n3068) );
  AO22X1 U3453 ( .IN1(EBX[26]), .IN2(n3175), .IN3(n3053), .IN4(n3047), .Q(
        n3065) );
  AO22X1 U3454 ( .IN1(EBX[27]), .IN2(n3175), .IN3(n3053), .IN4(n3048), .Q(
        n3062) );
  AO22X1 U3455 ( .IN1(EBX[28]), .IN2(n3175), .IN3(n3053), .IN4(n3049), .Q(
        n3059) );
  AO22X1 U3456 ( .IN1(EBX[29]), .IN2(n3175), .IN3(n3053), .IN4(n3050), .Q(
        n3056) );
  AO22X1 U3457 ( .IN1(EBX[30]), .IN2(n3175), .IN3(n3053), .IN4(n3051), .Q(
        n3171) );
  AO21X1 U3458 ( .IN1(n3053), .IN2(n3052), .IN3(n3175), .Q(n3054) );
  AND2X1 U3459 ( .IN1(n4445), .IN2(n3054), .Q(n3081) );
  INVX0 U3460 ( .INP(n3081), .ZN(n3169) );
  MUX21X1 U3461 ( .IN1(n3055), .IN2(EBX[30]), .S(n3169), .Q(n1858) );
  HADDX1 U3462 ( .A0(n3057), .B0(n3056), .C1(n3172), .SO(n3058) );
  MUX21X1 U3463 ( .IN1(n3058), .IN2(EBX[29]), .S(n3169), .Q(n1859) );
  HADDX1 U3464 ( .A0(n3060), .B0(n3059), .C1(n3057), .SO(n3061) );
  MUX21X1 U3465 ( .IN1(n3061), .IN2(EBX[28]), .S(n3169), .Q(n1860) );
  HADDX1 U3466 ( .A0(n3063), .B0(n3062), .C1(n3060), .SO(n3064) );
  MUX21X1 U3467 ( .IN1(n3064), .IN2(EBX[27]), .S(n3169), .Q(n1861) );
  HADDX1 U3468 ( .A0(n3066), .B0(n3065), .C1(n3063), .SO(n3067) );
  MUX21X1 U3469 ( .IN1(n3067), .IN2(EBX[26]), .S(n3169), .Q(n1862) );
  HADDX1 U3470 ( .A0(n3069), .B0(n3068), .C1(n3066), .SO(n3070) );
  MUX21X1 U3471 ( .IN1(n3070), .IN2(EBX[25]), .S(n3169), .Q(n1863) );
  XOR2X1 U3472 ( .IN1(n3072), .IN2(n3071), .Q(n3073) );
  MUX21X1 U3473 ( .IN1(n3073), .IN2(EBX[24]), .S(n3169), .Q(n1864) );
  FADDX1 U3474 ( .A(n3076), .B(n3075), .CI(n3074), .CO(n3072), .S(n3077) );
  MUX21X1 U3475 ( .IN1(n3077), .IN2(EBX[23]), .S(n3169), .Q(n1865) );
  FADDX1 U3476 ( .A(n3080), .B(n3079), .CI(n3078), .CO(n3074), .S(n3082) );
  INVX0 U3477 ( .INP(n3081), .ZN(n3176) );
  MUX21X1 U3478 ( .IN1(n3082), .IN2(EBX[22]), .S(n3176), .Q(n1866) );
  FADDX1 U3479 ( .A(n3085), .B(n3084), .CI(n3083), .CO(n3078), .S(n3086) );
  MUX21X1 U3480 ( .IN1(n3086), .IN2(EBX[21]), .S(n3176), .Q(n1867) );
  FADDX1 U3481 ( .A(n3089), .B(n3088), .CI(n3087), .CO(n3083), .S(n3090) );
  MUX21X1 U3482 ( .IN1(n3090), .IN2(EBX[20]), .S(n3176), .Q(n1868) );
  FADDX1 U3483 ( .A(n3093), .B(n3092), .CI(n3091), .CO(n3087), .S(n3094) );
  MUX21X1 U3484 ( .IN1(n3094), .IN2(EBX[19]), .S(n3176), .Q(n1869) );
  FADDX1 U3485 ( .A(n3097), .B(n3096), .CI(n3095), .CO(n3091), .S(n3098) );
  MUX21X1 U3486 ( .IN1(n3098), .IN2(EBX[18]), .S(n3176), .Q(n1870) );
  FADDX1 U3487 ( .A(n3101), .B(n3100), .CI(n3099), .CO(n3095), .S(n3102) );
  MUX21X1 U3488 ( .IN1(n3102), .IN2(EBX[17]), .S(n3176), .Q(n1871) );
  FADDX1 U3489 ( .A(n3105), .B(n3104), .CI(n3103), .CO(n3099), .S(n3106) );
  MUX21X1 U3490 ( .IN1(n3106), .IN2(EBX[16]), .S(n3176), .Q(n1872) );
  FADDX1 U3491 ( .A(n3109), .B(n3108), .CI(n3107), .CO(n3103), .S(n3110) );
  MUX21X1 U3492 ( .IN1(n3110), .IN2(EBX[15]), .S(n3176), .Q(n1873) );
  FADDX1 U3493 ( .A(n3113), .B(n3112), .CI(n3111), .CO(n3107), .S(n3114) );
  MUX21X1 U3494 ( .IN1(n3114), .IN2(EBX[14]), .S(n3176), .Q(n1874) );
  FADDX1 U3495 ( .A(n3117), .B(n3116), .CI(n3115), .CO(n3111), .S(n3118) );
  MUX21X1 U3496 ( .IN1(n3118), .IN2(EBX[13]), .S(n3176), .Q(n1875) );
  FADDX1 U3497 ( .A(n3121), .B(n3120), .CI(n3119), .CO(n3115), .S(n3122) );
  MUX21X1 U3498 ( .IN1(n3122), .IN2(EBX[12]), .S(n3176), .Q(n1876) );
  FADDX1 U3499 ( .A(n3125), .B(n3124), .CI(n3123), .CO(n3119), .S(n3126) );
  MUX21X1 U3500 ( .IN1(n3126), .IN2(EBX[11]), .S(n3176), .Q(n1877) );
  FADDX1 U3501 ( .A(n3129), .B(n3128), .CI(n3127), .CO(n3123), .S(n3130) );
  MUX21X1 U3502 ( .IN1(n3130), .IN2(EBX[10]), .S(n3169), .Q(n1878) );
  FADDX1 U3503 ( .A(n3133), .B(n3132), .CI(n3131), .CO(n3127), .S(n3134) );
  MUX21X1 U3504 ( .IN1(n3134), .IN2(EBX[9]), .S(n3169), .Q(n1879) );
  FADDX1 U3505 ( .A(n3137), .B(n3136), .CI(n3135), .CO(n3131), .S(n3138) );
  MUX21X1 U3506 ( .IN1(n3138), .IN2(EBX[8]), .S(n3169), .Q(n1880) );
  FADDX1 U3507 ( .A(n3141), .B(n3140), .CI(n3139), .CO(n3135), .S(n3142) );
  MUX21X1 U3508 ( .IN1(n3142), .IN2(EBX[7]), .S(n3169), .Q(n1881) );
  FADDX1 U3509 ( .A(n3145), .B(n3144), .CI(n3143), .CO(n3139), .S(n3146) );
  MUX21X1 U3510 ( .IN1(n3146), .IN2(EBX[6]), .S(n3169), .Q(n1882) );
  FADDX1 U3511 ( .A(n3149), .B(n3148), .CI(n3147), .CO(n3143), .S(n3150) );
  MUX21X1 U3512 ( .IN1(n3150), .IN2(EBX[5]), .S(n3176), .Q(n1883) );
  FADDX1 U3513 ( .A(n3153), .B(n3152), .CI(n3151), .CO(n3147), .S(n3154) );
  MUX21X1 U3514 ( .IN1(n3154), .IN2(EBX[4]), .S(n3169), .Q(n1884) );
  FADDX1 U3515 ( .A(n3157), .B(n3156), .CI(n3155), .CO(n3151), .S(n3158) );
  MUX21X1 U3516 ( .IN1(n3158), .IN2(EBX[3]), .S(n3176), .Q(n1885) );
  FADDX1 U3517 ( .A(n3161), .B(n3160), .CI(n3159), .CO(n3155), .S(n3162) );
  MUX21X1 U3518 ( .IN1(n3162), .IN2(EBX[2]), .S(n3169), .Q(n1886) );
  FADDX1 U3519 ( .A(n3165), .B(n3164), .CI(n3163), .CO(n3159), .S(n3166) );
  MUX21X1 U3520 ( .IN1(n3166), .IN2(EBX[1]), .S(n3176), .Q(n1887) );
  HADDX1 U3521 ( .A0(n3168), .B0(n3167), .C1(n3164), .SO(n3170) );
  MUX21X1 U3522 ( .IN1(n3170), .IN2(EBX[0]), .S(n3169), .Q(n1888) );
  HADDX1 U3523 ( .A0(n3172), .B0(n3171), .C1(n3173), .SO(n3055) );
  XOR2X1 U3524 ( .IN1(n3173), .IN2(N1989), .Q(n3174) );
  AND2X1 U3525 ( .IN1(n3175), .IN2(n3174), .Q(n3177) );
  MUX21X1 U3526 ( .IN1(n3177), .IN2(N1989), .S(n3176), .Q(n1857) );
  INVX0 U3527 ( .INP(n4104), .ZN(n4147) );
  NAND2X0 U3528 ( .IN1(n4515), .IN2(n3178), .QN(n4488) );
  NAND4X0 U3529 ( .IN1(n4147), .IN2(n4470), .IN3(n3288), .IN4(n4488), .QN(
        n4280) );
  HADDX1 U3530 ( .A0(n3179), .B0(PhyAddrPointer[30]), .C1(n3180), .SO(n3315)
         );
  XOR2X1 U3531 ( .IN1(n3180), .IN2(PhyAddrPointer[31]), .Q(n4254) );
  NAND2X0 U3532 ( .IN1(n4977), .IN2(n4254), .QN(n3186) );
  INVX0 U3533 ( .INP(n3186), .ZN(n3279) );
  INVX0 U3534 ( .INP(n3286), .ZN(n3183) );
  INVX0 U3535 ( .INP(n3284), .ZN(n3181) );
  NAND2X0 U3536 ( .IN1(n3181), .IN2(N1989), .QN(n3182) );
  OR2X1 U3537 ( .IN1(n3183), .IN2(n3182), .Q(n3185) );
  INVX0 U3538 ( .INP(n3185), .ZN(n3277) );
  OAI21X1 U3539 ( .IN1(n3286), .IN2(n3284), .IN3(n4446), .QN(n4229) );
  AO22X1 U3540 ( .IN1(n3277), .IN2(EBX[30]), .IN3(rEIP[30]), .IN4(n4229), .Q(
        n3184) );
  AO21X1 U3541 ( .IN1(n3315), .IN2(n3279), .IN3(n3184), .Q(n3187) );
  NAND2X1 U3542 ( .IN1(n3186), .IN2(n3185), .QN(n4278) );
  XOR2X1 U3543 ( .IN1(n3187), .IN2(n4278), .Q(n3312) );
  HADDX1 U3544 ( .A0(n3188), .B0(PhyAddrPointer[29]), .C1(n3179), .SO(n3368)
         );
  AO22X1 U3545 ( .IN1(n3277), .IN2(EBX[29]), .IN3(rEIP[29]), .IN4(n4229), .Q(
        n3189) );
  AO21X1 U3546 ( .IN1(n3368), .IN2(n3279), .IN3(n3189), .Q(n3190) );
  XOR2X1 U3547 ( .IN1(n3190), .IN2(n4278), .Q(n3366) );
  HADDX1 U3548 ( .A0(n3191), .B0(PhyAddrPointer[28]), .C1(n3188), .SO(n3404)
         );
  AO22X1 U3549 ( .IN1(n3277), .IN2(EBX[28]), .IN3(rEIP[28]), .IN4(n4229), .Q(
        n3192) );
  AO21X1 U3550 ( .IN1(n3404), .IN2(n3279), .IN3(n3192), .Q(n3193) );
  XOR2X1 U3551 ( .IN1(n3193), .IN2(n4278), .Q(n3402) );
  HADDX1 U3552 ( .A0(n3194), .B0(PhyAddrPointer[27]), .C1(n3191), .SO(n3385)
         );
  AO22X1 U3553 ( .IN1(n3277), .IN2(EBX[27]), .IN3(rEIP[27]), .IN4(n4229), .Q(
        n3195) );
  AO21X1 U3554 ( .IN1(n3385), .IN2(n3279), .IN3(n3195), .Q(n3196) );
  XOR2X1 U3555 ( .IN1(n3196), .IN2(n4278), .Q(n3374) );
  HADDX1 U3556 ( .A0(n3197), .B0(PhyAddrPointer[26]), .C1(n3194), .SO(n3440)
         );
  AO22X1 U3557 ( .IN1(n3277), .IN2(EBX[26]), .IN3(rEIP[26]), .IN4(n4229), .Q(
        n3198) );
  AO21X1 U3558 ( .IN1(n3440), .IN2(n3279), .IN3(n3198), .Q(n3199) );
  XOR2X1 U3559 ( .IN1(n3199), .IN2(n4278), .Q(n3438) );
  HADDX1 U3560 ( .A0(n3200), .B0(PhyAddrPointer[25]), .C1(n3197), .SO(n3421)
         );
  AO22X1 U3561 ( .IN1(n3277), .IN2(EBX[25]), .IN3(rEIP[25]), .IN4(n4229), .Q(
        n3201) );
  AO21X1 U3562 ( .IN1(n3421), .IN2(n3279), .IN3(n3201), .Q(n3202) );
  XOR2X1 U3563 ( .IN1(n3202), .IN2(n4278), .Q(n3410) );
  HADDX1 U3564 ( .A0(n3203), .B0(PhyAddrPointer[24]), .C1(n3200), .SO(n3476)
         );
  AO22X1 U3565 ( .IN1(n3277), .IN2(EBX[24]), .IN3(rEIP[24]), .IN4(n4229), .Q(
        n3204) );
  AO21X1 U3566 ( .IN1(n3476), .IN2(n3279), .IN3(n3204), .Q(n3205) );
  XOR2X1 U3567 ( .IN1(n3205), .IN2(n4278), .Q(n3474) );
  HADDX1 U3568 ( .A0(n3206), .B0(PhyAddrPointer[23]), .C1(n3203), .SO(n3457)
         );
  AO22X1 U3569 ( .IN1(n3277), .IN2(EBX[23]), .IN3(rEIP[23]), .IN4(n4229), .Q(
        n3207) );
  AO21X1 U3570 ( .IN1(n3457), .IN2(n3279), .IN3(n3207), .Q(n3208) );
  XOR2X1 U3571 ( .IN1(n3208), .IN2(n4278), .Q(n3446) );
  HADDX1 U3572 ( .A0(n3209), .B0(PhyAddrPointer[22]), .C1(n3206), .SO(n3512)
         );
  AO22X1 U3573 ( .IN1(n3277), .IN2(EBX[22]), .IN3(rEIP[22]), .IN4(n4229), .Q(
        n3210) );
  AO21X1 U3574 ( .IN1(n3512), .IN2(n3279), .IN3(n3210), .Q(n3211) );
  XOR2X1 U3575 ( .IN1(n3211), .IN2(n4278), .Q(n3510) );
  HADDX1 U3576 ( .A0(n3212), .B0(PhyAddrPointer[21]), .C1(n3209), .SO(n3493)
         );
  AO22X1 U3577 ( .IN1(n3277), .IN2(EBX[21]), .IN3(rEIP[21]), .IN4(n4229), .Q(
        n3213) );
  AO21X1 U3578 ( .IN1(n3493), .IN2(n3279), .IN3(n3213), .Q(n3214) );
  XOR2X1 U3579 ( .IN1(n3214), .IN2(n4278), .Q(n3482) );
  HADDX1 U3580 ( .A0(n3215), .B0(PhyAddrPointer[20]), .C1(n3212), .SO(n3548)
         );
  AO22X1 U3581 ( .IN1(n3277), .IN2(EBX[20]), .IN3(rEIP[20]), .IN4(n4229), .Q(
        n3216) );
  AO21X1 U3582 ( .IN1(n3548), .IN2(n3279), .IN3(n3216), .Q(n3217) );
  XOR2X1 U3583 ( .IN1(n3217), .IN2(n4278), .Q(n3546) );
  HADDX1 U3584 ( .A0(n3218), .B0(PhyAddrPointer[19]), .C1(n3215), .SO(n3530)
         );
  AO22X1 U3585 ( .IN1(n3277), .IN2(EBX[19]), .IN3(rEIP[19]), .IN4(n4229), .Q(
        n3219) );
  AO21X1 U3586 ( .IN1(n3530), .IN2(n3279), .IN3(n3219), .Q(n3220) );
  XOR2X1 U3587 ( .IN1(n3220), .IN2(n4278), .Q(n3520) );
  HADDX1 U3588 ( .A0(n3221), .B0(PhyAddrPointer[18]), .C1(n3218), .SO(n3709)
         );
  AO22X1 U3589 ( .IN1(n3277), .IN2(EBX[18]), .IN3(rEIP[18]), .IN4(n4229), .Q(
        n3222) );
  AO21X1 U3590 ( .IN1(n3709), .IN2(n3279), .IN3(n3222), .Q(n3223) );
  XOR2X1 U3591 ( .IN1(n3223), .IN2(n4278), .Q(n3708) );
  HADDX1 U3592 ( .A0(n3224), .B0(PhyAddrPointer[17]), .C1(n3221), .SO(n3692)
         );
  AO22X1 U3593 ( .IN1(n3277), .IN2(EBX[17]), .IN3(rEIP[17]), .IN4(n4229), .Q(
        n3225) );
  AO21X1 U3594 ( .IN1(n3692), .IN2(n3279), .IN3(n3225), .Q(n3226) );
  XOR2X1 U3595 ( .IN1(n3226), .IN2(n4278), .Q(n3681) );
  HADDX1 U3596 ( .A0(n3227), .B0(PhyAddrPointer[16]), .C1(n3224), .SO(n3771)
         );
  AO22X1 U3597 ( .IN1(n3277), .IN2(EBX[16]), .IN3(rEIP[16]), .IN4(n4229), .Q(
        n3228) );
  AO21X1 U3598 ( .IN1(n3771), .IN2(n3279), .IN3(n3228), .Q(n3229) );
  XOR2X1 U3599 ( .IN1(n3229), .IN2(n4278), .Q(n3770) );
  HADDX1 U3600 ( .A0(n3230), .B0(PhyAddrPointer[15]), .C1(n3227), .SO(n3754)
         );
  AO22X1 U3601 ( .IN1(n3277), .IN2(EBX[15]), .IN3(rEIP[15]), .IN4(n4229), .Q(
        n3231) );
  AO21X1 U3602 ( .IN1(n3754), .IN2(n3279), .IN3(n3231), .Q(n3232) );
  XOR2X1 U3603 ( .IN1(n3232), .IN2(n4278), .Q(n3744) );
  HADDX1 U3604 ( .A0(n3233), .B0(PhyAddrPointer[14]), .C1(n3230), .SO(n3833)
         );
  AO22X1 U3605 ( .IN1(n3277), .IN2(EBX[14]), .IN3(rEIP[14]), .IN4(n4229), .Q(
        n3234) );
  AO21X1 U3606 ( .IN1(n3833), .IN2(n3279), .IN3(n3234), .Q(n3235) );
  XOR2X1 U3607 ( .IN1(n3235), .IN2(n4278), .Q(n3832) );
  HADDX1 U3608 ( .A0(n3236), .B0(PhyAddrPointer[13]), .C1(n3233), .SO(n3815)
         );
  AO22X1 U3609 ( .IN1(n3277), .IN2(EBX[13]), .IN3(rEIP[13]), .IN4(n4229), .Q(
        n3237) );
  AO21X1 U3610 ( .IN1(n3815), .IN2(n3279), .IN3(n3237), .Q(n3238) );
  XOR2X1 U3611 ( .IN1(n3238), .IN2(n4278), .Q(n3805) );
  HADDX1 U3612 ( .A0(n3239), .B0(PhyAddrPointer[12]), .C1(n3236), .SO(n3895)
         );
  AO22X1 U3613 ( .IN1(n3277), .IN2(EBX[12]), .IN3(rEIP[12]), .IN4(n4229), .Q(
        n3240) );
  AO21X1 U3614 ( .IN1(n3895), .IN2(n3279), .IN3(n3240), .Q(n3241) );
  XOR2X1 U3615 ( .IN1(n3241), .IN2(n4278), .Q(n3894) );
  HADDX1 U3616 ( .A0(n3242), .B0(PhyAddrPointer[11]), .C1(n3239), .SO(n3877)
         );
  AO22X1 U3617 ( .IN1(n3277), .IN2(EBX[11]), .IN3(rEIP[11]), .IN4(n4229), .Q(
        n3243) );
  AO21X1 U3618 ( .IN1(n3877), .IN2(n3279), .IN3(n3243), .Q(n3244) );
  XOR2X1 U3619 ( .IN1(n3244), .IN2(n4278), .Q(n3867) );
  HADDX1 U3620 ( .A0(n3245), .B0(PhyAddrPointer[10]), .C1(n3242), .SO(n3958)
         );
  AO22X1 U3621 ( .IN1(n3277), .IN2(EBX[10]), .IN3(rEIP[10]), .IN4(n4229), .Q(
        n3246) );
  AO21X1 U3622 ( .IN1(n3958), .IN2(n3279), .IN3(n3246), .Q(n3247) );
  XOR2X1 U3623 ( .IN1(n3247), .IN2(n4278), .Q(n3957) );
  HADDX1 U3624 ( .A0(n3248), .B0(PhyAddrPointer[9]), .C1(n3245), .SO(n3939) );
  AO22X1 U3625 ( .IN1(n3277), .IN2(EBX[9]), .IN3(rEIP[9]), .IN4(n4229), .Q(
        n3249) );
  AO21X1 U3626 ( .IN1(n3939), .IN2(n3279), .IN3(n3249), .Q(n3250) );
  XOR2X1 U3627 ( .IN1(n3250), .IN2(n4278), .Q(n3929) );
  HADDX1 U3628 ( .A0(n3251), .B0(PhyAddrPointer[8]), .C1(n3248), .SO(n4003) );
  AO22X1 U3629 ( .IN1(n3277), .IN2(EBX[8]), .IN3(rEIP[8]), .IN4(n4229), .Q(
        n3252) );
  AO21X1 U3630 ( .IN1(n4003), .IN2(n3279), .IN3(n3252), .Q(n3253) );
  XOR2X1 U3631 ( .IN1(n3253), .IN2(n4278), .Q(n4002) );
  HADDX1 U3632 ( .A0(n3254), .B0(PhyAddrPointer[7]), .C1(n3251), .SO(n4144) );
  AO22X1 U3633 ( .IN1(rEIP[7]), .IN2(n4229), .IN3(EBX[7]), .IN4(n3277), .Q(
        n3255) );
  AO21X1 U3634 ( .IN1(n4144), .IN2(n3279), .IN3(n3255), .Q(n3256) );
  XOR2X1 U3635 ( .IN1(n3256), .IN2(n4278), .Q(n4143) );
  HADDX1 U3636 ( .A0(n3257), .B0(PhyAddrPointer[6]), .C1(n3254), .SO(n4126) );
  AO22X1 U3637 ( .IN1(rEIP[6]), .IN2(n4229), .IN3(EBX[6]), .IN4(n3277), .Q(
        n3258) );
  AO21X1 U3638 ( .IN1(n4126), .IN2(n3279), .IN3(n3258), .Q(n3259) );
  XOR2X1 U3639 ( .IN1(n3259), .IN2(n4278), .Q(n4110) );
  HADDX1 U3640 ( .A0(n3260), .B0(PhyAddrPointer[5]), .C1(n3257), .SO(n4103) );
  AO22X1 U3641 ( .IN1(rEIP[5]), .IN2(n4229), .IN3(EBX[5]), .IN4(n3277), .Q(
        n3261) );
  AO21X1 U3642 ( .IN1(n4103), .IN2(n3279), .IN3(n3261), .Q(n3262) );
  XOR2X1 U3643 ( .IN1(n3262), .IN2(n4278), .Q(n4092) );
  HADDX1 U3644 ( .A0(n3263), .B0(PhyAddrPointer[4]), .C1(n3260), .SO(n4086) );
  NAND2X0 U3645 ( .IN1(n4229), .IN2(rEIP[4]), .QN(n3265) );
  NAND2X0 U3646 ( .IN1(EBX[4]), .IN2(n3277), .QN(n3264) );
  NAND2X0 U3647 ( .IN1(n3265), .IN2(n3264), .QN(n3266) );
  AO21X1 U3648 ( .IN1(n4086), .IN2(n3279), .IN3(n3266), .Q(n3267) );
  XOR2X1 U3649 ( .IN1(n3267), .IN2(n4278), .Q(n4072) );
  HADDX1 U3650 ( .A0(n3268), .B0(PhyAddrPointer[3]), .C1(n3263), .SO(n4053) );
  AO222X1 U3651 ( .IN1(n4229), .IN2(rEIP[3]), .IN3(n4277), .IN4(
        InstQueueRd_Addr[3]), .IN5(EBX[3]), .IN6(n3277), .Q(n3269) );
  AO21X1 U3652 ( .IN1(n4053), .IN2(n3279), .IN3(n3269), .Q(n3270) );
  XOR2X1 U3653 ( .IN1(n3270), .IN2(n4278), .Q(n4051) );
  HADDX1 U3654 ( .A0(PhyAddrPointer[1]), .B0(PhyAddrPointer[2]), .C1(n3268), 
        .SO(n4036) );
  AO222X1 U3655 ( .IN1(n4229), .IN2(rEIP[2]), .IN3(n4277), .IN4(
        InstQueueRd_Addr[2]), .IN5(n3277), .IN6(EBX[2]), .Q(n3271) );
  AO21X1 U3656 ( .IN1(n4036), .IN2(n3279), .IN3(n3271), .Q(n3272) );
  XOR2X1 U3657 ( .IN1(n3272), .IN2(n4278), .Q(n4023) );
  AO222X1 U3658 ( .IN1(n4229), .IN2(N4154), .IN3(EBX[1]), .IN4(n3277), .IN5(
        InstQueueRd_Addr[1]), .IN6(n4277), .Q(n3273) );
  AO21X1 U3659 ( .IN1(n5201), .IN2(n3279), .IN3(n3273), .Q(n3274) );
  XOR2X1 U3660 ( .IN1(n3274), .IN2(n4278), .Q(n4228) );
  AO222X1 U3661 ( .IN1(n4229), .IN2(rEIP[0]), .IN3(EBX[0]), .IN4(n3277), .IN5(
        N2884), .IN6(n4277), .Q(n3275) );
  AO21X1 U3662 ( .IN1(N1009), .IN2(n3279), .IN3(n3275), .Q(n3276) );
  XOR2X1 U3663 ( .IN1(n3276), .IN2(n4278), .Q(n4276) );
  AND2X1 U3664 ( .IN1(n4023), .IN2(n4022), .Q(n4050) );
  AND2X1 U3665 ( .IN1(n4051), .IN2(n4050), .Q(n4071) );
  AND2X1 U3666 ( .IN1(n4072), .IN2(n4071), .Q(n4091) );
  AND2X1 U3667 ( .IN1(n4092), .IN2(n4091), .Q(n4109) );
  AND2X1 U3668 ( .IN1(n4110), .IN2(n4109), .Q(n4142) );
  AND2X1 U3669 ( .IN1(n4143), .IN2(n4142), .Q(n4001) );
  AND2X1 U3670 ( .IN1(n4002), .IN2(n4001), .Q(n3928) );
  AND2X1 U3671 ( .IN1(n3929), .IN2(n3928), .Q(n3956) );
  AND2X1 U3672 ( .IN1(n3957), .IN2(n3956), .Q(n3866) );
  AND2X1 U3673 ( .IN1(n3867), .IN2(n3866), .Q(n3893) );
  AND2X1 U3674 ( .IN1(n3894), .IN2(n3893), .Q(n3804) );
  AND2X1 U3675 ( .IN1(n3805), .IN2(n3804), .Q(n3831) );
  AND2X1 U3676 ( .IN1(n3832), .IN2(n3831), .Q(n3743) );
  AND2X1 U3677 ( .IN1(n3744), .IN2(n3743), .Q(n3769) );
  AND2X1 U3678 ( .IN1(n3770), .IN2(n3769), .Q(n3680) );
  AND2X1 U3679 ( .IN1(n3681), .IN2(n3680), .Q(n3707) );
  AND2X1 U3680 ( .IN1(n3708), .IN2(n3707), .Q(n3519) );
  AND2X1 U3681 ( .IN1(n3520), .IN2(n3519), .Q(n3545) );
  AND2X1 U3682 ( .IN1(n3546), .IN2(n3545), .Q(n3481) );
  AND2X1 U3683 ( .IN1(n3482), .IN2(n3481), .Q(n3509) );
  AND2X1 U3684 ( .IN1(n3510), .IN2(n3509), .Q(n3445) );
  AND2X1 U3685 ( .IN1(n3446), .IN2(n3445), .Q(n3473) );
  AND2X1 U3686 ( .IN1(n3474), .IN2(n3473), .Q(n3409) );
  AND2X1 U3687 ( .IN1(n3410), .IN2(n3409), .Q(n3437) );
  AND2X1 U3688 ( .IN1(n3438), .IN2(n3437), .Q(n3373) );
  AND2X1 U3689 ( .IN1(n3374), .IN2(n3373), .Q(n3401) );
  AND2X1 U3690 ( .IN1(n3402), .IN2(n3401), .Q(n3365) );
  AND2X1 U3691 ( .IN1(n3366), .IN2(n3365), .Q(n3311) );
  AND2X1 U3692 ( .IN1(n3312), .IN2(n3311), .Q(n3282) );
  AO21X1 U3693 ( .IN1(rEIP[31]), .IN2(n4229), .IN3(n3277), .Q(n3278) );
  OR2X1 U3694 ( .IN1(n3279), .IN2(n3278), .Q(n3280) );
  XOR2X1 U3695 ( .IN1(n3280), .IN2(n4278), .Q(n3281) );
  XOR2X1 U3696 ( .IN1(n3282), .IN2(n3281), .Q(n3283) );
  NAND2X0 U3697 ( .IN1(n4280), .IN2(n3283), .QN(n3292) );
  INVX0 U3698 ( .INP(n4280), .ZN(n4281) );
  NAND2X0 U3699 ( .IN1(rEIP[31]), .IN2(n4281), .QN(n3291) );
  NOR2X0 U3700 ( .IN1(N1989), .IN2(n3284), .QN(n3285) );
  AO222X1 U3701 ( .IN1(n4443), .IN2(n3286), .IN3(n4443), .IN4(n4518), .IN5(
        n3286), .IN6(n3285), .Q(n3287) );
  AND2X1 U3702 ( .IN1(n4280), .IN2(n3287), .Q(n4275) );
  NAND2X0 U3703 ( .IN1(N1989), .IN2(n4275), .QN(n3290) );
  INVX0 U3704 ( .INP(n3288), .ZN(n4274) );
  NAND2X0 U3705 ( .IN1(n4274), .IN2(PhyAddrPointer[31]), .QN(n3289) );
  NAND4X0 U3706 ( .IN1(n3292), .IN2(n3291), .IN3(n3290), .IN4(n3289), .QN(
        n2071) );
  OAI21X1 U3707 ( .IN1(n3293), .IN2(n4519), .IN3(n4450), .QN(n4221) );
  NAND2X0 U3708 ( .IN1(n4445), .IN2(n4221), .QN(n3294) );
  NOR2X0 U3709 ( .IN1(n3295), .IN2(n3294), .QN(n4266) );
  HADDX1 U3710 ( .A0(n3296), .B0(InstAddrPointer[29]), .C1(n3336), .SO(n2927)
         );
  HADDX1 U3711 ( .A0(n3297), .B0(InstAddrPointer[29]), .C1(n3338), .SO(n2829)
         );
  AO22X1 U3712 ( .IN1(n4132), .IN2(n3323), .IN3(n3298), .IN4(n2916), .Q(n3343)
         );
  FADDX1 U3713 ( .A(n3993), .B(n3300), .CI(n3299), .CO(n3342), .S(n2921) );
  NAND3X0 U3714 ( .IN1(n4445), .IN2(n3301), .IN3(n4221), .QN(n4252) );
  NOR2X0 U3715 ( .IN1(n3302), .IN2(n5223), .QN(n3332) );
  MUX21X1 U3716 ( .IN1(n5230), .IN2(InstAddrPointer[30]), .S(n3332), .Q(n3321)
         );
  NOR2X0 U3717 ( .IN1(n3321), .IN2(n3303), .QN(n3334) );
  AO21X1 U3718 ( .IN1(n3321), .IN2(n3303), .IN3(n3334), .Q(n3320) );
  NOR2X0 U3719 ( .IN1(n4252), .IN2(n3320), .QN(n3304) );
  AOI21X1 U3720 ( .IN1(n4266), .IN2(n3322), .IN3(n3304), .QN(n3310) );
  AND3X1 U3721 ( .IN1(PhyAddrPointer[3]), .IN2(PhyAddrPointer[2]), .IN3(
        PhyAddrPointer[4]), .Q(n4122) );
  NAND2X0 U3722 ( .IN1(n4122), .IN2(PhyAddrPointer[5]), .QN(n3305) );
  NOR2X0 U3723 ( .IN1(n3305), .IN2(n5184), .QN(n4136) );
  NAND2X0 U3724 ( .IN1(n4136), .IN2(PhyAddrPointer[7]), .QN(n3996) );
  NOR2X0 U3725 ( .IN1(n3996), .IN2(n5189), .QN(n3937) );
  AND3X1 U3726 ( .IN1(n3937), .IN2(PhyAddrPointer[10]), .IN3(PhyAddrPointer[9]), .Q(n3875) );
  AND3X1 U3727 ( .IN1(n3875), .IN2(PhyAddrPointer[12]), .IN3(
        PhyAddrPointer[11]), .Q(n3813) );
  AND3X1 U3728 ( .IN1(n3813), .IN2(PhyAddrPointer[14]), .IN3(
        PhyAddrPointer[13]), .Q(n3764) );
  AND3X1 U3729 ( .IN1(n3764), .IN2(PhyAddrPointer[16]), .IN3(
        PhyAddrPointer[15]), .Q(n3703) );
  AND3X1 U3730 ( .IN1(n3703), .IN2(PhyAddrPointer[18]), .IN3(
        PhyAddrPointer[17]), .Q(n3541) );
  AND3X1 U3731 ( .IN1(n3541), .IN2(PhyAddrPointer[20]), .IN3(
        PhyAddrPointer[19]), .Q(n3504) );
  AND3X1 U3732 ( .IN1(n3504), .IN2(PhyAddrPointer[22]), .IN3(
        PhyAddrPointer[21]), .Q(n3468) );
  AND3X1 U3733 ( .IN1(n3468), .IN2(PhyAddrPointer[24]), .IN3(
        PhyAddrPointer[23]), .Q(n3432) );
  AND3X1 U3734 ( .IN1(n3432), .IN2(PhyAddrPointer[26]), .IN3(
        PhyAddrPointer[25]), .Q(n3396) );
  AND3X1 U3735 ( .IN1(n3396), .IN2(PhyAddrPointer[28]), .IN3(
        PhyAddrPointer[27]), .Q(n3306) );
  NAND2X0 U3736 ( .IN1(n5098), .IN2(n3306), .QN(n3360) );
  NOR2X0 U3737 ( .IN1(n5240), .IN2(n3360), .QN(n4253) );
  INVX0 U3738 ( .INP(n4253), .ZN(n3307) );
  OA21X1 U3739 ( .IN1(n3306), .IN2(n5020), .IN3(n4221), .Q(n3359) );
  OA21X1 U3740 ( .IN1(PhyAddrPointer[29]), .IN2(n5020), .IN3(n3359), .Q(n4245)
         );
  MUX21X1 U3741 ( .IN1(n3307), .IN2(n4245), .S(PhyAddrPointer[30]), .Q(n3309)
         );
  NAND2X0 U3742 ( .IN1(n4104), .IN2(rEIP[30]), .QN(n3329) );
  NAND2X0 U3743 ( .IN1(n4255), .IN2(n3315), .QN(n3308) );
  NAND4X0 U3744 ( .IN1(n3310), .IN2(n3309), .IN3(n3329), .IN4(n3308), .QN(
        n1706) );
  AOI22X1 U3745 ( .IN1(n4275), .IN2(EBX[30]), .IN3(n4274), .IN4(
        PhyAddrPointer[30]), .QN(n3319) );
  XOR2X1 U3746 ( .IN1(n3312), .IN2(n3311), .Q(n3313) );
  NAND2X0 U3747 ( .IN1(n4280), .IN2(n3313), .QN(n3318) );
  INVX0 U3748 ( .INP(n4254), .ZN(n3314) );
  NAND2X0 U3749 ( .IN1(n2090), .IN2(n3315), .QN(n3317) );
  NAND2X0 U3750 ( .IN1(rEIP[30]), .IN2(n4281), .QN(n3316) );
  NAND4X0 U3751 ( .IN1(n3319), .IN2(n3318), .IN3(n3317), .IN4(n3316), .QN(
        n2035) );
  OA22X1 U3752 ( .IN1(n3321), .IN2(n4206), .IN3(n4208), .IN4(n3320), .Q(n3326)
         );
  INVX0 U3753 ( .INP(n4060), .ZN(n4288) );
  NAND2X0 U3754 ( .IN1(n3322), .IN2(n4288), .QN(n3325) );
  NAND2X0 U3755 ( .IN1(n4290), .IN2(n3323), .QN(n3324) );
  AND3X1 U3756 ( .IN1(n3326), .IN2(n3325), .IN3(n3324), .Q(n3331) );
  NAND2X0 U3757 ( .IN1(InstAddrPointer[29]), .IN2(n3327), .QN(n3350) );
  OA21X1 U3758 ( .IN1(InstAddrPointer[29]), .IN2(n4205), .IN3(n3328), .Q(n3351) );
  MUX21X1 U3759 ( .IN1(n3350), .IN2(n3351), .S(InstAddrPointer[30]), .Q(n3330)
         );
  NAND3X0 U3760 ( .IN1(n3331), .IN2(n3330), .IN3(n3329), .QN(n1991) );
  NAND2X0 U3761 ( .IN1(n3332), .IN2(InstAddrPointer[30]), .QN(n3333) );
  MUX21X1 U3762 ( .IN1(N3678), .IN2(n5224), .S(n3333), .Q(n3335) );
  XOR2X1 U3763 ( .IN1(n3334), .IN2(n3335), .Q(n4251) );
  OA22X1 U3764 ( .IN1(n3335), .IN2(n4206), .IN3(n4251), .IN4(n4208), .Q(n3349)
         );
  HADDX1 U3765 ( .A0(n3336), .B0(InstAddrPointer[30]), .C1(n3337), .SO(n3323)
         );
  XOR2X1 U3766 ( .IN1(n3337), .IN2(N3678), .Q(n3346) );
  HADDX1 U3767 ( .A0(n3338), .B0(InstAddrPointer[30]), .C1(n3339), .SO(n3298)
         );
  XOR2X1 U3768 ( .IN1(n3339), .IN2(N3678), .Q(n3340) );
  AO22X1 U3769 ( .IN1(n4132), .IN2(n3346), .IN3(n3340), .IN4(n2916), .Q(n3341)
         );
  XOR2X1 U3770 ( .IN1(n3341), .IN2(n3947), .Q(n3345) );
  FADDX1 U3771 ( .A(n3993), .B(n3343), .CI(n3342), .CO(n3344), .S(n3322) );
  XOR2X1 U3772 ( .IN1(n3345), .IN2(n3344), .Q(n4246) );
  NAND2X0 U3773 ( .IN1(n4246), .IN2(n4288), .QN(n3348) );
  NAND2X0 U3774 ( .IN1(n4290), .IN2(n3346), .QN(n3347) );
  AND3X1 U3775 ( .IN1(n3349), .IN2(n3348), .IN3(n3347), .Q(n3355) );
  NAND2X0 U3776 ( .IN1(n4104), .IN2(rEIP[31]), .QN(n4250) );
  OR3X1 U3777 ( .IN1(N3678), .IN2(n3350), .IN3(n5230), .Q(n3354) );
  OAI21X1 U3778 ( .IN1(n4205), .IN2(InstAddrPointer[30]), .IN3(n3351), .QN(
        n3352) );
  NAND2X0 U3779 ( .IN1(N3678), .IN2(n3352), .QN(n3353) );
  NAND4X0 U3780 ( .IN1(n3355), .IN2(n4250), .IN3(n3354), .IN4(n3353), .QN(
        n2070) );
  INVX0 U3781 ( .INP(n4266), .ZN(n4248) );
  OA22X1 U3782 ( .IN1(n4252), .IN2(n3357), .IN3(n3356), .IN4(n4248), .Q(n3358)
         );
  OA21X1 U3783 ( .IN1(n3359), .IN2(n5240), .IN3(n3358), .Q(n3364) );
  NAND2X0 U3784 ( .IN1(n4255), .IN2(n3368), .QN(n3362) );
  OR2X1 U3785 ( .IN1(PhyAddrPointer[29]), .IN2(n3360), .Q(n3361) );
  NAND4X0 U3786 ( .IN1(n3364), .IN2(n3363), .IN3(n3362), .IN4(n3361), .QN(
        n1707) );
  AOI22X1 U3787 ( .IN1(n4275), .IN2(EBX[29]), .IN3(n4274), .IN4(
        PhyAddrPointer[29]), .QN(n3372) );
  XOR2X1 U3788 ( .IN1(n3366), .IN2(n3365), .Q(n3367) );
  NAND2X0 U3789 ( .IN1(n4280), .IN2(n3367), .QN(n3371) );
  NAND2X0 U3790 ( .IN1(n2090), .IN2(n3368), .QN(n3370) );
  NAND2X0 U3791 ( .IN1(rEIP[29]), .IN2(n4281), .QN(n3369) );
  NAND4X0 U3792 ( .IN1(n3372), .IN2(n3371), .IN3(n3370), .IN4(n3369), .QN(
        n2036) );
  AOI22X1 U3793 ( .IN1(n4275), .IN2(EBX[27]), .IN3(n4274), .IN4(
        PhyAddrPointer[27]), .QN(n3379) );
  XOR2X1 U3794 ( .IN1(n3374), .IN2(n3373), .Q(n3375) );
  NAND2X0 U3795 ( .IN1(n4280), .IN2(n3375), .QN(n3378) );
  NAND2X0 U3796 ( .IN1(n2090), .IN2(n3385), .QN(n3377) );
  NAND2X0 U3797 ( .IN1(rEIP[27]), .IN2(n4281), .QN(n3376) );
  NAND4X0 U3798 ( .IN1(n3379), .IN2(n3378), .IN3(n3377), .IN4(n3376), .QN(
        n2038) );
  OAI21X1 U3799 ( .IN1(n3427), .IN2(n3642), .IN3(n3392), .QN(n3644) );
  FADDX1 U3800 ( .A(n3993), .B(n3381), .CI(n3380), .CO(n3393), .S(n3640) );
  INVX0 U3801 ( .INP(n3640), .ZN(n3382) );
  OA22X1 U3802 ( .IN1(n4252), .IN2(n3644), .IN3(n3382), .IN4(n4248), .Q(n3389)
         );
  NAND2X0 U3803 ( .IN1(n5098), .IN2(n3396), .QN(n3384) );
  OA21X1 U3804 ( .IN1(n3396), .IN2(n5020), .IN3(n4221), .Q(n3383) );
  MUX21X1 U3805 ( .IN1(n3384), .IN2(n3383), .S(PhyAddrPointer[27]), .Q(n3388)
         );
  NOR2X0 U3806 ( .IN1(n4147), .IN2(n5186), .QN(n3650) );
  INVX0 U3807 ( .INP(n3650), .ZN(n3387) );
  NAND2X0 U3808 ( .IN1(n4255), .IN2(n3385), .QN(n3386) );
  NAND4X0 U3809 ( .IN1(n3389), .IN2(n3388), .IN3(n3387), .IN4(n3386), .QN(
        n1709) );
  OA221X1 U3810 ( .IN1(n5020), .IN2(n3396), .IN3(n5020), .IN4(
        PhyAddrPointer[27]), .IN5(n4221), .Q(n3390) );
  NAND2X0 U3811 ( .IN1(n4104), .IN2(rEIP[28]), .QN(n3663) );
  OA21X1 U3812 ( .IN1(n3390), .IN2(n5243), .IN3(n3663), .Q(n3400) );
  AO21X1 U3813 ( .IN1(n3652), .IN2(n3392), .IN3(n3391), .Q(n3651) );
  FADDX1 U3814 ( .A(n3993), .B(n3394), .CI(n3393), .CO(n3299), .S(n3653) );
  INVX0 U3815 ( .INP(n3653), .ZN(n3395) );
  OA22X1 U3816 ( .IN1(n4252), .IN2(n3651), .IN3(n3395), .IN4(n4248), .Q(n3399)
         );
  NAND4X0 U3817 ( .IN1(PhyAddrPointer[27]), .IN2(n5098), .IN3(n3396), .IN4(
        n5243), .QN(n3398) );
  NAND2X0 U3818 ( .IN1(n4255), .IN2(n3404), .QN(n3397) );
  NAND4X0 U3819 ( .IN1(n3400), .IN2(n3399), .IN3(n3398), .IN4(n3397), .QN(
        n1708) );
  AOI22X1 U3820 ( .IN1(n4275), .IN2(EBX[28]), .IN3(n4274), .IN4(
        PhyAddrPointer[28]), .QN(n3408) );
  XOR2X1 U3821 ( .IN1(n3402), .IN2(n3401), .Q(n3403) );
  NAND2X0 U3822 ( .IN1(n4280), .IN2(n3403), .QN(n3407) );
  NAND2X0 U3823 ( .IN1(n2090), .IN2(n3404), .QN(n3406) );
  NAND2X0 U3824 ( .IN1(rEIP[28]), .IN2(n4281), .QN(n3405) );
  NAND4X0 U3825 ( .IN1(n3408), .IN2(n3407), .IN3(n3406), .IN4(n3405), .QN(
        n2037) );
  AOI22X1 U3826 ( .IN1(n4275), .IN2(EBX[25]), .IN3(n4274), .IN4(
        PhyAddrPointer[25]), .QN(n3415) );
  XOR2X1 U3827 ( .IN1(n3410), .IN2(n3409), .Q(n3411) );
  NAND2X0 U3828 ( .IN1(n4280), .IN2(n3411), .QN(n3414) );
  NAND2X0 U3829 ( .IN1(n2090), .IN2(n3421), .QN(n3413) );
  NAND2X0 U3830 ( .IN1(rEIP[25]), .IN2(n4281), .QN(n3412) );
  NAND4X0 U3831 ( .IN1(n3415), .IN2(n3414), .IN3(n3413), .IN4(n3412), .QN(
        n2040) );
  OAI21X1 U3832 ( .IN1(n3463), .IN2(n3617), .IN3(n3428), .QN(n3619) );
  FADDX1 U3833 ( .A(n3993), .B(n3417), .CI(n3416), .CO(n3429), .S(n3615) );
  INVX0 U3834 ( .INP(n3615), .ZN(n3418) );
  OA22X1 U3835 ( .IN1(n4252), .IN2(n3619), .IN3(n3418), .IN4(n4248), .Q(n3425)
         );
  NAND2X0 U3836 ( .IN1(n5098), .IN2(n3432), .QN(n3420) );
  OA21X1 U3837 ( .IN1(n3432), .IN2(n5020), .IN3(n4221), .Q(n3419) );
  MUX21X1 U3838 ( .IN1(n3420), .IN2(n3419), .S(PhyAddrPointer[25]), .Q(n3424)
         );
  NOR2X0 U3839 ( .IN1(n4147), .IN2(n5187), .QN(n3625) );
  INVX0 U3840 ( .INP(n3625), .ZN(n3423) );
  NAND2X0 U3841 ( .IN1(n4255), .IN2(n3421), .QN(n3422) );
  NAND4X0 U3842 ( .IN1(n3425), .IN2(n3424), .IN3(n3423), .IN4(n3422), .QN(
        n1711) );
  OA221X1 U3843 ( .IN1(n5020), .IN2(n3432), .IN3(n5020), .IN4(
        PhyAddrPointer[25]), .IN5(n4221), .Q(n3426) );
  NAND2X0 U3844 ( .IN1(n4104), .IN2(rEIP[26]), .QN(n3638) );
  OA21X1 U3845 ( .IN1(n3426), .IN2(n5244), .IN3(n3638), .Q(n3436) );
  AO21X1 U3846 ( .IN1(n3627), .IN2(n3428), .IN3(n3427), .Q(n3626) );
  FADDX1 U3847 ( .A(n3993), .B(n3430), .CI(n3429), .CO(n3380), .S(n3628) );
  INVX0 U3848 ( .INP(n3628), .ZN(n3431) );
  OA22X1 U3849 ( .IN1(n4252), .IN2(n3626), .IN3(n3431), .IN4(n4248), .Q(n3435)
         );
  NAND4X0 U3850 ( .IN1(PhyAddrPointer[25]), .IN2(n5098), .IN3(n3432), .IN4(
        n5244), .QN(n3434) );
  NAND2X0 U3851 ( .IN1(n4255), .IN2(n3440), .QN(n3433) );
  NAND4X0 U3852 ( .IN1(n3436), .IN2(n3435), .IN3(n3434), .IN4(n3433), .QN(
        n1710) );
  AOI22X1 U3853 ( .IN1(n4275), .IN2(EBX[26]), .IN3(n4274), .IN4(
        PhyAddrPointer[26]), .QN(n3444) );
  XOR2X1 U3854 ( .IN1(n3438), .IN2(n3437), .Q(n3439) );
  NAND2X0 U3855 ( .IN1(n4280), .IN2(n3439), .QN(n3443) );
  NAND2X0 U3856 ( .IN1(n2090), .IN2(n3440), .QN(n3442) );
  NAND2X0 U3857 ( .IN1(rEIP[26]), .IN2(n4281), .QN(n3441) );
  NAND4X0 U3858 ( .IN1(n3444), .IN2(n3443), .IN3(n3442), .IN4(n3441), .QN(
        n2039) );
  AOI22X1 U3859 ( .IN1(n4275), .IN2(EBX[23]), .IN3(n4274), .IN4(
        PhyAddrPointer[23]), .QN(n3451) );
  XOR2X1 U3860 ( .IN1(n3446), .IN2(n3445), .Q(n3447) );
  NAND2X0 U3861 ( .IN1(n4280), .IN2(n3447), .QN(n3450) );
  NAND2X0 U3862 ( .IN1(n2090), .IN2(n3457), .QN(n3449) );
  NAND2X0 U3863 ( .IN1(rEIP[23]), .IN2(n4281), .QN(n3448) );
  NAND4X0 U3864 ( .IN1(n3451), .IN2(n3450), .IN3(n3449), .IN4(n3448), .QN(
        n2042) );
  OAI21X1 U3865 ( .IN1(n3499), .IN2(n3592), .IN3(n3464), .QN(n3594) );
  FADDX1 U3866 ( .A(n3993), .B(n3453), .CI(n3452), .CO(n3465), .S(n3590) );
  INVX0 U3867 ( .INP(n3590), .ZN(n3454) );
  OA22X1 U3868 ( .IN1(n4252), .IN2(n3594), .IN3(n3454), .IN4(n4248), .Q(n3461)
         );
  NAND2X0 U3869 ( .IN1(n5098), .IN2(n3468), .QN(n3456) );
  OA21X1 U3870 ( .IN1(n3468), .IN2(n5020), .IN3(n4221), .Q(n3455) );
  MUX21X1 U3871 ( .IN1(n3456), .IN2(n3455), .S(PhyAddrPointer[23]), .Q(n3460)
         );
  NOR2X0 U3872 ( .IN1(n4147), .IN2(n5216), .QN(n3600) );
  INVX0 U3873 ( .INP(n3600), .ZN(n3459) );
  NAND2X0 U3874 ( .IN1(n4255), .IN2(n3457), .QN(n3458) );
  NAND4X0 U3875 ( .IN1(n3461), .IN2(n3460), .IN3(n3459), .IN4(n3458), .QN(
        n1713) );
  OA221X1 U3876 ( .IN1(n5020), .IN2(n3468), .IN3(n5020), .IN4(
        PhyAddrPointer[23]), .IN5(n4221), .Q(n3462) );
  NAND2X0 U3877 ( .IN1(n4104), .IN2(rEIP[24]), .QN(n3613) );
  OA21X1 U3878 ( .IN1(n3462), .IN2(n5245), .IN3(n3613), .Q(n3472) );
  AO21X1 U3879 ( .IN1(n3602), .IN2(n3464), .IN3(n3463), .Q(n3601) );
  FADDX1 U3880 ( .A(n3993), .B(n3466), .CI(n3465), .CO(n3416), .S(n3603) );
  INVX0 U3881 ( .INP(n3603), .ZN(n3467) );
  OA22X1 U3882 ( .IN1(n4252), .IN2(n3601), .IN3(n3467), .IN4(n4248), .Q(n3471)
         );
  NAND4X0 U3883 ( .IN1(PhyAddrPointer[23]), .IN2(n5098), .IN3(n3468), .IN4(
        n5245), .QN(n3470) );
  NAND2X0 U3884 ( .IN1(n4255), .IN2(n3476), .QN(n3469) );
  NAND4X0 U3885 ( .IN1(n3472), .IN2(n3471), .IN3(n3470), .IN4(n3469), .QN(
        n1712) );
  AOI22X1 U3886 ( .IN1(n4275), .IN2(EBX[24]), .IN3(n4274), .IN4(
        PhyAddrPointer[24]), .QN(n3480) );
  XOR2X1 U3887 ( .IN1(n3474), .IN2(n3473), .Q(n3475) );
  NAND2X0 U3888 ( .IN1(n4280), .IN2(n3475), .QN(n3479) );
  NAND2X0 U3889 ( .IN1(n2090), .IN2(n3476), .QN(n3478) );
  NAND2X0 U3890 ( .IN1(rEIP[24]), .IN2(n4281), .QN(n3477) );
  NAND4X0 U3891 ( .IN1(n3480), .IN2(n3479), .IN3(n3478), .IN4(n3477), .QN(
        n2041) );
  AOI22X1 U3892 ( .IN1(n4275), .IN2(EBX[21]), .IN3(n4274), .IN4(
        PhyAddrPointer[21]), .QN(n3487) );
  XOR2X1 U3893 ( .IN1(n3482), .IN2(n3481), .Q(n3483) );
  NAND2X0 U3894 ( .IN1(n4280), .IN2(n3483), .QN(n3486) );
  NAND2X0 U3895 ( .IN1(n2090), .IN2(n3493), .QN(n3485) );
  NAND2X0 U3896 ( .IN1(rEIP[21]), .IN2(n4281), .QN(n3484) );
  NAND4X0 U3897 ( .IN1(n3487), .IN2(n3486), .IN3(n3485), .IN4(n3484), .QN(
        n2044) );
  OAI21X1 U3898 ( .IN1(n3534), .IN2(n3567), .IN3(n3500), .QN(n3569) );
  FADDX1 U3899 ( .A(n3993), .B(n3489), .CI(n3488), .CO(n3501), .S(n3565) );
  INVX0 U3900 ( .INP(n3565), .ZN(n3490) );
  OA22X1 U3901 ( .IN1(n4252), .IN2(n3569), .IN3(n3490), .IN4(n4248), .Q(n3497)
         );
  NAND2X0 U3902 ( .IN1(n5098), .IN2(n3504), .QN(n3492) );
  INVX0 U3903 ( .INP(n5098), .ZN(n4222) );
  OA21X1 U3904 ( .IN1(n3504), .IN2(n4222), .IN3(n4221), .Q(n3491) );
  MUX21X1 U3905 ( .IN1(n3492), .IN2(n3491), .S(PhyAddrPointer[21]), .Q(n3496)
         );
  NOR2X0 U3906 ( .IN1(n4147), .IN2(n5188), .QN(n3575) );
  INVX0 U3907 ( .INP(n3575), .ZN(n3495) );
  NAND2X0 U3908 ( .IN1(n4255), .IN2(n3493), .QN(n3494) );
  NAND4X0 U3909 ( .IN1(n3497), .IN2(n3496), .IN3(n3495), .IN4(n3494), .QN(
        n1715) );
  OA221X1 U3910 ( .IN1(n5020), .IN2(n3504), .IN3(n5020), .IN4(
        PhyAddrPointer[21]), .IN5(n4221), .Q(n3498) );
  NAND2X0 U3911 ( .IN1(n4104), .IN2(rEIP[22]), .QN(n3588) );
  OA21X1 U3912 ( .IN1(n3498), .IN2(n5246), .IN3(n3588), .Q(n3508) );
  AO21X1 U3913 ( .IN1(n3577), .IN2(n3500), .IN3(n3499), .Q(n3576) );
  FADDX1 U3914 ( .A(n3993), .B(n3502), .CI(n3501), .CO(n3452), .S(n3578) );
  INVX0 U3915 ( .INP(n3578), .ZN(n3503) );
  OA22X1 U3916 ( .IN1(n4252), .IN2(n3576), .IN3(n3503), .IN4(n4248), .Q(n3507)
         );
  NAND4X0 U3917 ( .IN1(PhyAddrPointer[21]), .IN2(n5098), .IN3(n3504), .IN4(
        n5246), .QN(n3506) );
  NAND2X0 U3918 ( .IN1(n4255), .IN2(n3512), .QN(n3505) );
  NAND4X0 U3919 ( .IN1(n3508), .IN2(n3507), .IN3(n3506), .IN4(n3505), .QN(
        n1714) );
  AOI22X1 U3920 ( .IN1(n4275), .IN2(EBX[22]), .IN3(n4274), .IN4(
        PhyAddrPointer[22]), .QN(n3516) );
  XOR2X1 U3921 ( .IN1(n3510), .IN2(n3509), .Q(n3511) );
  NAND2X0 U3922 ( .IN1(n4280), .IN2(n3511), .QN(n3515) );
  NAND2X0 U3923 ( .IN1(n2090), .IN2(n3512), .QN(n3514) );
  NAND2X0 U3924 ( .IN1(rEIP[22]), .IN2(n4281), .QN(n3513) );
  NAND4X0 U3925 ( .IN1(n3516), .IN2(n3515), .IN3(n3514), .IN4(n3513), .QN(
        n2043) );
  NAND2X0 U3926 ( .IN1(rEIP[19]), .IN2(n4281), .QN(n3518) );
  NAND2X0 U3927 ( .IN1(n4275), .IN2(EBX[19]), .QN(n3517) );
  AND3X1 U3928 ( .IN1(n4147), .IN2(n3518), .IN3(n3517), .Q(n3525) );
  XOR2X1 U3929 ( .IN1(n3520), .IN2(n3519), .Q(n3521) );
  NAND2X0 U3930 ( .IN1(n4280), .IN2(n3521), .QN(n3524) );
  NAND2X0 U3931 ( .IN1(n2090), .IN2(n3530), .QN(n3523) );
  NAND2X0 U3932 ( .IN1(PhyAddrPointer[19]), .IN2(n4274), .QN(n3522) );
  NAND4X0 U3933 ( .IN1(n3525), .IN2(n3524), .IN3(n3523), .IN4(n3522), .QN(
        n2046) );
  FADDX1 U3934 ( .A(n3993), .B(n3527), .CI(n3526), .CO(n3536), .S(n3669) );
  OA21X1 U3935 ( .IN1(n3696), .IN2(n3677), .IN3(n3535), .Q(n3671) );
  INVX0 U3936 ( .INP(n4252), .ZN(n4262) );
  AOI22X1 U3937 ( .IN1(n3669), .IN2(n4266), .IN3(n3671), .IN4(n4262), .QN(
        n3533) );
  NAND2X0 U3938 ( .IN1(n5098), .IN2(n3541), .QN(n3529) );
  OA21X1 U3939 ( .IN1(n3541), .IN2(n4222), .IN3(n4221), .Q(n3528) );
  MUX21X1 U3940 ( .IN1(n3529), .IN2(n3528), .S(PhyAddrPointer[19]), .Q(n3532)
         );
  NAND2X0 U3941 ( .IN1(n4104), .IN2(rEIP[19]), .QN(n3673) );
  INVX0 U3942 ( .INP(n4431), .ZN(n4255) );
  NAND2X0 U3943 ( .IN1(n4255), .IN2(n3530), .QN(n3531) );
  NAND4X0 U3944 ( .IN1(n3533), .IN2(n3532), .IN3(n3673), .IN4(n3531), .QN(
        n1717) );
  OA221X1 U3945 ( .IN1(n5020), .IN2(n3541), .IN3(n5020), .IN4(
        PhyAddrPointer[19]), .IN5(n4221), .Q(n3540) );
  AO21X1 U3946 ( .IN1(n3557), .IN2(n3535), .IN3(n3534), .Q(n3556) );
  FADDX1 U3947 ( .A(n3993), .B(n3537), .CI(n3536), .CO(n3488), .S(n3538) );
  INVX0 U3948 ( .INP(n3538), .ZN(n3554) );
  OA22X1 U3949 ( .IN1(n4252), .IN2(n3556), .IN3(n3554), .IN4(n4248), .Q(n3539)
         );
  OA21X1 U3950 ( .IN1(n3540), .IN2(n5247), .IN3(n3539), .Q(n3544) );
  NAND4X0 U3951 ( .IN1(PhyAddrPointer[19]), .IN2(n5098), .IN3(n3541), .IN4(
        n5247), .QN(n3543) );
  NAND2X0 U3952 ( .IN1(n4104), .IN2(rEIP[20]), .QN(n3555) );
  NAND2X0 U3953 ( .IN1(n4255), .IN2(n3548), .QN(n3542) );
  NAND4X0 U3954 ( .IN1(n3544), .IN2(n3543), .IN3(n3555), .IN4(n3542), .QN(
        n1716) );
  AOI22X1 U3955 ( .IN1(n4275), .IN2(EBX[20]), .IN3(n4274), .IN4(
        PhyAddrPointer[20]), .QN(n3552) );
  XOR2X1 U3956 ( .IN1(n3546), .IN2(n3545), .Q(n3547) );
  NAND2X0 U3957 ( .IN1(n4280), .IN2(n3547), .QN(n3551) );
  NAND2X0 U3958 ( .IN1(n2090), .IN2(n3548), .QN(n3550) );
  NAND2X0 U3959 ( .IN1(rEIP[20]), .IN2(n4281), .QN(n3549) );
  NAND4X0 U3960 ( .IN1(n3552), .IN2(n3551), .IN3(n3550), .IN4(n3549), .QN(
        n2045) );
  NOR2X0 U3961 ( .IN1(InstAddrPointer[19]), .IN2(n4205), .QN(n3667) );
  AO21X1 U3962 ( .IN1(n4236), .IN2(n3665), .IN3(n4217), .Q(n3670) );
  NOR2X0 U3963 ( .IN1(n3667), .IN2(n3670), .QN(n3553) );
  OA22X1 U3964 ( .IN1(n4060), .IN2(n3554), .IN3(n3553), .IN4(n5215), .Q(n3564)
         );
  OA21X1 U3965 ( .IN1(n4208), .IN2(n3556), .IN3(n3555), .Q(n3563) );
  NOR2X0 U3966 ( .IN1(n3557), .IN2(n4206), .QN(n3558) );
  AOI21X1 U3967 ( .IN1(n4290), .IN2(n3559), .IN3(n3558), .QN(n3562) );
  NAND3X0 U3968 ( .IN1(n4236), .IN2(n3560), .IN3(n5215), .QN(n3561) );
  NAND4X0 U3969 ( .IN1(n3564), .IN2(n3563), .IN3(n3562), .IN4(n3561), .QN(
        n2001) );
  AO21X1 U3970 ( .IN1(n4236), .IN2(n3566), .IN3(n4217), .Q(n3584) );
  AO22X1 U3971 ( .IN1(n3584), .IN2(InstAddrPointer[21]), .IN3(n3565), .IN4(
        n4288), .Q(n3574) );
  INVX0 U3972 ( .INP(n3566), .ZN(n3568) );
  NOR2X0 U3973 ( .IN1(InstAddrPointer[21]), .IN2(n4205), .QN(n3585) );
  AO22X1 U3974 ( .IN1(n3568), .IN2(n3585), .IN3(n3567), .IN4(n4237), .Q(n3573)
         );
  NOR2X0 U3975 ( .IN1(n4208), .IN2(n3569), .QN(n3570) );
  AO21X1 U3976 ( .IN1(n4290), .IN2(n3571), .IN3(n3570), .Q(n3572) );
  OR4X1 U3977 ( .IN1(n3575), .IN2(n3574), .IN3(n3573), .IN4(n3572), .Q(n2000)
         );
  OA22X1 U3978 ( .IN1(n3577), .IN2(n4206), .IN3(n4208), .IN4(n3576), .Q(n3582)
         );
  NAND2X0 U3979 ( .IN1(n3578), .IN2(n4288), .QN(n3581) );
  NAND2X0 U3980 ( .IN1(n4290), .IN2(n3579), .QN(n3580) );
  AND3X1 U3981 ( .IN1(n3582), .IN2(n3581), .IN3(n3580), .Q(n3589) );
  NAND3X0 U3982 ( .IN1(n4236), .IN2(n3583), .IN3(n5231), .QN(n3587) );
  OAI21X1 U3983 ( .IN1(n3585), .IN2(n3584), .IN3(InstAddrPointer[22]), .QN(
        n3586) );
  NAND4X0 U3984 ( .IN1(n3589), .IN2(n3588), .IN3(n3587), .IN4(n3586), .QN(
        n1999) );
  AO21X1 U3985 ( .IN1(n4236), .IN2(n3591), .IN3(n4217), .Q(n3609) );
  AO22X1 U3986 ( .IN1(n3609), .IN2(InstAddrPointer[23]), .IN3(n3590), .IN4(
        n4288), .Q(n3599) );
  INVX0 U3987 ( .INP(n3591), .ZN(n3593) );
  NOR2X0 U3988 ( .IN1(n4205), .IN2(InstAddrPointer[23]), .QN(n3610) );
  AO22X1 U3989 ( .IN1(n3593), .IN2(n3610), .IN3(n3592), .IN4(n4237), .Q(n3598)
         );
  NOR2X0 U3990 ( .IN1(n4208), .IN2(n3594), .QN(n3595) );
  AO21X1 U3991 ( .IN1(n4290), .IN2(n3596), .IN3(n3595), .Q(n3597) );
  OR4X1 U3992 ( .IN1(n3600), .IN2(n3599), .IN3(n3598), .IN4(n3597), .Q(n1998)
         );
  OA22X1 U3993 ( .IN1(n3602), .IN2(n4206), .IN3(n4208), .IN4(n3601), .Q(n3607)
         );
  NAND2X0 U3994 ( .IN1(n3603), .IN2(n4288), .QN(n3606) );
  NAND2X0 U3995 ( .IN1(n4290), .IN2(n3604), .QN(n3605) );
  AND3X1 U3996 ( .IN1(n3607), .IN2(n3606), .IN3(n3605), .Q(n3614) );
  NAND3X0 U3997 ( .IN1(n4236), .IN2(n3608), .IN3(n5232), .QN(n3612) );
  OAI21X1 U3998 ( .IN1(n3610), .IN2(n3609), .IN3(InstAddrPointer[24]), .QN(
        n3611) );
  NAND4X0 U3999 ( .IN1(n3614), .IN2(n3613), .IN3(n3612), .IN4(n3611), .QN(
        n1997) );
  AO21X1 U4000 ( .IN1(n4236), .IN2(n3616), .IN3(n4217), .Q(n3634) );
  AO22X1 U4001 ( .IN1(n3634), .IN2(InstAddrPointer[25]), .IN3(n3615), .IN4(
        n4288), .Q(n3624) );
  INVX0 U4002 ( .INP(n3616), .ZN(n3618) );
  NOR2X0 U4003 ( .IN1(n4205), .IN2(InstAddrPointer[25]), .QN(n3635) );
  AO22X1 U4004 ( .IN1(n3618), .IN2(n3635), .IN3(n3617), .IN4(n4237), .Q(n3623)
         );
  NOR2X0 U4005 ( .IN1(n4208), .IN2(n3619), .QN(n3620) );
  AO21X1 U4006 ( .IN1(n4290), .IN2(n3621), .IN3(n3620), .Q(n3622) );
  OR4X1 U4007 ( .IN1(n3625), .IN2(n3624), .IN3(n3623), .IN4(n3622), .Q(n1996)
         );
  OA22X1 U4008 ( .IN1(n3627), .IN2(n4206), .IN3(n4208), .IN4(n3626), .Q(n3632)
         );
  NAND2X0 U4009 ( .IN1(n3628), .IN2(n4288), .QN(n3631) );
  NAND2X0 U4010 ( .IN1(n4290), .IN2(n3629), .QN(n3630) );
  AND3X1 U4011 ( .IN1(n3632), .IN2(n3631), .IN3(n3630), .Q(n3639) );
  NAND3X0 U4012 ( .IN1(n4236), .IN2(n3633), .IN3(n5233), .QN(n3637) );
  OAI21X1 U4013 ( .IN1(n3635), .IN2(n3634), .IN3(InstAddrPointer[26]), .QN(
        n3636) );
  NAND4X0 U4014 ( .IN1(n3639), .IN2(n3638), .IN3(n3637), .IN4(n3636), .QN(
        n1995) );
  AO21X1 U4015 ( .IN1(n4236), .IN2(n3641), .IN3(n4217), .Q(n3659) );
  AO22X1 U4016 ( .IN1(n3659), .IN2(InstAddrPointer[27]), .IN3(n3640), .IN4(
        n4288), .Q(n3649) );
  INVX0 U4017 ( .INP(n3641), .ZN(n3643) );
  NOR2X0 U4018 ( .IN1(n4205), .IN2(InstAddrPointer[27]), .QN(n3660) );
  AO22X1 U4019 ( .IN1(n3643), .IN2(n3660), .IN3(n3642), .IN4(n4237), .Q(n3648)
         );
  NOR2X0 U4020 ( .IN1(n4208), .IN2(n3644), .QN(n3645) );
  AO21X1 U4021 ( .IN1(n4290), .IN2(n3646), .IN3(n3645), .Q(n3647) );
  OR4X1 U4022 ( .IN1(n3650), .IN2(n3649), .IN3(n3648), .IN4(n3647), .Q(n1994)
         );
  OA22X1 U4023 ( .IN1(n3652), .IN2(n4206), .IN3(n4208), .IN4(n3651), .Q(n3657)
         );
  NAND2X0 U4024 ( .IN1(n3653), .IN2(n4288), .QN(n3656) );
  NAND2X0 U4025 ( .IN1(n4290), .IN2(n3654), .QN(n3655) );
  AND3X1 U4026 ( .IN1(n3657), .IN2(n3656), .IN3(n3655), .Q(n3664) );
  NAND3X0 U4027 ( .IN1(n4236), .IN2(n3658), .IN3(n5237), .QN(n3662) );
  OAI21X1 U4028 ( .IN1(n3660), .IN2(n3659), .IN3(InstAddrPointer[28]), .QN(
        n3661) );
  NAND4X0 U4029 ( .IN1(n3664), .IN2(n3663), .IN3(n3662), .IN4(n3661), .QN(
        n1993) );
  INVX0 U4030 ( .INP(n3665), .ZN(n3666) );
  AOI22X1 U4031 ( .IN1(n4290), .IN2(n3668), .IN3(n3667), .IN4(n3666), .QN(
        n3675) );
  AOI22X1 U4032 ( .IN1(n3670), .IN2(InstAddrPointer[19]), .IN3(n3669), .IN4(
        n4288), .QN(n3674) );
  INVX0 U4033 ( .INP(n4208), .ZN(n4287) );
  NAND2X0 U4034 ( .IN1(n3671), .IN2(n4287), .QN(n3672) );
  NAND4X0 U4035 ( .IN1(n3675), .IN2(n3674), .IN3(n3673), .IN4(n3672), .QN(
        n3676) );
  AO21X1 U4036 ( .IN1(n4237), .IN2(n3677), .IN3(n3676), .Q(n2002) );
  NAND2X0 U4037 ( .IN1(rEIP[17]), .IN2(n4281), .QN(n3679) );
  NAND2X0 U4038 ( .IN1(n4275), .IN2(EBX[17]), .QN(n3678) );
  AND3X1 U4039 ( .IN1(n4147), .IN2(n3679), .IN3(n3678), .Q(n3686) );
  XOR2X1 U4040 ( .IN1(n3681), .IN2(n3680), .Q(n3682) );
  NAND2X0 U4041 ( .IN1(n4280), .IN2(n3682), .QN(n3685) );
  NAND2X0 U4042 ( .IN1(n2090), .IN2(n3692), .QN(n3684) );
  NAND2X0 U4043 ( .IN1(PhyAddrPointer[17]), .IN2(n4274), .QN(n3683) );
  NAND4X0 U4044 ( .IN1(n3686), .IN2(n3685), .IN3(n3684), .IN4(n3683), .QN(
        n2048) );
  OA21X1 U4045 ( .IN1(n3703), .IN2(n4222), .IN3(n4221), .Q(n3690) );
  FADDX1 U4046 ( .A(n3993), .B(n3688), .CI(n3687), .CO(n3698), .S(n3728) );
  INVX0 U4047 ( .INP(n3728), .ZN(n3689) );
  OA22X1 U4048 ( .IN1(n3690), .IN2(n5241), .IN3(n4248), .IN4(n3689), .Q(n3695)
         );
  AND2X1 U4049 ( .IN1(n5098), .IN2(n3703), .Q(n3691) );
  OA21X1 U4050 ( .IN1(n3759), .IN2(n3736), .IN3(n3697), .Q(n3733) );
  AOI22X1 U4051 ( .IN1(n3691), .IN2(n5241), .IN3(n3733), .IN4(n4262), .QN(
        n3694) );
  NAND2X0 U4052 ( .IN1(n4104), .IN2(rEIP[17]), .QN(n3737) );
  NAND2X0 U4053 ( .IN1(n4255), .IN2(n3692), .QN(n3693) );
  NAND4X0 U4054 ( .IN1(n3695), .IN2(n3694), .IN3(n3737), .IN4(n3693), .QN(
        n1719) );
  OA221X1 U4055 ( .IN1(n5020), .IN2(n3703), .IN3(n5020), .IN4(
        PhyAddrPointer[17]), .IN5(n4221), .Q(n3702) );
  AO21X1 U4056 ( .IN1(n3722), .IN2(n3697), .IN3(n3696), .Q(n3721) );
  FADDX1 U4057 ( .A(n3993), .B(n3699), .CI(n3698), .CO(n3526), .S(n3700) );
  INVX0 U4058 ( .INP(n3700), .ZN(n3719) );
  OA22X1 U4059 ( .IN1(n4252), .IN2(n3721), .IN3(n3719), .IN4(n4248), .Q(n3701)
         );
  OA21X1 U4060 ( .IN1(n3702), .IN2(n5191), .IN3(n3701), .Q(n3706) );
  NAND2X0 U4061 ( .IN1(n4104), .IN2(rEIP[18]), .QN(n3718) );
  NAND4X0 U4062 ( .IN1(PhyAddrPointer[17]), .IN2(n5098), .IN3(n3703), .IN4(
        n5191), .QN(n3705) );
  NAND2X0 U4063 ( .IN1(n4255), .IN2(n3709), .QN(n3704) );
  NAND4X0 U4064 ( .IN1(n3706), .IN2(n3718), .IN3(n3705), .IN4(n3704), .QN(
        n1718) );
  XOR2X1 U4065 ( .IN1(n3708), .IN2(n3707), .Q(n3714) );
  OA22X1 U4066 ( .IN1(n4280), .IN2(n5254), .IN3(n5191), .IN4(n3288), .Q(n3712)
         );
  NAND2X0 U4067 ( .IN1(n2090), .IN2(n3709), .QN(n3711) );
  NAND2X0 U4068 ( .IN1(n4275), .IN2(EBX[18]), .QN(n3710) );
  NAND4X0 U4069 ( .IN1(n3712), .IN2(n4147), .IN3(n3711), .IN4(n3710), .QN(
        n3713) );
  AO21X1 U4070 ( .IN1(n4280), .IN2(n3714), .IN3(n3713), .Q(n2047) );
  NOR2X0 U4071 ( .IN1(InstAddrPointer[17]), .IN2(n4205), .QN(n3731) );
  AO21X1 U4072 ( .IN1(n4236), .IN2(n3730), .IN3(n4217), .Q(n3729) );
  NOR2X0 U4073 ( .IN1(n3731), .IN2(n3729), .QN(n3717) );
  NAND2X0 U4074 ( .IN1(n4290), .IN2(n3715), .QN(n3716) );
  OA21X1 U4075 ( .IN1(n3717), .IN2(n5238), .IN3(n3716), .Q(n3727) );
  OA21X1 U4076 ( .IN1(n4060), .IN2(n3719), .IN3(n3718), .Q(n3720) );
  OA21X1 U4077 ( .IN1(n4208), .IN2(n3721), .IN3(n3720), .Q(n3726) );
  OR2X1 U4078 ( .IN1(n4206), .IN2(n3722), .Q(n3725) );
  NAND3X0 U4079 ( .IN1(n4236), .IN2(n3723), .IN3(n5238), .QN(n3724) );
  NAND4X0 U4080 ( .IN1(n3727), .IN2(n3726), .IN3(n3725), .IN4(n3724), .QN(
        n2003) );
  AOI22X1 U4081 ( .IN1(n3729), .IN2(InstAddrPointer[17]), .IN3(n3728), .IN4(
        n4288), .QN(n3740) );
  INVX0 U4082 ( .INP(n3730), .ZN(n3732) );
  AO22X1 U4083 ( .IN1(n4287), .IN2(n3733), .IN3(n3732), .IN4(n3731), .Q(n3734)
         );
  AOI21X1 U4084 ( .IN1(n4290), .IN2(n3735), .IN3(n3734), .QN(n3739) );
  NAND2X0 U4085 ( .IN1(n4237), .IN2(n3736), .QN(n3738) );
  NAND4X0 U4086 ( .IN1(n3740), .IN2(n3739), .IN3(n3738), .IN4(n3737), .QN(
        n2004) );
  NAND2X0 U4087 ( .IN1(rEIP[15]), .IN2(n4281), .QN(n3742) );
  NAND2X0 U4088 ( .IN1(n4275), .IN2(EBX[15]), .QN(n3741) );
  AND3X1 U4089 ( .IN1(n4147), .IN2(n3742), .IN3(n3741), .Q(n3749) );
  XOR2X1 U4090 ( .IN1(n3744), .IN2(n3743), .Q(n3745) );
  NAND2X0 U4091 ( .IN1(n4280), .IN2(n3745), .QN(n3748) );
  NAND2X0 U4092 ( .IN1(n2090), .IN2(n3754), .QN(n3747) );
  NAND2X0 U4093 ( .IN1(PhyAddrPointer[15]), .IN2(n4274), .QN(n3746) );
  NAND4X0 U4094 ( .IN1(n3749), .IN2(n3748), .IN3(n3747), .IN4(n3746), .QN(
        n2050) );
  FADDX1 U4095 ( .A(n3993), .B(n3751), .CI(n3750), .CO(n3761), .S(n3795) );
  OA21X1 U4096 ( .IN1(n3819), .IN2(n3792), .IN3(n3760), .Q(n3797) );
  AOI22X1 U4097 ( .IN1(n3795), .IN2(n4266), .IN3(n3797), .IN4(n4262), .QN(
        n3757) );
  NAND2X0 U4098 ( .IN1(n5098), .IN2(n3764), .QN(n3753) );
  OA21X1 U4099 ( .IN1(n3764), .IN2(n4222), .IN3(n4221), .Q(n3752) );
  MUX21X1 U4100 ( .IN1(n3753), .IN2(n3752), .S(PhyAddrPointer[15]), .Q(n3756)
         );
  NAND2X0 U4101 ( .IN1(n4104), .IN2(rEIP[15]), .QN(n3799) );
  NAND2X0 U4102 ( .IN1(n4255), .IN2(n3754), .QN(n3755) );
  NAND4X0 U4103 ( .IN1(n3757), .IN2(n3756), .IN3(n3799), .IN4(n3755), .QN(
        n1721) );
  OA221X1 U4104 ( .IN1(n5020), .IN2(n3764), .IN3(n5020), .IN4(
        PhyAddrPointer[15]), .IN5(n4221), .Q(n3758) );
  NAND2X0 U4105 ( .IN1(n4104), .IN2(rEIP[16]), .QN(n3786) );
  OA21X1 U4106 ( .IN1(n3758), .IN2(n5192), .IN3(n3786), .Q(n3768) );
  AO21X1 U4107 ( .IN1(n3778), .IN2(n3760), .IN3(n3759), .Q(n3777) );
  FADDX1 U4108 ( .A(n3993), .B(n3762), .CI(n3761), .CO(n3687), .S(n3763) );
  INVX0 U4109 ( .INP(n3763), .ZN(n3785) );
  OA22X1 U4110 ( .IN1(n4252), .IN2(n3777), .IN3(n3785), .IN4(n4248), .Q(n3767)
         );
  NAND4X0 U4111 ( .IN1(PhyAddrPointer[15]), .IN2(n5098), .IN3(n3764), .IN4(
        n5192), .QN(n3766) );
  NAND2X0 U4112 ( .IN1(n4255), .IN2(n3771), .QN(n3765) );
  NAND4X0 U4113 ( .IN1(n3768), .IN2(n3767), .IN3(n3766), .IN4(n3765), .QN(
        n1720) );
  XOR2X1 U4114 ( .IN1(n3770), .IN2(n3769), .Q(n3776) );
  OA22X1 U4115 ( .IN1(n4280), .IN2(n5255), .IN3(n5192), .IN4(n3288), .Q(n3774)
         );
  NAND2X0 U4116 ( .IN1(n2090), .IN2(n3771), .QN(n3773) );
  NAND2X0 U4117 ( .IN1(n4275), .IN2(EBX[16]), .QN(n3772) );
  NAND4X0 U4118 ( .IN1(n3774), .IN2(n4147), .IN3(n3773), .IN4(n3772), .QN(
        n3775) );
  AO21X1 U4119 ( .IN1(n4280), .IN2(n3776), .IN3(n3775), .Q(n2049) );
  OA22X1 U4120 ( .IN1(n3778), .IN2(n4206), .IN3(n4208), .IN4(n3777), .Q(n3783)
         );
  NAND3X0 U4121 ( .IN1(n4236), .IN2(n3779), .IN3(n5226), .QN(n3782) );
  NAND2X0 U4122 ( .IN1(n4290), .IN2(n3780), .QN(n3781) );
  AND3X1 U4123 ( .IN1(n3783), .IN2(n3782), .IN3(n3781), .Q(n3788) );
  AO21X1 U4124 ( .IN1(n4236), .IN2(n3789), .IN3(n4217), .Q(n3796) );
  NOR2X0 U4125 ( .IN1(InstAddrPointer[15]), .IN2(n4205), .QN(n3790) );
  NOR2X0 U4126 ( .IN1(n3796), .IN2(n3790), .QN(n3784) );
  OA22X1 U4127 ( .IN1(n4060), .IN2(n3785), .IN3(n3784), .IN4(n5226), .Q(n3787)
         );
  NAND3X0 U4128 ( .IN1(n3788), .IN2(n3787), .IN3(n3786), .QN(n2005) );
  INVX0 U4129 ( .INP(n3789), .ZN(n3791) );
  AO22X1 U4130 ( .IN1(n3792), .IN2(n4237), .IN3(n3791), .IN4(n3790), .Q(n3793)
         );
  AOI21X1 U4131 ( .IN1(n4290), .IN2(n3794), .IN3(n3793), .QN(n3801) );
  AOI22X1 U4132 ( .IN1(InstAddrPointer[15]), .IN2(n3796), .IN3(n3795), .IN4(
        n4288), .QN(n3800) );
  NAND2X0 U4133 ( .IN1(n3797), .IN2(n4287), .QN(n3798) );
  NAND4X0 U4134 ( .IN1(n3801), .IN2(n3800), .IN3(n3799), .IN4(n3798), .QN(
        n2006) );
  NAND2X0 U4135 ( .IN1(rEIP[13]), .IN2(n4281), .QN(n3803) );
  NAND2X0 U4136 ( .IN1(n4275), .IN2(EBX[13]), .QN(n3802) );
  AND3X1 U4137 ( .IN1(n4147), .IN2(n3803), .IN3(n3802), .Q(n3810) );
  XOR2X1 U4138 ( .IN1(n3805), .IN2(n3804), .Q(n3806) );
  NAND2X0 U4139 ( .IN1(n4280), .IN2(n3806), .QN(n3809) );
  NAND2X0 U4140 ( .IN1(n2090), .IN2(n3815), .QN(n3808) );
  NAND2X0 U4141 ( .IN1(PhyAddrPointer[13]), .IN2(n4274), .QN(n3807) );
  NAND4X0 U4142 ( .IN1(n3810), .IN2(n3809), .IN3(n3808), .IN4(n3807), .QN(
        n2052) );
  FADDX1 U4143 ( .A(n3947), .B(n3812), .CI(n3811), .CO(n3821), .S(n3857) );
  OA21X1 U4144 ( .IN1(n3881), .IN2(n3854), .IN3(n3820), .Q(n3859) );
  AOI22X1 U4145 ( .IN1(n3857), .IN2(n4266), .IN3(n3859), .IN4(n4262), .QN(
        n3818) );
  AND2X1 U4146 ( .IN1(n5098), .IN2(n3813), .Q(n3826) );
  INVX0 U4147 ( .INP(n3826), .ZN(n3814) );
  OA21X1 U4148 ( .IN1(n3813), .IN2(n4222), .IN3(n4221), .Q(n3824) );
  MUX21X1 U4149 ( .IN1(n3814), .IN2(n3824), .S(PhyAddrPointer[13]), .Q(n3817)
         );
  NAND2X0 U4150 ( .IN1(n4104), .IN2(rEIP[13]), .QN(n3861) );
  NAND2X0 U4151 ( .IN1(n4255), .IN2(n3815), .QN(n3816) );
  NAND4X0 U4152 ( .IN1(n3818), .IN2(n3817), .IN3(n3861), .IN4(n3816), .QN(
        n1723) );
  AO21X1 U4153 ( .IN1(n3840), .IN2(n3820), .IN3(n3819), .Q(n3839) );
  FADDX1 U4154 ( .A(n3947), .B(n3822), .CI(n3821), .CO(n3750), .S(n3823) );
  INVX0 U4155 ( .INP(n3823), .ZN(n3847) );
  OA22X1 U4156 ( .IN1(n4252), .IN2(n3839), .IN3(n3847), .IN4(n4248), .Q(n3830)
         );
  OA21X1 U4157 ( .IN1(PhyAddrPointer[13]), .IN2(n5020), .IN3(n3824), .Q(n3825)
         );
  NAND2X0 U4158 ( .IN1(n4104), .IN2(rEIP[14]), .QN(n3848) );
  OA21X1 U4159 ( .IN1(n3825), .IN2(n5193), .IN3(n3848), .Q(n3829) );
  NAND3X0 U4160 ( .IN1(PhyAddrPointer[13]), .IN2(n3826), .IN3(n5193), .QN(
        n3828) );
  NAND2X0 U4161 ( .IN1(n4255), .IN2(n3833), .QN(n3827) );
  NAND4X0 U4162 ( .IN1(n3830), .IN2(n3829), .IN3(n3828), .IN4(n3827), .QN(
        n1722) );
  XOR2X1 U4163 ( .IN1(n3832), .IN2(n3831), .Q(n3838) );
  OA22X1 U4164 ( .IN1(n4280), .IN2(n5256), .IN3(n5193), .IN4(n3288), .Q(n3836)
         );
  NAND2X0 U4165 ( .IN1(n2090), .IN2(n3833), .QN(n3835) );
  NAND2X0 U4166 ( .IN1(n4275), .IN2(EBX[14]), .QN(n3834) );
  NAND4X0 U4167 ( .IN1(n3836), .IN2(n4147), .IN3(n3835), .IN4(n3834), .QN(
        n3837) );
  AO21X1 U4168 ( .IN1(n4280), .IN2(n3838), .IN3(n3837), .Q(n2051) );
  OA22X1 U4169 ( .IN1(n3840), .IN2(n4206), .IN3(n4208), .IN4(n3839), .Q(n3845)
         );
  NAND3X0 U4170 ( .IN1(n4236), .IN2(n3841), .IN3(n5227), .QN(n3844) );
  NAND2X0 U4171 ( .IN1(n4290), .IN2(n3842), .QN(n3843) );
  AND3X1 U4172 ( .IN1(n3845), .IN2(n3844), .IN3(n3843), .Q(n3850) );
  AO21X1 U4173 ( .IN1(n4236), .IN2(n3851), .IN3(n4217), .Q(n3858) );
  NOR2X0 U4174 ( .IN1(InstAddrPointer[13]), .IN2(n4205), .QN(n3852) );
  NOR2X0 U4175 ( .IN1(n3858), .IN2(n3852), .QN(n3846) );
  OA22X1 U4176 ( .IN1(n4060), .IN2(n3847), .IN3(n3846), .IN4(n5227), .Q(n3849)
         );
  NAND3X0 U4177 ( .IN1(n3850), .IN2(n3849), .IN3(n3848), .QN(n2007) );
  INVX0 U4178 ( .INP(n3851), .ZN(n3853) );
  AO22X1 U4179 ( .IN1(n3854), .IN2(n4237), .IN3(n3853), .IN4(n3852), .Q(n3855)
         );
  AOI21X1 U4180 ( .IN1(n4290), .IN2(n3856), .IN3(n3855), .QN(n3863) );
  AOI22X1 U4181 ( .IN1(InstAddrPointer[13]), .IN2(n3858), .IN3(n3857), .IN4(
        n4288), .QN(n3862) );
  NAND2X0 U4182 ( .IN1(n3859), .IN2(n4287), .QN(n3860) );
  NAND4X0 U4183 ( .IN1(n3863), .IN2(n3862), .IN3(n3861), .IN4(n3860), .QN(
        n2008) );
  NAND2X0 U4184 ( .IN1(rEIP[11]), .IN2(n4281), .QN(n3865) );
  NAND2X0 U4185 ( .IN1(n4275), .IN2(EBX[11]), .QN(n3864) );
  AND3X1 U4186 ( .IN1(n4147), .IN2(n3865), .IN3(n3864), .Q(n3872) );
  XOR2X1 U4187 ( .IN1(n3867), .IN2(n3866), .Q(n3868) );
  NAND2X0 U4188 ( .IN1(n4280), .IN2(n3868), .QN(n3871) );
  NAND2X0 U4189 ( .IN1(n2090), .IN2(n3877), .QN(n3870) );
  NAND2X0 U4190 ( .IN1(PhyAddrPointer[11]), .IN2(n4274), .QN(n3869) );
  NAND4X0 U4191 ( .IN1(n3872), .IN2(n3871), .IN3(n3870), .IN4(n3869), .QN(
        n2054) );
  FADDX1 U4192 ( .A(n3947), .B(n3874), .CI(n3873), .CO(n3883), .S(n3919) );
  OA21X1 U4193 ( .IN1(n3943), .IN2(n3916), .IN3(n3882), .Q(n3921) );
  AOI22X1 U4194 ( .IN1(n3919), .IN2(n4266), .IN3(n3921), .IN4(n4262), .QN(
        n3880) );
  AND2X1 U4195 ( .IN1(n5098), .IN2(n3875), .Q(n3888) );
  INVX0 U4196 ( .INP(n3888), .ZN(n3876) );
  OA21X1 U4197 ( .IN1(n3875), .IN2(n4222), .IN3(n4221), .Q(n3886) );
  MUX21X1 U4198 ( .IN1(n3876), .IN2(n3886), .S(PhyAddrPointer[11]), .Q(n3879)
         );
  NAND2X0 U4199 ( .IN1(n4104), .IN2(rEIP[11]), .QN(n3923) );
  NAND2X0 U4200 ( .IN1(n4255), .IN2(n3877), .QN(n3878) );
  NAND4X0 U4201 ( .IN1(n3880), .IN2(n3879), .IN3(n3923), .IN4(n3878), .QN(
        n1725) );
  AO21X1 U4202 ( .IN1(n3902), .IN2(n3882), .IN3(n3881), .Q(n3901) );
  FADDX1 U4203 ( .A(n3947), .B(n3884), .CI(n3883), .CO(n3811), .S(n3885) );
  INVX0 U4204 ( .INP(n3885), .ZN(n3909) );
  OA22X1 U4205 ( .IN1(n4252), .IN2(n3901), .IN3(n3909), .IN4(n4248), .Q(n3892)
         );
  OA21X1 U4206 ( .IN1(PhyAddrPointer[11]), .IN2(n5020), .IN3(n3886), .Q(n3887)
         );
  NAND2X0 U4207 ( .IN1(n4104), .IN2(rEIP[12]), .QN(n3910) );
  OA21X1 U4208 ( .IN1(n3887), .IN2(n5194), .IN3(n3910), .Q(n3891) );
  NAND3X0 U4209 ( .IN1(PhyAddrPointer[11]), .IN2(n3888), .IN3(n5194), .QN(
        n3890) );
  NAND2X0 U4210 ( .IN1(n4255), .IN2(n3895), .QN(n3889) );
  NAND4X0 U4211 ( .IN1(n3892), .IN2(n3891), .IN3(n3890), .IN4(n3889), .QN(
        n1724) );
  XOR2X1 U4212 ( .IN1(n3894), .IN2(n3893), .Q(n3900) );
  OA22X1 U4213 ( .IN1(n4280), .IN2(n5257), .IN3(n5194), .IN4(n3288), .Q(n3898)
         );
  NAND2X0 U4214 ( .IN1(n2090), .IN2(n3895), .QN(n3897) );
  NAND2X0 U4215 ( .IN1(n4275), .IN2(EBX[12]), .QN(n3896) );
  NAND4X0 U4216 ( .IN1(n3898), .IN2(n4147), .IN3(n3897), .IN4(n3896), .QN(
        n3899) );
  AO21X1 U4217 ( .IN1(n4280), .IN2(n3900), .IN3(n3899), .Q(n2053) );
  OA22X1 U4218 ( .IN1(n3902), .IN2(n4206), .IN3(n4208), .IN4(n3901), .Q(n3907)
         );
  NAND3X0 U4219 ( .IN1(n4236), .IN2(n3903), .IN3(n5228), .QN(n3906) );
  NAND2X0 U4220 ( .IN1(n4290), .IN2(n3904), .QN(n3905) );
  AND3X1 U4221 ( .IN1(n3907), .IN2(n3906), .IN3(n3905), .Q(n3912) );
  AO21X1 U4222 ( .IN1(n4236), .IN2(n3913), .IN3(n4217), .Q(n3920) );
  NOR2X0 U4223 ( .IN1(InstAddrPointer[11]), .IN2(n4205), .QN(n3914) );
  NOR2X0 U4224 ( .IN1(n3920), .IN2(n3914), .QN(n3908) );
  OA22X1 U4225 ( .IN1(n4060), .IN2(n3909), .IN3(n3908), .IN4(n5228), .Q(n3911)
         );
  NAND3X0 U4226 ( .IN1(n3912), .IN2(n3911), .IN3(n3910), .QN(n2009) );
  INVX0 U4227 ( .INP(n3913), .ZN(n3915) );
  AO22X1 U4228 ( .IN1(n3916), .IN2(n4237), .IN3(n3915), .IN4(n3914), .Q(n3917)
         );
  AOI21X1 U4229 ( .IN1(n4290), .IN2(n3918), .IN3(n3917), .QN(n3925) );
  AOI22X1 U4230 ( .IN1(InstAddrPointer[11]), .IN2(n3920), .IN3(n3919), .IN4(
        n4288), .QN(n3924) );
  NAND2X0 U4231 ( .IN1(n3921), .IN2(n4287), .QN(n3922) );
  NAND4X0 U4232 ( .IN1(n3925), .IN2(n3924), .IN3(n3923), .IN4(n3922), .QN(
        n2010) );
  NAND2X0 U4233 ( .IN1(rEIP[9]), .IN2(n4281), .QN(n3927) );
  NAND2X0 U4234 ( .IN1(n4275), .IN2(EBX[9]), .QN(n3926) );
  AND3X1 U4235 ( .IN1(n4147), .IN2(n3927), .IN3(n3926), .Q(n3934) );
  XOR2X1 U4236 ( .IN1(n3929), .IN2(n3928), .Q(n3930) );
  NAND2X0 U4237 ( .IN1(n4280), .IN2(n3930), .QN(n3933) );
  NAND2X0 U4238 ( .IN1(n2090), .IN2(n3939), .QN(n3932) );
  NAND2X0 U4239 ( .IN1(PhyAddrPointer[9]), .IN2(n4274), .QN(n3931) );
  NAND4X0 U4240 ( .IN1(n3934), .IN2(n3933), .IN3(n3932), .IN4(n3931), .QN(
        n2056) );
  FADDX1 U4241 ( .A(n3993), .B(n3936), .CI(n3935), .CO(n3945), .S(n3982) );
  OA21X1 U4242 ( .IN1(n3989), .IN2(n3979), .IN3(n3944), .Q(n3984) );
  AOI22X1 U4243 ( .IN1(n3982), .IN2(n4266), .IN3(n3984), .IN4(n4262), .QN(
        n3942) );
  AND2X1 U4244 ( .IN1(n5098), .IN2(n3937), .Q(n3951) );
  INVX0 U4245 ( .INP(n3951), .ZN(n3938) );
  OA21X1 U4246 ( .IN1(n3937), .IN2(n5020), .IN3(n4221), .Q(n3949) );
  MUX21X1 U4247 ( .IN1(n3938), .IN2(n3949), .S(PhyAddrPointer[9]), .Q(n3941)
         );
  NAND2X0 U4248 ( .IN1(n4104), .IN2(rEIP[9]), .QN(n3986) );
  NAND2X0 U4249 ( .IN1(n4255), .IN2(n3939), .QN(n3940) );
  NAND4X0 U4250 ( .IN1(n3942), .IN2(n3941), .IN3(n3986), .IN4(n3940), .QN(
        n1727) );
  AO21X1 U4251 ( .IN1(n3965), .IN2(n3944), .IN3(n3943), .Q(n3964) );
  FADDX1 U4252 ( .A(n3947), .B(n3946), .CI(n3945), .CO(n3873), .S(n3948) );
  INVX0 U4253 ( .INP(n3948), .ZN(n3972) );
  OA22X1 U4254 ( .IN1(n4252), .IN2(n3964), .IN3(n3972), .IN4(n4248), .Q(n3955)
         );
  OA21X1 U4255 ( .IN1(PhyAddrPointer[9]), .IN2(n5020), .IN3(n3949), .Q(n3950)
         );
  NAND2X0 U4256 ( .IN1(n4104), .IN2(rEIP[10]), .QN(n3973) );
  OA21X1 U4257 ( .IN1(n3950), .IN2(n5195), .IN3(n3973), .Q(n3954) );
  NAND3X0 U4258 ( .IN1(PhyAddrPointer[9]), .IN2(n3951), .IN3(n5195), .QN(n3953) );
  NAND2X0 U4259 ( .IN1(n4255), .IN2(n3958), .QN(n3952) );
  NAND4X0 U4260 ( .IN1(n3955), .IN2(n3954), .IN3(n3953), .IN4(n3952), .QN(
        n1726) );
  XOR2X1 U4261 ( .IN1(n3957), .IN2(n3956), .Q(n3963) );
  OA22X1 U4262 ( .IN1(n4280), .IN2(n5258), .IN3(n5195), .IN4(n3288), .Q(n3961)
         );
  NAND2X0 U4263 ( .IN1(n2090), .IN2(n3958), .QN(n3960) );
  NAND2X0 U4264 ( .IN1(n4275), .IN2(EBX[10]), .QN(n3959) );
  NAND4X0 U4265 ( .IN1(n3961), .IN2(n4147), .IN3(n3960), .IN4(n3959), .QN(
        n3962) );
  AO21X1 U4266 ( .IN1(n4280), .IN2(n3963), .IN3(n3962), .Q(n2055) );
  OA22X1 U4267 ( .IN1(n3965), .IN2(n4206), .IN3(n4208), .IN4(n3964), .Q(n3970)
         );
  NAND3X0 U4268 ( .IN1(n4236), .IN2(n3966), .IN3(n5229), .QN(n3969) );
  NAND2X0 U4269 ( .IN1(n4290), .IN2(n3967), .QN(n3968) );
  AND3X1 U4270 ( .IN1(n3970), .IN2(n3969), .IN3(n3968), .Q(n3975) );
  AO21X1 U4271 ( .IN1(n4236), .IN2(n3976), .IN3(n4217), .Q(n3983) );
  NOR2X0 U4272 ( .IN1(InstAddrPointer[9]), .IN2(n4205), .QN(n3977) );
  NOR2X0 U4273 ( .IN1(n3983), .IN2(n3977), .QN(n3971) );
  OA22X1 U4274 ( .IN1(n4060), .IN2(n3972), .IN3(n3971), .IN4(n5229), .Q(n3974)
         );
  NAND3X0 U4275 ( .IN1(n3975), .IN2(n3974), .IN3(n3973), .QN(n2011) );
  INVX0 U4276 ( .INP(n3976), .ZN(n3978) );
  AO22X1 U4277 ( .IN1(n3979), .IN2(n4237), .IN3(n3978), .IN4(n3977), .Q(n3980)
         );
  AOI21X1 U4278 ( .IN1(n4290), .IN2(n3981), .IN3(n3980), .QN(n3988) );
  AOI22X1 U4279 ( .IN1(InstAddrPointer[9]), .IN2(n3983), .IN3(n3982), .IN4(
        n4288), .QN(n3987) );
  NAND2X0 U4280 ( .IN1(n3984), .IN2(n4287), .QN(n3985) );
  NAND4X0 U4281 ( .IN1(n3988), .IN2(n3987), .IN3(n3986), .IN4(n3985), .QN(
        n2012) );
  AO21X1 U4282 ( .IN1(n3990), .IN2(n4010), .IN3(n3989), .Q(n4009) );
  NAND2X0 U4283 ( .IN1(n4104), .IN2(rEIP[8]), .QN(n4020) );
  OA21X1 U4284 ( .IN1(n4252), .IN2(n4009), .IN3(n4020), .Q(n4000) );
  NOR2X0 U4285 ( .IN1(PhyAddrPointer[7]), .IN2(n5020), .QN(n4137) );
  OAI21X1 U4286 ( .IN1(n4136), .IN2(n4222), .IN3(n4221), .QN(n4135) );
  NOR2X0 U4287 ( .IN1(n4137), .IN2(n4135), .QN(n3995) );
  FADDX1 U4288 ( .A(n3993), .B(n3992), .CI(n3991), .CO(n3935), .S(n4011) );
  INVX0 U4289 ( .INP(n4011), .ZN(n3994) );
  OA22X1 U4290 ( .IN1(n3995), .IN2(n5189), .IN3(n4248), .IN4(n3994), .Q(n3999)
         );
  OR3X1 U4291 ( .IN1(PhyAddrPointer[8]), .IN2(n3996), .IN3(n5020), .Q(n3998)
         );
  NAND2X0 U4292 ( .IN1(n4255), .IN2(n4003), .QN(n3997) );
  NAND4X0 U4293 ( .IN1(n4000), .IN2(n3999), .IN3(n3998), .IN4(n3997), .QN(
        n1728) );
  XOR2X1 U4294 ( .IN1(n4002), .IN2(n4001), .Q(n4008) );
  OA22X1 U4295 ( .IN1(n4280), .IN2(n5259), .IN3(n5189), .IN4(n3288), .Q(n4006)
         );
  NAND2X0 U4296 ( .IN1(n2090), .IN2(n4003), .QN(n4005) );
  NAND2X0 U4297 ( .IN1(n4275), .IN2(EBX[8]), .QN(n4004) );
  NAND4X0 U4298 ( .IN1(n4006), .IN2(n4147), .IN3(n4005), .IN4(n4004), .QN(
        n4007) );
  AO21X1 U4299 ( .IN1(n4280), .IN2(n4008), .IN3(n4007), .Q(n2057) );
  OA22X1 U4300 ( .IN1(n4010), .IN2(n4206), .IN3(n4208), .IN4(n4009), .Q(n4015)
         );
  NAND2X0 U4301 ( .IN1(n4011), .IN2(n4288), .QN(n4014) );
  NAND2X0 U4302 ( .IN1(n4290), .IN2(n4012), .QN(n4013) );
  AND3X1 U4303 ( .IN1(n4015), .IN2(n4014), .IN3(n4013), .Q(n4021) );
  NAND2X0 U4304 ( .IN1(n5209), .IN2(n4236), .QN(n4153) );
  AO21X1 U4305 ( .IN1(n4236), .IN2(n4154), .IN3(n4217), .Q(n4151) );
  INVX0 U4306 ( .INP(n4151), .ZN(n4016) );
  AO21X1 U4307 ( .IN1(n4153), .IN2(n4016), .IN3(n5225), .Q(n4019) );
  NAND3X0 U4308 ( .IN1(n4236), .IN2(n4017), .IN3(n5225), .QN(n4018) );
  NAND4X0 U4309 ( .IN1(n4021), .IN2(n4020), .IN3(n4019), .IN4(n4018), .QN(
        n2013) );
  AOI22X1 U4310 ( .IN1(PhyAddrPointer[2]), .IN2(n4274), .IN3(n4275), .IN4(
        EBX[2]), .QN(n4028) );
  XOR2X1 U4311 ( .IN1(n4023), .IN2(n4022), .Q(n4024) );
  NAND2X0 U4312 ( .IN1(n4280), .IN2(n4024), .QN(n4027) );
  NAND2X0 U4313 ( .IN1(n2090), .IN2(n4036), .QN(n4026) );
  NAND2X0 U4314 ( .IN1(rEIP[2]), .IN2(n4281), .QN(n4025) );
  NAND4X0 U4315 ( .IN1(n4028), .IN2(n4027), .IN3(n4026), .IN4(n4025), .QN(
        n2063) );
  FADDX1 U4316 ( .A(n4030), .B(n4029), .CI(n4204), .CO(n4045), .S(n4209) );
  FADDX1 U4317 ( .A(n4033), .B(n4032), .CI(n4031), .CO(n4039), .S(n4210) );
  INVX0 U4318 ( .INP(n4221), .ZN(n4034) );
  AOI22X1 U4319 ( .IN1(n4266), .IN2(n4210), .IN3(PhyAddrPointer[2]), .IN4(
        n4034), .QN(n4035) );
  OA21X1 U4320 ( .IN1(n4252), .IN2(n4209), .IN3(n4035), .Q(n4038) );
  OR2X1 U4321 ( .IN1(PhyAddrPointer[2]), .IN2(n5020), .Q(n4042) );
  NAND2X0 U4322 ( .IN1(n4104), .IN2(rEIP[2]), .QN(n4207) );
  NAND2X0 U4323 ( .IN1(n4255), .IN2(n4036), .QN(n4037) );
  NAND4X0 U4324 ( .IN1(n4038), .IN2(n4042), .IN3(n4207), .IN4(n4037), .QN(
        n1734) );
  NOR2X0 U4325 ( .IN1(n4147), .IN2(n5217), .QN(n4063) );
  FADDX1 U4326 ( .A(n4041), .B(n4040), .CI(n4039), .CO(n4080), .S(n4058) );
  NAND2X0 U4327 ( .IN1(n4221), .IN2(n4042), .QN(n4083) );
  AO22X1 U4328 ( .IN1(n4266), .IN2(n4058), .IN3(PhyAddrPointer[3]), .IN4(n4083), .Q(n4043) );
  NOR2X0 U4329 ( .IN1(n4063), .IN2(n4043), .QN(n4049) );
  XNOR3X1 U4330 ( .IN1(n4070), .IN2(n4045), .IN3(n4044), .Q(n4062) );
  OR2X1 U4331 ( .IN1(n4252), .IN2(n4062), .Q(n4048) );
  NAND3X0 U4332 ( .IN1(n5098), .IN2(PhyAddrPointer[2]), .IN3(n5253), .QN(n4047) );
  NAND2X0 U4333 ( .IN1(n4255), .IN2(n4053), .QN(n4046) );
  NAND4X0 U4334 ( .IN1(n4049), .IN2(n4048), .IN3(n4047), .IN4(n4046), .QN(
        n1733) );
  AOI22X1 U4335 ( .IN1(PhyAddrPointer[3]), .IN2(n4274), .IN3(n4275), .IN4(
        EBX[3]), .QN(n4057) );
  XOR2X1 U4336 ( .IN1(n4051), .IN2(n4050), .Q(n4052) );
  NAND2X0 U4337 ( .IN1(n4280), .IN2(n4052), .QN(n4056) );
  NAND2X0 U4338 ( .IN1(n4053), .IN2(n2090), .QN(n4055) );
  NAND2X0 U4339 ( .IN1(rEIP[3]), .IN2(n4281), .QN(n4054) );
  NAND4X0 U4340 ( .IN1(n4057), .IN2(n4056), .IN3(n4055), .IN4(n4054), .QN(
        n2062) );
  INVX0 U4341 ( .INP(n4058), .ZN(n4059) );
  OA21X1 U4342 ( .IN1(n4189), .IN2(n4205), .IN3(n4294), .Q(n4194) );
  OA22X1 U4343 ( .IN1(n4060), .IN2(n4059), .IN3(n4194), .IN4(n5222), .Q(n4068)
         );
  NAND2X0 U4344 ( .IN1(n4236), .IN2(n5222), .QN(n4193) );
  OA22X1 U4345 ( .IN1(n4062), .IN2(n4208), .IN3(n4061), .IN4(n4193), .Q(n4067)
         );
  INVX0 U4346 ( .INP(n4063), .ZN(n4066) );
  NAND2X0 U4347 ( .IN1(n4290), .IN2(n4064), .QN(n4065) );
  NAND4X0 U4348 ( .IN1(n4068), .IN2(n4067), .IN3(n4066), .IN4(n4065), .QN(
        n4069) );
  AO21X1 U4349 ( .IN1(n4070), .IN2(n4237), .IN3(n4069), .Q(n2018) );
  XOR2X1 U4350 ( .IN1(n4072), .IN2(n4071), .Q(n4077) );
  AOI22X1 U4351 ( .IN1(PhyAddrPointer[4]), .IN2(n4274), .IN3(rEIP[4]), .IN4(
        n4281), .QN(n4075) );
  NAND2X0 U4352 ( .IN1(n4086), .IN2(n2090), .QN(n4074) );
  NAND2X0 U4353 ( .IN1(n4275), .IN2(EBX[4]), .QN(n4073) );
  NAND4X0 U4354 ( .IN1(n4075), .IN2(n4147), .IN3(n4074), .IN4(n4073), .QN(
        n4076) );
  AO21X1 U4355 ( .IN1(n4280), .IN2(n4077), .IN3(n4076), .Q(n2061) );
  XNOR3X1 U4356 ( .IN1(n4079), .IN2(n4198), .IN3(n4078), .Q(n4199) );
  FADDX1 U4357 ( .A(n4082), .B(n4081), .CI(n4080), .CO(n4100), .S(n4195) );
  AOI22X1 U4358 ( .IN1(n4266), .IN2(n4195), .IN3(PhyAddrPointer[4]), .IN4(
        n4083), .QN(n4089) );
  NOR2X0 U4359 ( .IN1(PhyAddrPointer[4]), .IN2(n5214), .QN(n4084) );
  MUX21X1 U4360 ( .IN1(PhyAddrPointer[4]), .IN2(n4084), .S(PhyAddrPointer[3]), 
        .Q(n4085) );
  NAND2X0 U4361 ( .IN1(n5098), .IN2(n4085), .QN(n4088) );
  NAND2X0 U4362 ( .IN1(n4255), .IN2(n4086), .QN(n4087) );
  NAND2X0 U4363 ( .IN1(n4104), .IN2(rEIP[4]), .QN(n4201) );
  NAND4X0 U4364 ( .IN1(n4089), .IN2(n4088), .IN3(n4087), .IN4(n4201), .QN(
        n4090) );
  AO21X1 U4365 ( .IN1(n4199), .IN2(n4262), .IN3(n4090), .Q(n1732) );
  XOR2X1 U4366 ( .IN1(n4092), .IN2(n4091), .Q(n4097) );
  OA22X1 U4367 ( .IN1(n4280), .IN2(n5260), .IN3(n5181), .IN4(n3288), .Q(n4095)
         );
  NAND2X0 U4368 ( .IN1(n4103), .IN2(n2090), .QN(n4094) );
  NAND2X0 U4369 ( .IN1(n4275), .IN2(EBX[5]), .QN(n4093) );
  NAND4X0 U4370 ( .IN1(n4095), .IN2(n4147), .IN3(n4094), .IN4(n4093), .QN(
        n4096) );
  AO21X1 U4371 ( .IN1(n4280), .IN2(n4097), .IN3(n4096), .Q(n2060) );
  XNOR3X1 U4372 ( .IN1(n4166), .IN2(n4099), .IN3(n4098), .Q(n4173) );
  FADDX1 U4373 ( .A(n4102), .B(n4101), .CI(n4100), .CO(n4118), .S(n4163) );
  OAI21X1 U4374 ( .IN1(n4122), .IN2(n4222), .IN3(n4221), .QN(n4121) );
  AOI22X1 U4375 ( .IN1(n4266), .IN2(n4163), .IN3(PhyAddrPointer[5]), .IN4(
        n4121), .QN(n4107) );
  NAND3X0 U4376 ( .IN1(n4122), .IN2(n5098), .IN3(n5181), .QN(n4106) );
  NAND2X0 U4377 ( .IN1(n4255), .IN2(n4103), .QN(n4105) );
  NAND2X0 U4378 ( .IN1(n4104), .IN2(rEIP[5]), .QN(n4169) );
  NAND4X0 U4379 ( .IN1(n4107), .IN2(n4106), .IN3(n4105), .IN4(n4169), .QN(
        n4108) );
  AO21X1 U4380 ( .IN1(n4173), .IN2(n4262), .IN3(n4108), .Q(n1731) );
  XOR2X1 U4381 ( .IN1(n4110), .IN2(n4109), .Q(n4115) );
  OA22X1 U4382 ( .IN1(n4280), .IN2(n5261), .IN3(n5184), .IN4(n3288), .Q(n4113)
         );
  NAND2X0 U4383 ( .IN1(n4126), .IN2(n2090), .QN(n4112) );
  NAND2X0 U4384 ( .IN1(n4275), .IN2(EBX[6]), .QN(n4111) );
  NAND4X0 U4385 ( .IN1(n4113), .IN2(n4147), .IN3(n4112), .IN4(n4111), .QN(
        n4114) );
  AO21X1 U4386 ( .IN1(n4280), .IN2(n4115), .IN3(n4114), .Q(n2059) );
  XNOR3X1 U4387 ( .IN1(n4179), .IN2(n4117), .IN3(n4116), .Q(n4188) );
  FADDX1 U4388 ( .A(n4120), .B(n4119), .CI(n4118), .CO(n4133), .S(n4182) );
  AOI22X1 U4389 ( .IN1(PhyAddrPointer[6]), .IN2(n4121), .IN3(n4266), .IN4(
        n4182), .QN(n4129) );
  INVX0 U4390 ( .INP(n4122), .ZN(n4123) );
  OA21X1 U4391 ( .IN1(PhyAddrPointer[6]), .IN2(n4123), .IN3(PhyAddrPointer[5]), 
        .Q(n4125) );
  NOR2X0 U4392 ( .IN1(PhyAddrPointer[6]), .IN2(PhyAddrPointer[5]), .QN(n4124)
         );
  OR3X1 U4393 ( .IN1(n4125), .IN2(n4124), .IN3(n5020), .Q(n4128) );
  NAND2X0 U4394 ( .IN1(n4255), .IN2(n4126), .QN(n4127) );
  NAND2X0 U4395 ( .IN1(n4104), .IN2(rEIP[6]), .QN(n4185) );
  NAND4X0 U4396 ( .IN1(n4129), .IN2(n4128), .IN3(n4127), .IN4(n4185), .QN(
        n4130) );
  AO21X1 U4397 ( .IN1(n4188), .IN2(n4262), .IN3(n4130), .Q(n1730) );
  XNOR3X1 U4398 ( .IN1(n4132), .IN2(n4155), .IN3(n4131), .Q(n4162) );
  XOR2X1 U4399 ( .IN1(n4134), .IN2(n4133), .Q(n4152) );
  AOI22X1 U4400 ( .IN1(PhyAddrPointer[7]), .IN2(n4135), .IN3(n4266), .IN4(
        n4152), .QN(n4140) );
  NAND2X0 U4401 ( .IN1(n4137), .IN2(n4136), .QN(n4139) );
  NAND2X0 U4402 ( .IN1(n4255), .IN2(n4144), .QN(n4138) );
  NAND2X0 U4403 ( .IN1(rEIP[7]), .IN2(n4104), .QN(n4158) );
  NAND4X0 U4404 ( .IN1(n4140), .IN2(n4139), .IN3(n4138), .IN4(n4158), .QN(
        n4141) );
  AO21X1 U4405 ( .IN1(n4162), .IN2(n4262), .IN3(n4141), .Q(n1729) );
  XOR2X1 U4406 ( .IN1(n4143), .IN2(n4142), .Q(n4150) );
  AOI22X1 U4407 ( .IN1(rEIP[7]), .IN2(n4281), .IN3(PhyAddrPointer[7]), .IN4(
        n4274), .QN(n4148) );
  NAND2X0 U4408 ( .IN1(n4144), .IN2(n2090), .QN(n4146) );
  NAND2X0 U4409 ( .IN1(n4275), .IN2(EBX[7]), .QN(n4145) );
  NAND4X0 U4410 ( .IN1(n4148), .IN2(n4147), .IN3(n4146), .IN4(n4145), .QN(
        n4149) );
  AO21X1 U4411 ( .IN1(n4280), .IN2(n4150), .IN3(n4149), .Q(n2058) );
  AOI22X1 U4412 ( .IN1(n4152), .IN2(n4288), .IN3(InstAddrPointer[7]), .IN4(
        n4151), .QN(n4160) );
  OA22X1 U4413 ( .IN1(n4206), .IN2(n4155), .IN3(n4154), .IN4(n4153), .Q(n4159)
         );
  NAND2X0 U4414 ( .IN1(n4290), .IN2(n4156), .QN(n4157) );
  NAND4X0 U4415 ( .IN1(n4160), .IN2(n4159), .IN3(n4158), .IN4(n4157), .QN(
        n4161) );
  AO21X1 U4416 ( .IN1(n4162), .IN2(n4287), .IN3(n4161), .Q(n2014) );
  AO21X1 U4417 ( .IN1(n4236), .IN2(n4180), .IN3(n4217), .Q(n4164) );
  AOI22X1 U4418 ( .IN1(n4164), .IN2(InstAddrPointer[5]), .IN3(n4163), .IN4(
        n4288), .QN(n4171) );
  NAND2X0 U4419 ( .IN1(n4236), .IN2(n5205), .QN(n4165) );
  OA22X1 U4420 ( .IN1(n4206), .IN2(n4166), .IN3(n4180), .IN4(n4165), .Q(n4170)
         );
  NAND2X0 U4421 ( .IN1(n4290), .IN2(n4167), .QN(n4168) );
  NAND4X0 U4422 ( .IN1(n4171), .IN2(n4170), .IN3(n4169), .IN4(n4168), .QN(
        n4172) );
  AO21X1 U4423 ( .IN1(n4173), .IN2(n4287), .IN3(n4172), .Q(n2016) );
  NAND2X0 U4424 ( .IN1(n4236), .IN2(n4174), .QN(n4177) );
  NAND2X0 U4425 ( .IN1(n4290), .IN2(n4175), .QN(n4176) );
  OA21X1 U4426 ( .IN1(InstAddrPointer[6]), .IN2(n4177), .IN3(n4176), .Q(n4178)
         );
  OA21X1 U4427 ( .IN1(n4179), .IN2(n4206), .IN3(n4178), .Q(n4186) );
  OA21X1 U4428 ( .IN1(n4180), .IN2(n5205), .IN3(n4236), .Q(n4181) );
  OAI21X1 U4429 ( .IN1(n4217), .IN2(n4181), .IN3(InstAddrPointer[6]), .QN(
        n4184) );
  NAND2X0 U4430 ( .IN1(n4182), .IN2(n4288), .QN(n4183) );
  NAND4X0 U4431 ( .IN1(n4186), .IN2(n4185), .IN3(n4184), .IN4(n4183), .QN(
        n4187) );
  AO21X1 U4432 ( .IN1(n4188), .IN2(n4287), .IN3(n4187), .Q(n2015) );
  NAND3X0 U4433 ( .IN1(InstAddrPointer[3]), .IN2(n4236), .IN3(n4189), .QN(
        n4192) );
  NAND2X0 U4434 ( .IN1(n4290), .IN2(n4190), .QN(n4191) );
  OA21X1 U4435 ( .IN1(n4192), .IN2(InstAddrPointer[4]), .IN3(n4191), .Q(n4203)
         );
  NAND2X0 U4436 ( .IN1(n4194), .IN2(n4193), .QN(n4196) );
  AOI22X1 U4437 ( .IN1(n4196), .IN2(InstAddrPointer[4]), .IN3(n4195), .IN4(
        n4288), .QN(n4197) );
  OA21X1 U4438 ( .IN1(n4198), .IN2(n4206), .IN3(n4197), .Q(n4202) );
  NAND2X0 U4439 ( .IN1(n4199), .IN2(n4287), .QN(n4200) );
  NAND4X0 U4440 ( .IN1(n4203), .IN2(n4202), .IN3(n4201), .IN4(n4200), .QN(
        n2017) );
  MUX21X1 U4441 ( .IN1(n4206), .IN2(n4205), .S(n4204), .Q(n4215) );
  OA21X1 U4442 ( .IN1(n4209), .IN2(n4208), .IN3(n4207), .Q(n4214) );
  NAND2X0 U4443 ( .IN1(n4210), .IN2(n4288), .QN(n4213) );
  NAND2X0 U4444 ( .IN1(n4290), .IN2(n4211), .QN(n4212) );
  NAND4X0 U4445 ( .IN1(n4215), .IN2(n4214), .IN3(n4213), .IN4(n4212), .QN(
        n4216) );
  AO21X1 U4446 ( .IN1(n4217), .IN2(InstAddrPointer[2]), .IN3(n4216), .Q(n2019)
         );
  FADDX1 U4447 ( .A(n4220), .B(n4219), .CI(n4218), .CO(n4031), .S(n4235) );
  NAND2X0 U4448 ( .IN1(n4222), .IN2(n4221), .QN(n4263) );
  AOI22X1 U4449 ( .IN1(n4266), .IN2(n4235), .IN3(n4263), .IN4(
        PhyAddrPointer[1]), .QN(n4226) );
  XOR3X1 U4450 ( .IN1(n4238), .IN2(n4260), .IN3(n4223), .Q(n4240) );
  NAND2X0 U4451 ( .IN1(n4262), .IN2(n4240), .QN(n4225) );
  NAND2X0 U4452 ( .IN1(n4255), .IN2(n5201), .QN(n4224) );
  NAND2X0 U4453 ( .IN1(n4104), .IN2(N4154), .QN(n4242) );
  NAND4X0 U4454 ( .IN1(n4226), .IN2(n4225), .IN3(n4224), .IN4(n4242), .QN(
        n1735) );
  AOI22X1 U4455 ( .IN1(PhyAddrPointer[1]), .IN2(n4274), .IN3(n4275), .IN4(
        EBX[1]), .QN(n4234) );
  FADDX1 U4456 ( .A(n4229), .B(n4228), .CI(n4227), .CO(n4022), .S(n4230) );
  NAND2X0 U4457 ( .IN1(n4280), .IN2(n4230), .QN(n4233) );
  NAND2X0 U4458 ( .IN1(n5201), .IN2(n2090), .QN(n4232) );
  NAND2X0 U4459 ( .IN1(N4154), .IN2(n4281), .QN(n4231) );
  NAND4X0 U4460 ( .IN1(n4234), .IN2(n4233), .IN3(n4232), .IN4(n4231), .QN(
        n2064) );
  AOI22X1 U4461 ( .IN1(n5185), .IN2(n4290), .IN3(n4235), .IN4(n4288), .QN(
        n4244) );
  NOR2X0 U4462 ( .IN1(n4237), .IN2(n4236), .QN(n4295) );
  OR2X1 U4463 ( .IN1(n4295), .IN2(n4238), .Q(n4239) );
  OA21X1 U4464 ( .IN1(n4294), .IN2(n5185), .IN3(n4239), .Q(n4243) );
  NAND2X0 U4465 ( .IN1(n4287), .IN2(n4240), .QN(n4241) );
  NAND4X0 U4466 ( .IN1(n4244), .IN2(n4243), .IN3(n4242), .IN4(n4241), .QN(
        n2020) );
  OA21X1 U4467 ( .IN1(PhyAddrPointer[30]), .IN2(n5020), .IN3(n4245), .Q(n4249)
         );
  INVX0 U4468 ( .INP(n4246), .ZN(n4247) );
  OA22X1 U4469 ( .IN1(n4249), .IN2(n5239), .IN3(n4248), .IN4(n4247), .Q(n4259)
         );
  OA21X1 U4470 ( .IN1(n4252), .IN2(n4251), .IN3(n4250), .Q(n4258) );
  NAND3X0 U4471 ( .IN1(PhyAddrPointer[30]), .IN2(n4253), .IN3(n5239), .QN(
        n4257) );
  NAND2X0 U4472 ( .IN1(n4255), .IN2(n4254), .QN(n4256) );
  NAND4X0 U4473 ( .IN1(n4259), .IN2(n4258), .IN3(n4257), .IN4(n4256), .QN(
        n1705) );
  OA21X1 U4474 ( .IN1(n4261), .IN2(n5204), .IN3(n4260), .Q(n4286) );
  NAND2X0 U4475 ( .IN1(n4262), .IN2(n4286), .QN(n4270) );
  NAND2X0 U4476 ( .IN1(n4104), .IN2(rEIP[0]), .QN(n4296) );
  OA21X1 U4477 ( .IN1(n5196), .IN2(n4431), .IN3(n4296), .Q(n4269) );
  NAND2X0 U4478 ( .IN1(n4263), .IN2(N1009), .QN(n4268) );
  HADDX1 U4479 ( .A0(n4265), .B0(n4264), .C1(n4219), .SO(n4289) );
  NAND2X0 U4480 ( .IN1(n4266), .IN2(n4289), .QN(n4267) );
  NAND4X0 U4481 ( .IN1(n4270), .IN2(n4269), .IN3(n4268), .IN4(n4267), .QN(
        n1736) );
  AO22X1 U4482 ( .IN1(n4445), .IN2(n4272), .IN3(n4271), .IN4(n5016), .Q(n4273)
         );
  MUX21X1 U4483 ( .IN1(n4273), .IN2(InstQueueRd_Addr[3]), .S(n4302), .Q(n2025)
         );
  AOI22X1 U4484 ( .IN1(n4275), .IN2(EBX[0]), .IN3(n4274), .IN4(N1009), .QN(
        n4285) );
  FADDX1 U4485 ( .A(n4278), .B(n4277), .CI(n4276), .CO(n4227), .S(n4279) );
  NAND2X0 U4486 ( .IN1(n4280), .IN2(n4279), .QN(n4284) );
  NAND2X0 U4487 ( .IN1(n2090), .IN2(N1009), .QN(n4283) );
  NAND2X0 U4488 ( .IN1(rEIP[0]), .IN2(n4281), .QN(n4282) );
  NAND4X0 U4489 ( .IN1(n4285), .IN2(n4284), .IN3(n4283), .IN4(n4282), .QN(
        n2065) );
  NAND2X0 U4490 ( .IN1(n4287), .IN2(n4286), .QN(n4293) );
  NAND2X0 U4491 ( .IN1(n4289), .IN2(n4288), .QN(n4292) );
  NAND2X0 U4492 ( .IN1(n4290), .IN2(N1868), .QN(n4291) );
  AND3X1 U4493 ( .IN1(n4293), .IN2(n4292), .IN3(n4291), .Q(n4298) );
  MUX21X1 U4494 ( .IN1(n4295), .IN2(n4294), .S(N1868), .Q(n4297) );
  NAND3X0 U4495 ( .IN1(n4298), .IN2(n4297), .IN3(n4296), .QN(n2021) );
  AO22X1 U4496 ( .IN1(n4299), .IN2(n4445), .IN3(n5016), .IN4(n5183), .Q(n4300)
         );
  AO21X1 U4497 ( .IN1(n4495), .IN2(n5204), .IN3(n4300), .Q(n4301) );
  MUX21X1 U4498 ( .IN1(n4301), .IN2(N2884), .S(n4302), .Q(n2028) );
  AO21X1 U4499 ( .IN1(n5016), .IN2(n4303), .IN3(n4302), .Q(n4312) );
  NAND2X0 U4500 ( .IN1(n4445), .IN2(n4304), .QN(n4309) );
  NAND3X0 U4501 ( .IN1(N1868), .IN2(n4495), .IN3(n4305), .QN(n4308) );
  NAND3X0 U4502 ( .IN1(n4306), .IN2(n5016), .IN3(n5180), .QN(n4307) );
  NAND3X0 U4503 ( .IN1(n4309), .IN2(n4308), .IN3(n4307), .QN(n4311) );
  AO22X1 U4504 ( .IN1(InstQueueRd_Addr[2]), .IN2(n4312), .IN3(n4311), .IN4(
        n4310), .Q(n2026) );
  NAND2X0 U4505 ( .IN1(READY_n), .IN2(State[1]), .QN(n4460) );
  OA22X1 U4506 ( .IN1(State[1]), .IN2(RequestPending), .IN3(NA_n), .IN4(n4460), 
        .Q(n4313) );
  NAND2X0 U4507 ( .IN1(n4313), .IN2(n5207), .QN(n4314) );
  NAND3X0 U4508 ( .IN1(n4314), .IN2(HOLD), .IN3(State[0]), .QN(n4317) );
  OR2X1 U4509 ( .IN1(n5207), .IN2(n4460), .Q(n4316) );
  NAND2X0 U4510 ( .IN1(State[2]), .IN2(n5202), .QN(n4462) );
  NAND2X0 U4511 ( .IN1(State[0]), .IN2(RequestPending), .QN(n4459) );
  AO221X1 U4512 ( .IN1(n4462), .IN2(n4460), .IN3(n4462), .IN4(n4459), .IN5(
        NA_n), .Q(n4315) );
  NOR2X1 U4513 ( .IN1(State[0]), .IN2(n5178), .QN(n5168) );
  NAND2X0 U4514 ( .IN1(n5168), .IN2(State[2]), .QN(n4334) );
  NAND4X0 U4515 ( .IN1(n4317), .IN2(n4316), .IN3(n4315), .IN4(n4334), .QN(
        n2074) );
  AO222X1 U4516 ( .IN1(Datai[15]), .IN2(n4320), .IN3(\C1/DATA2_15 ), .IN4(
        n4319), .IN5(EAX[15]), .IN6(n4318), .Q(n1928) );
  NAND2X0 U4517 ( .IN1(EAX[31]), .IN2(n4321), .QN(n4331) );
  NAND2X0 U4518 ( .IN1(n4322), .IN2(Datai[31]), .QN(n4330) );
  HADDX1 U4519 ( .A0(n4324), .B0(n4323), .C1(n4325), .SO(n2601) );
  XOR2X1 U4520 ( .IN1(n4325), .IN2(EAX[31]), .Q(n4326) );
  NAND3X0 U4521 ( .IN1(n4328), .IN2(n4327), .IN3(n4326), .QN(n4329) );
  NAND3X0 U4522 ( .IN1(n4331), .IN2(n4330), .IN3(n4329), .QN(n1959) );
  OR2X1 U4523 ( .IN1(n5190), .IN2(n5248), .Q(n4333) );
  NAND2X0 U4524 ( .IN1(rEIP[31]), .IN2(rEIP[0]), .QN(n4332) );
  OAI21X1 U4525 ( .IN1(n4333), .IN2(State[2]), .IN3(n4332), .QN(n4337) );
  INVX0 U4526 ( .INP(n4334), .ZN(n4422) );
  AO22X1 U4527 ( .IN1(N4154), .IN2(n4422), .IN3(rEIP[2]), .IN4(n5207), .Q(
        n4336) );
  MUX21X1 U4528 ( .IN1(Address[0]), .IN2(n4335), .S(n5168), .Q(n1702) );
  HADDX1 U4529 ( .A0(n4337), .B0(n4336), .C1(n4340), .SO(n4335) );
  AO22X1 U4530 ( .IN1(rEIP[3]), .IN2(n5207), .IN3(rEIP[2]), .IN4(n4422), .Q(
        n4339) );
  MUX21X1 U4531 ( .IN1(Address[1]), .IN2(n4338), .S(n5168), .Q(n1701) );
  HADDX1 U4532 ( .A0(n4340), .B0(n4339), .C1(n4343), .SO(n4338) );
  AO22X1 U4533 ( .IN1(rEIP[4]), .IN2(n5207), .IN3(rEIP[3]), .IN4(n4422), .Q(
        n4342) );
  MUX21X1 U4534 ( .IN1(Address[2]), .IN2(n4341), .S(n5168), .Q(n1700) );
  HADDX1 U4535 ( .A0(n4343), .B0(n4342), .C1(n4346), .SO(n4341) );
  AO22X1 U4536 ( .IN1(rEIP[4]), .IN2(n4422), .IN3(rEIP[5]), .IN4(n5207), .Q(
        n4345) );
  MUX21X1 U4537 ( .IN1(Address[3]), .IN2(n4344), .S(n5168), .Q(n1699) );
  HADDX1 U4538 ( .A0(n4346), .B0(n4345), .C1(n4349), .SO(n4344) );
  AO22X1 U4539 ( .IN1(rEIP[6]), .IN2(n5207), .IN3(rEIP[5]), .IN4(n4422), .Q(
        n4348) );
  MUX21X1 U4540 ( .IN1(Address[4]), .IN2(n4347), .S(n5168), .Q(n1698) );
  HADDX1 U4541 ( .A0(n4349), .B0(n4348), .C1(n4352), .SO(n4347) );
  AO22X1 U4542 ( .IN1(rEIP[7]), .IN2(n5207), .IN3(rEIP[6]), .IN4(n4422), .Q(
        n4351) );
  MUX21X1 U4543 ( .IN1(Address[5]), .IN2(n4350), .S(n5168), .Q(n1697) );
  HADDX1 U4544 ( .A0(n4352), .B0(n4351), .C1(n4355), .SO(n4350) );
  AO22X1 U4545 ( .IN1(rEIP[7]), .IN2(n4422), .IN3(rEIP[8]), .IN4(n5207), .Q(
        n4354) );
  MUX21X1 U4546 ( .IN1(Address[6]), .IN2(n4353), .S(n5168), .Q(n1696) );
  HADDX1 U4547 ( .A0(n4355), .B0(n4354), .C1(n4358), .SO(n4353) );
  AO22X1 U4548 ( .IN1(rEIP[9]), .IN2(n5207), .IN3(rEIP[8]), .IN4(n4422), .Q(
        n4357) );
  MUX21X1 U4549 ( .IN1(Address[7]), .IN2(n4356), .S(n5168), .Q(n1695) );
  HADDX1 U4550 ( .A0(n4358), .B0(n4357), .C1(n4361), .SO(n4356) );
  AO22X1 U4551 ( .IN1(rEIP[9]), .IN2(n4422), .IN3(rEIP[10]), .IN4(n5207), .Q(
        n4360) );
  MUX21X1 U4552 ( .IN1(Address[8]), .IN2(n4359), .S(n5168), .Q(n1694) );
  HADDX1 U4553 ( .A0(n4361), .B0(n4360), .C1(n4364), .SO(n4359) );
  AO22X1 U4554 ( .IN1(rEIP[11]), .IN2(n5207), .IN3(rEIP[10]), .IN4(n4422), .Q(
        n4363) );
  MUX21X1 U4555 ( .IN1(Address[9]), .IN2(n4362), .S(n5168), .Q(n1693) );
  HADDX1 U4556 ( .A0(n4364), .B0(n4363), .C1(n4367), .SO(n4362) );
  AO22X1 U4557 ( .IN1(rEIP[11]), .IN2(n4422), .IN3(rEIP[12]), .IN4(n5207), .Q(
        n4366) );
  MUX21X1 U4558 ( .IN1(Address[10]), .IN2(n4365), .S(n5168), .Q(n1692) );
  HADDX1 U4559 ( .A0(n4367), .B0(n4366), .C1(n4370), .SO(n4365) );
  AO22X1 U4560 ( .IN1(rEIP[13]), .IN2(n5207), .IN3(rEIP[12]), .IN4(n4422), .Q(
        n4369) );
  MUX21X1 U4561 ( .IN1(Address[11]), .IN2(n4368), .S(n5168), .Q(n1691) );
  HADDX1 U4562 ( .A0(n4370), .B0(n4369), .C1(n4373), .SO(n4368) );
  AO22X1 U4563 ( .IN1(rEIP[13]), .IN2(n4422), .IN3(rEIP[14]), .IN4(n5207), .Q(
        n4372) );
  MUX21X1 U4564 ( .IN1(Address[12]), .IN2(n4371), .S(n5168), .Q(n1690) );
  HADDX1 U4565 ( .A0(n4373), .B0(n4372), .C1(n4376), .SO(n4371) );
  AO22X1 U4566 ( .IN1(rEIP[15]), .IN2(n5207), .IN3(rEIP[14]), .IN4(n4422), .Q(
        n4375) );
  MUX21X1 U4567 ( .IN1(Address[13]), .IN2(n4374), .S(n5168), .Q(n1689) );
  HADDX1 U4568 ( .A0(n4376), .B0(n4375), .C1(n4379), .SO(n4374) );
  AO22X1 U4569 ( .IN1(rEIP[15]), .IN2(n4422), .IN3(rEIP[16]), .IN4(n5207), .Q(
        n4378) );
  MUX21X1 U4570 ( .IN1(Address[14]), .IN2(n4377), .S(n5168), .Q(n1688) );
  HADDX1 U4571 ( .A0(n4379), .B0(n4378), .C1(n4382), .SO(n4377) );
  AO22X1 U4572 ( .IN1(rEIP[17]), .IN2(n5207), .IN3(rEIP[16]), .IN4(n4422), .Q(
        n4381) );
  MUX21X1 U4573 ( .IN1(Address[15]), .IN2(n4380), .S(n5168), .Q(n1687) );
  HADDX1 U4574 ( .A0(n4382), .B0(n4381), .C1(n4385), .SO(n4380) );
  AO22X1 U4575 ( .IN1(rEIP[17]), .IN2(n4422), .IN3(rEIP[18]), .IN4(n5207), .Q(
        n4384) );
  MUX21X1 U4576 ( .IN1(Address[16]), .IN2(n4383), .S(n5168), .Q(n1686) );
  HADDX1 U4577 ( .A0(n4385), .B0(n4384), .C1(n4388), .SO(n4383) );
  AO22X1 U4578 ( .IN1(rEIP[19]), .IN2(n5207), .IN3(rEIP[18]), .IN4(n4422), .Q(
        n4387) );
  MUX21X1 U4579 ( .IN1(Address[17]), .IN2(n4386), .S(n5168), .Q(n1685) );
  HADDX1 U4580 ( .A0(n4388), .B0(n4387), .C1(n4391), .SO(n4386) );
  AO22X1 U4581 ( .IN1(rEIP[19]), .IN2(n4422), .IN3(rEIP[20]), .IN4(n5207), .Q(
        n4390) );
  MUX21X1 U4582 ( .IN1(Address[18]), .IN2(n4389), .S(n5168), .Q(n1684) );
  HADDX1 U4583 ( .A0(n4391), .B0(n4390), .C1(n4394), .SO(n4389) );
  AO22X1 U4584 ( .IN1(rEIP[21]), .IN2(n5207), .IN3(rEIP[20]), .IN4(n4422), .Q(
        n4393) );
  MUX21X1 U4585 ( .IN1(Address[19]), .IN2(n4392), .S(n5168), .Q(n1683) );
  HADDX1 U4586 ( .A0(n4394), .B0(n4393), .C1(n4397), .SO(n4392) );
  AO22X1 U4587 ( .IN1(rEIP[21]), .IN2(n4422), .IN3(rEIP[22]), .IN4(n5207), .Q(
        n4396) );
  MUX21X1 U4588 ( .IN1(Address[20]), .IN2(n4395), .S(n5168), .Q(n1682) );
  HADDX1 U4589 ( .A0(n4397), .B0(n4396), .C1(n4400), .SO(n4395) );
  AO22X1 U4590 ( .IN1(rEIP[23]), .IN2(n5207), .IN3(rEIP[22]), .IN4(n4422), .Q(
        n4399) );
  MUX21X1 U4591 ( .IN1(Address[21]), .IN2(n4398), .S(n5168), .Q(n1681) );
  HADDX1 U4592 ( .A0(n4400), .B0(n4399), .C1(n4403), .SO(n4398) );
  AO22X1 U4593 ( .IN1(rEIP[23]), .IN2(n4422), .IN3(rEIP[24]), .IN4(n5207), .Q(
        n4402) );
  MUX21X1 U4594 ( .IN1(Address[22]), .IN2(n4401), .S(n5168), .Q(n1680) );
  HADDX1 U4595 ( .A0(n4403), .B0(n4402), .C1(n4406), .SO(n4401) );
  AO22X1 U4596 ( .IN1(rEIP[25]), .IN2(n5207), .IN3(rEIP[24]), .IN4(n4422), .Q(
        n4405) );
  MUX21X1 U4597 ( .IN1(Address[23]), .IN2(n4404), .S(n5168), .Q(n1679) );
  HADDX1 U4598 ( .A0(n4406), .B0(n4405), .C1(n4409), .SO(n4404) );
  AO22X1 U4599 ( .IN1(rEIP[25]), .IN2(n4422), .IN3(rEIP[26]), .IN4(n5207), .Q(
        n4408) );
  MUX21X1 U4600 ( .IN1(Address[24]), .IN2(n4407), .S(n5168), .Q(n1678) );
  HADDX1 U4601 ( .A0(n4409), .B0(n4408), .C1(n4412), .SO(n4407) );
  AO22X1 U4602 ( .IN1(rEIP[27]), .IN2(n5207), .IN3(rEIP[26]), .IN4(n4422), .Q(
        n4411) );
  MUX21X1 U4603 ( .IN1(Address[25]), .IN2(n4410), .S(n5168), .Q(n1677) );
  HADDX1 U4604 ( .A0(n4412), .B0(n4411), .C1(n4415), .SO(n4410) );
  AO22X1 U4605 ( .IN1(rEIP[27]), .IN2(n4422), .IN3(rEIP[28]), .IN4(n5207), .Q(
        n4414) );
  MUX21X1 U4606 ( .IN1(Address[26]), .IN2(n4413), .S(n5168), .Q(n1676) );
  HADDX1 U4607 ( .A0(n4415), .B0(n4414), .C1(n4418), .SO(n4413) );
  AO22X1 U4608 ( .IN1(rEIP[29]), .IN2(n5207), .IN3(rEIP[28]), .IN4(n4422), .Q(
        n4417) );
  MUX21X1 U4609 ( .IN1(Address[27]), .IN2(n4416), .S(n5168), .Q(n1675) );
  HADDX1 U4610 ( .A0(n4418), .B0(n4417), .C1(n4421), .SO(n4416) );
  AO22X1 U4611 ( .IN1(rEIP[30]), .IN2(n5207), .IN3(rEIP[29]), .IN4(n4422), .Q(
        n4420) );
  MUX21X1 U4612 ( .IN1(Address[28]), .IN2(n4419), .S(n5168), .Q(n1674) );
  HADDX1 U4613 ( .A0(n4421), .B0(n4420), .C1(n4424), .SO(n4419) );
  AO22X1 U4614 ( .IN1(rEIP[31]), .IN2(n5207), .IN3(rEIP[30]), .IN4(n4422), .Q(
        n4423) );
  XOR2X1 U4615 ( .IN1(n4424), .IN2(n4423), .Q(n4425) );
  MUX21X1 U4616 ( .IN1(Address[29]), .IN2(n4425), .S(n5168), .Q(n1673) );
  INVX0 U4617 ( .INP(n5097), .ZN(n4428) );
  NOR2X0 U4618 ( .IN1(N4188), .IN2(n4426), .QN(n5102) );
  NOR2X0 U4619 ( .IN1(n5200), .IN2(N4187), .QN(n4849) );
  NAND2X0 U4620 ( .IN1(n4604), .IN2(n4849), .QN(n5019) );
  INVX0 U4621 ( .INP(n5019), .ZN(n4432) );
  NOR2X0 U4622 ( .IN1(n5102), .IN2(n4432), .QN(n4427) );
  AO222X1 U4623 ( .IN1(n5020), .IN2(n4428), .IN3(n5020), .IN4(n4485), .IN5(
        n4428), .IN6(n4427), .Q(n4429) );
  OA21X1 U4624 ( .IN1(n4431), .IN2(n4430), .IN3(n4429), .Q(n5089) );
  INVX0 U4625 ( .INP(n5089), .ZN(n5069) );
  NAND2X0 U4626 ( .IN1(n4432), .IN2(n5069), .QN(n5086) );
  OA22X1 U4627 ( .IN1(n5089), .IN2(n5156), .IN3(n5086), .IN4(n5155), .Q(n4437)
         );
  NAND2X0 U4628 ( .IN1(n5102), .IN2(n5199), .QN(n4971) );
  NAND3X0 U4629 ( .IN1(n5098), .IN2(n5019), .IN3(n5069), .QN(n4433) );
  NOR2X0 U4630 ( .IN1(n4971), .IN2(n4433), .QN(n5087) );
  NAND2X0 U4631 ( .IN1(n5158), .IN2(n5087), .QN(n4436) );
  INVX0 U4632 ( .INP(n4971), .ZN(n5099) );
  NOR2X0 U4633 ( .IN1(n5099), .IN2(n4433), .QN(n5088) );
  NAND2X0 U4634 ( .IN1(Datai[7]), .IN2(n5088), .QN(n4435) );
  NAND2X0 U4635 ( .IN1(\InstQueue[14][7] ), .IN2(n5089), .QN(n4434) );
  NAND4X0 U4636 ( .IN1(n4437), .IN2(n4436), .IN3(n4435), .IN4(n4434), .QN(
        n1745) );
  NOR4X0 U4637 ( .IN1(EAX[12]), .IN2(EAX[13]), .IN3(EAX[14]), .IN4(EAX[15]), 
        .QN(n4441) );
  NOR4X0 U4638 ( .IN1(EAX[8]), .IN2(EAX[9]), .IN3(EAX[10]), .IN4(EAX[11]), 
        .QN(n4440) );
  NOR4X0 U4639 ( .IN1(EAX[4]), .IN2(EAX[5]), .IN3(EAX[6]), .IN4(EAX[7]), .QN(
        n4439) );
  NOR4X0 U4640 ( .IN1(EAX[0]), .IN2(EAX[1]), .IN3(EAX[2]), .IN4(EAX[3]), .QN(
        n4438) );
  NAND4X0 U4641 ( .IN1(n4441), .IN2(n4440), .IN3(n4439), .IN4(n4438), .QN(
        n4442) );
  AND2X1 U4642 ( .IN1(EAX[31]), .IN2(n4442), .Q(N1753) );
  AO21X1 U4643 ( .IN1(n4444), .IN2(n4445), .IN3(n4443), .Q(n4514) );
  AOI22X1 U4644 ( .IN1(n4445), .IN2(READY_n), .IN3(n4518), .IN4(n4514), .QN(
        n4448) );
  NAND4X0 U4645 ( .IN1(n4448), .IN2(n4447), .IN3(n4468), .IN4(n4446), .QN(
        n4452) );
  INVX0 U4646 ( .INP(n4516), .ZN(n4525) );
  NAND2X0 U4647 ( .IN1(n4525), .IN2(n4469), .QN(n4449) );
  NAND4X0 U4648 ( .IN1(n4450), .IN2(n4488), .IN3(n4468), .IN4(n4449), .QN(
        n4451) );
  MUX21X1 U4649 ( .IN1(RequestPending), .IN2(n4452), .S(n4451), .Q(n2077) );
  NAND2X0 U4650 ( .IN1(State[1]), .IN2(HOLD), .QN(n4453) );
  NAND2X0 U4651 ( .IN1(RequestPending), .IN2(n4453), .QN(n4457) );
  AOI22X1 U4652 ( .IN1(HOLD), .IN2(State[2]), .IN3(NA_n), .IN4(n5202), .QN(
        n4454) );
  NAND2X0 U4653 ( .IN1(RequestPending), .IN2(n4454), .QN(n4456) );
  NAND2X0 U4654 ( .IN1(State[0]), .IN2(n4460), .QN(n4455) );
  AO222X1 U4655 ( .IN1(n4457), .IN2(State[0]), .IN3(n5178), .IN4(n4456), .IN5(
        n4455), .IN6(n5207), .Q(n2076) );
  INVX0 U4656 ( .INP(HOLD), .ZN(n4458) );
  AO222X1 U4657 ( .IN1(n4459), .IN2(n5178), .IN3(n4459), .IN4(n4458), .IN5(
        HOLD), .IN6(State[2]), .Q(n4461) );
  NAND3X0 U4658 ( .IN1(n4518), .IN2(n4461), .IN3(n4460), .QN(n2075) );
  NOR2X0 U4659 ( .IN1(State[1]), .IN2(n4462), .QN(n4463) );
  NOR3X0 U4660 ( .IN1(n5202), .IN2(n5178), .IN3(State[2]), .QN(n4464) );
  NOR2X0 U4661 ( .IN1(n4463), .IN2(n4464), .QN(n5166) );
  AO21X1 U4662 ( .IN1(n5178), .IN2(n5202), .IN3(n4464), .Q(n5169) );
  NOR2X0 U4663 ( .IN1(State[0]), .IN2(n4465), .QN(n5167) );
  AO21X1 U4664 ( .IN1(BS16_n), .IN2(n5169), .IN3(n5167), .Q(n5165) );
  AO21X1 U4665 ( .IN1(StateBS16), .IN2(n5166), .IN3(n5165), .Q(n2073) );
  NAND2X0 U4666 ( .IN1(n4474), .IN2(State2[3]), .QN(n4467) );
  NAND3X0 U4667 ( .IN1(n4467), .IN2(n4466), .IN3(n4485), .QN(n2072) );
  NOR3X0 U4668 ( .IN1(n5176), .IN2(n4469), .IN3(State2[2]), .QN(n4475) );
  NOR2X0 U4669 ( .IN1(State2[1]), .IN2(n4468), .QN(n4476) );
  NAND2X0 U4670 ( .IN1(n4476), .IN2(n4469), .QN(n4471) );
  NAND3X0 U4671 ( .IN1(n4471), .IN2(n4519), .IN3(n4470), .QN(n4472) );
  AO222X1 U4672 ( .IN1(State2[1]), .IN2(n4475), .IN3(State2[1]), .IN4(n4474), 
        .IN5(n4473), .IN6(n4472), .Q(n2067) );
  AO21X1 U4673 ( .IN1(CodeFetch), .IN2(n4488), .IN3(n4476), .Q(n2034) );
  OA21X1 U4674 ( .IN1(Flush), .IN2(n4493), .IN3(n4495), .Q(n4477) );
  NOR2X0 U4675 ( .IN1(n5094), .IN2(n4477), .QN(n4497) );
  INVX0 U4676 ( .INP(n4497), .ZN(n4499) );
  OA21X1 U4677 ( .IN1(n4604), .IN2(n4485), .IN3(n4499), .Q(n4513) );
  INVX0 U4678 ( .INP(n4849), .ZN(n4890) );
  NOR2X0 U4679 ( .IN1(N4186), .IN2(n5198), .QN(n4726) );
  NAND2X0 U4680 ( .IN1(n4604), .IN2(n4726), .QN(n4893) );
  NAND4X0 U4681 ( .IN1(StateBS16), .IN2(n4977), .IN3(N4187), .IN4(n5182), .QN(
        n4482) );
  NAND3X0 U4682 ( .IN1(N4187), .IN2(StateBS16), .IN3(n5182), .QN(n4478) );
  NAND2X0 U4683 ( .IN1(n4977), .IN2(n4478), .QN(n4502) );
  AND2X1 U4684 ( .IN1(n4479), .IN2(n4502), .Q(n4505) );
  OA21X1 U4685 ( .IN1(N4186), .IN2(n4504), .IN3(n4480), .Q(n4481) );
  MUX21X1 U4686 ( .IN1(n4482), .IN2(n4505), .S(n4481), .Q(n4483) );
  OA21X1 U4687 ( .IN1(n4485), .IN2(n4893), .IN3(n4483), .Q(n4484) );
  OAI221X1 U4688 ( .IN1(n4513), .IN2(n5200), .IN3(n4485), .IN4(n4890), .IN5(
        n4484), .QN(n2033) );
  INVX0 U4689 ( .INP(n4488), .ZN(n4490) );
  AO221X1 U4690 ( .IN1(n4490), .IN2(n4486), .IN3(n4488), .IN4(MemoryFetch), 
        .IN5(n4487), .Q(n2032) );
  AO221X1 U4691 ( .IN1(n4490), .IN2(n4489), .IN3(n4488), .IN4(ReadRequest), 
        .IN5(n4487), .Q(n2031) );
  MUX21X1 U4692 ( .IN1(Flush), .IN2(n4492), .S(n4491), .Q(n2030) );
  INVX0 U4693 ( .INP(n4493), .ZN(n4494) );
  AO22X1 U4694 ( .IN1(n4495), .IN2(n4494), .IN3(n5016), .IN4(n5199), .Q(n4496)
         );
  AO222X1 U4695 ( .IN1(N1351), .IN2(n4497), .IN3(N1351), .IN4(n5096), .IN5(
        n4499), .IN6(n4496), .Q(n2024) );
  NAND2X0 U4696 ( .IN1(n5016), .IN2(n5199), .QN(n4498) );
  NAND3X0 U4697 ( .IN1(n5020), .IN2(n4499), .IN3(n4498), .QN(n4501) );
  AO22X1 U4698 ( .IN1(n4848), .IN2(n5016), .IN3(n4255), .IN4(n5182), .Q(n4500)
         );
  AO21X1 U4699 ( .IN1(N4188), .IN2(n4501), .IN3(n4500), .Q(n2023) );
  NAND2X0 U4701 ( .IN1(StateBS16), .IN2(n5182), .QN(n4503) );
  NOR2X0 U4702 ( .IN1(n4503), .IN2(n4502), .QN(n4511) );
  NAND3X0 U4703 ( .IN1(n4604), .IN2(n5016), .IN3(n5198), .QN(n4509) );
  NOR2X0 U4704 ( .IN1(n4505), .IN2(n4504), .QN(n4507) );
  NAND2X0 U4705 ( .IN1(n5198), .IN2(n5182), .QN(n4506) );
  NAND2X0 U4706 ( .IN1(n4507), .IN2(n4506), .QN(n4508) );
  NAND2X0 U4707 ( .IN1(n4509), .IN2(n4508), .QN(n4510) );
  NOR2X0 U4708 ( .IN1(n4511), .IN2(n4510), .QN(n4512) );
  OAI21X1 U4709 ( .IN1(n4513), .IN2(n5198), .IN3(n4512), .QN(n2022) );
  NAND2X0 U4710 ( .IN1(n4515), .IN2(n4514), .QN(n4517) );
  OA21X1 U4711 ( .IN1(n4518), .IN2(n4517), .IN3(n4516), .Q(n4522) );
  NOR2X0 U4712 ( .IN1(n4522), .IN2(n4519), .QN(n4520) );
  AO222X1 U4713 ( .IN1(n4525), .IN2(\C1/DATA2_0 ), .IN3(EAX[0]), .IN4(n4520), 
        .IN5(n4522), .IN6(Datao[0]), .Q(n1927) );
  AO222X1 U4714 ( .IN1(n4525), .IN2(\C1/DATA2_1 ), .IN3(EAX[1]), .IN4(n4520), 
        .IN5(n4522), .IN6(Datao[1]), .Q(n1926) );
  AO222X1 U4715 ( .IN1(n4525), .IN2(\C1/DATA2_2 ), .IN3(EAX[2]), .IN4(n4520), 
        .IN5(n4522), .IN6(Datao[2]), .Q(n1925) );
  AO222X1 U4716 ( .IN1(n4525), .IN2(\C1/DATA2_3 ), .IN3(EAX[3]), .IN4(n4520), 
        .IN5(n4522), .IN6(Datao[3]), .Q(n1924) );
  AO222X1 U4717 ( .IN1(n4525), .IN2(\C1/DATA2_4 ), .IN3(EAX[4]), .IN4(n4520), 
        .IN5(n4522), .IN6(Datao[4]), .Q(n1923) );
  AO222X1 U4718 ( .IN1(n4525), .IN2(\C1/DATA2_5 ), .IN3(EAX[5]), .IN4(n4520), 
        .IN5(n4522), .IN6(Datao[5]), .Q(n1922) );
  AO222X1 U4719 ( .IN1(n4525), .IN2(\C1/DATA2_6 ), .IN3(EAX[6]), .IN4(n4520), 
        .IN5(n4522), .IN6(Datao[6]), .Q(n1921) );
  AO222X1 U4720 ( .IN1(n4525), .IN2(\C1/DATA2_7 ), .IN3(EAX[7]), .IN4(n4520), 
        .IN5(n4522), .IN6(Datao[7]), .Q(n1920) );
  AO222X1 U4721 ( .IN1(n4525), .IN2(\C1/DATA2_8 ), .IN3(EAX[8]), .IN4(n4520), 
        .IN5(n4522), .IN6(Datao[8]), .Q(n1919) );
  AO222X1 U4722 ( .IN1(n4525), .IN2(\C1/DATA2_9 ), .IN3(EAX[9]), .IN4(n4520), 
        .IN5(n4522), .IN6(Datao[9]), .Q(n1918) );
  AO222X1 U4723 ( .IN1(n4525), .IN2(\C1/DATA2_10 ), .IN3(EAX[10]), .IN4(n4520), 
        .IN5(n4522), .IN6(Datao[10]), .Q(n1917) );
  AO222X1 U4724 ( .IN1(n4525), .IN2(\C1/DATA2_11 ), .IN3(EAX[11]), .IN4(n4520), 
        .IN5(n4522), .IN6(Datao[11]), .Q(n1916) );
  AO222X1 U4725 ( .IN1(n4525), .IN2(\C1/DATA2_12 ), .IN3(EAX[12]), .IN4(n4520), 
        .IN5(n4522), .IN6(Datao[12]), .Q(n1915) );
  AO222X1 U4726 ( .IN1(n4525), .IN2(\C1/DATA2_13 ), .IN3(EAX[13]), .IN4(n4520), 
        .IN5(n4522), .IN6(Datao[13]), .Q(n1914) );
  AO222X1 U4727 ( .IN1(n4525), .IN2(\C1/DATA2_14 ), .IN3(EAX[14]), .IN4(n4520), 
        .IN5(n4522), .IN6(Datao[14]), .Q(n1913) );
  AO222X1 U4728 ( .IN1(n4525), .IN2(\C1/DATA2_15 ), .IN3(EAX[15]), .IN4(n4520), 
        .IN5(n4522), .IN6(Datao[15]), .Q(n1912) );
  NOR2X0 U4729 ( .IN1(n4522), .IN2(n4521), .QN(n4523) );
  AO222X1 U4730 ( .IN1(n4525), .IN2(\C1/DATA2_16 ), .IN3(\C1/DATA1_16 ), .IN4(
        n4523), .IN5(n4522), .IN6(Datao[16]), .Q(n1911) );
  AO222X1 U4731 ( .IN1(n4525), .IN2(\C1/DATA2_17 ), .IN3(\C1/DATA1_17 ), .IN4(
        n4523), .IN5(n4522), .IN6(Datao[17]), .Q(n1910) );
  AO222X1 U4732 ( .IN1(n4525), .IN2(\C1/DATA2_18 ), .IN3(\C1/DATA1_18 ), .IN4(
        n4523), .IN5(n4522), .IN6(Datao[18]), .Q(n1909) );
  AO222X1 U4733 ( .IN1(n4525), .IN2(\C1/DATA2_19 ), .IN3(\C1/DATA1_19 ), .IN4(
        n4523), .IN5(n4522), .IN6(Datao[19]), .Q(n1908) );
  AO222X1 U4734 ( .IN1(n4525), .IN2(\C1/DATA2_20 ), .IN3(\C1/DATA1_20 ), .IN4(
        n4523), .IN5(n4522), .IN6(Datao[20]), .Q(n1907) );
  AO222X1 U4735 ( .IN1(n4525), .IN2(\C1/DATA2_21 ), .IN3(\C1/DATA1_21 ), .IN4(
        n4523), .IN5(n4522), .IN6(Datao[21]), .Q(n1906) );
  AO222X1 U4736 ( .IN1(n4525), .IN2(\C1/DATA2_22 ), .IN3(\C1/DATA1_22 ), .IN4(
        n4523), .IN5(n4522), .IN6(Datao[22]), .Q(n1905) );
  AO222X1 U4737 ( .IN1(n4525), .IN2(\C1/DATA2_23 ), .IN3(\C1/DATA1_23 ), .IN4(
        n4523), .IN5(n4522), .IN6(Datao[23]), .Q(n1904) );
  AO222X1 U4738 ( .IN1(n4525), .IN2(\C1/DATA2_24 ), .IN3(\C1/DATA1_24 ), .IN4(
        n4523), .IN5(n4522), .IN6(Datao[24]), .Q(n1903) );
  AO222X1 U4739 ( .IN1(n4525), .IN2(\C1/DATA2_25 ), .IN3(\C1/DATA1_25 ), .IN4(
        n4523), .IN5(n4522), .IN6(Datao[25]), .Q(n1902) );
  AO222X1 U4740 ( .IN1(n4525), .IN2(\C1/DATA2_26 ), .IN3(\C1/DATA1_26 ), .IN4(
        n4523), .IN5(n4522), .IN6(Datao[26]), .Q(n1901) );
  AO222X1 U4741 ( .IN1(n4525), .IN2(\C1/DATA2_27 ), .IN3(\C1/DATA1_27 ), .IN4(
        n4523), .IN5(n4522), .IN6(Datao[27]), .Q(n1900) );
  AO222X1 U4742 ( .IN1(n4525), .IN2(\C1/DATA2_28 ), .IN3(\C1/DATA1_28 ), .IN4(
        n4523), .IN5(n4522), .IN6(Datao[28]), .Q(n1899) );
  AO222X1 U4743 ( .IN1(n4525), .IN2(\C1/DATA2_29 ), .IN3(\C1/DATA1_29 ), .IN4(
        n4523), .IN5(n4522), .IN6(Datao[29]), .Q(n1898) );
  AO222X1 U4744 ( .IN1(n4525), .IN2(\C1/DATA2_30 ), .IN3(n4524), .IN4(n4523), 
        .IN5(n4522), .IN6(Datao[30]), .Q(n1897) );
  NAND2X0 U4745 ( .IN1(n4605), .IN2(n4848), .QN(n4648) );
  OA22X1 U4746 ( .IN1(n4972), .IN2(n4648), .IN3(n4973), .IN4(n4608), .Q(n4526)
         );
  NOR2X0 U4747 ( .IN1(n5020), .IN2(n4566), .QN(n4557) );
  INVX0 U4748 ( .INP(n4557), .ZN(n4564) );
  NAND3X0 U4749 ( .IN1(n4526), .IN2(n4556), .IN3(n4564), .QN(n4547) );
  INVX0 U4750 ( .INP(n4547), .ZN(n4559) );
  OA22X1 U4751 ( .IN1(n4559), .IN2(n5105), .IN3(n5100), .IN4(n4556), .Q(n4530)
         );
  NOR4X0 U4752 ( .IN1(n5101), .IN2(n5095), .IN3(n5097), .IN4(n4559), .QN(n4558) );
  NAND2X0 U4753 ( .IN1(Datai[0]), .IN2(n4558), .QN(n4529) );
  NAND2X0 U4754 ( .IN1(\InstQueue[1][0] ), .IN2(n4559), .QN(n4528) );
  NAND2X0 U4755 ( .IN1(n4557), .IN2(n5108), .QN(n4527) );
  NAND4X0 U4756 ( .IN1(n4530), .IN2(n4529), .IN3(n4528), .IN4(n4527), .QN(
        n1856) );
  INVX0 U4757 ( .INP(n5068), .ZN(n5113) );
  OA22X1 U4758 ( .IN1(n4559), .IN2(n5113), .IN3(n5112), .IN4(n4556), .Q(n4534)
         );
  NAND2X0 U4759 ( .IN1(Datai[1]), .IN2(n4558), .QN(n4533) );
  NAND2X0 U4760 ( .IN1(\InstQueue[1][1] ), .IN2(n4559), .QN(n4532) );
  INVX0 U4761 ( .INP(n5063), .ZN(n5114) );
  NAND2X0 U4762 ( .IN1(n4557), .IN2(n5114), .QN(n4531) );
  NAND4X0 U4763 ( .IN1(n4534), .IN2(n4533), .IN3(n4532), .IN4(n4531), .QN(
        n1855) );
  OA22X1 U4764 ( .IN1(n4559), .IN2(n5120), .IN3(n5119), .IN4(n4556), .Q(n4538)
         );
  NAND2X0 U4765 ( .IN1(n4557), .IN2(n5121), .QN(n4537) );
  NAND2X0 U4766 ( .IN1(\InstQueue[1][2] ), .IN2(n4559), .QN(n4536) );
  NAND2X0 U4767 ( .IN1(Datai[2]), .IN2(n4558), .QN(n4535) );
  NAND4X0 U4768 ( .IN1(n4538), .IN2(n4537), .IN3(n4536), .IN4(n4535), .QN(
        n1854) );
  OA22X1 U4769 ( .IN1(n4559), .IN2(n5127), .IN3(n5126), .IN4(n4556), .Q(n4542)
         );
  NAND2X0 U4770 ( .IN1(n4557), .IN2(n5128), .QN(n4541) );
  NAND2X0 U4771 ( .IN1(\InstQueue[1][3] ), .IN2(n4559), .QN(n4540) );
  NAND2X0 U4772 ( .IN1(Datai[3]), .IN2(n4558), .QN(n4539) );
  NAND4X0 U4773 ( .IN1(n4542), .IN2(n4541), .IN3(n4540), .IN4(n4539), .QN(
        n1853) );
  OA22X1 U4774 ( .IN1(n4559), .IN2(n5134), .IN3(n5133), .IN4(n4556), .Q(n4546)
         );
  NAND2X0 U4775 ( .IN1(n4557), .IN2(n5135), .QN(n4545) );
  NAND2X0 U4776 ( .IN1(Datai[4]), .IN2(n4558), .QN(n4544) );
  NAND2X0 U4777 ( .IN1(\InstQueue[1][4] ), .IN2(n4559), .QN(n4543) );
  NAND4X0 U4778 ( .IN1(n4546), .IN2(n4545), .IN3(n4544), .IN4(n4543), .QN(
        n1852) );
  OA22X1 U4779 ( .IN1(n4564), .IN2(n5042), .IN3(n4556), .IN4(n5140), .Q(n4551)
         );
  NAND2X0 U4780 ( .IN1(n4547), .IN2(n5041), .QN(n4550) );
  NAND2X0 U4781 ( .IN1(Datai[5]), .IN2(n4558), .QN(n4549) );
  NAND2X0 U4782 ( .IN1(\InstQueue[1][5] ), .IN2(n4559), .QN(n4548) );
  NAND4X0 U4783 ( .IN1(n4551), .IN2(n4550), .IN3(n4549), .IN4(n4548), .QN(
        n1851) );
  OA22X1 U4784 ( .IN1(n4559), .IN2(n5148), .IN3(n5147), .IN4(n4556), .Q(n4555)
         );
  NAND2X0 U4785 ( .IN1(n4557), .IN2(n5149), .QN(n4554) );
  NAND2X0 U4786 ( .IN1(Datai[6]), .IN2(n4558), .QN(n4553) );
  NAND2X0 U4787 ( .IN1(\InstQueue[1][6] ), .IN2(n4559), .QN(n4552) );
  NAND4X0 U4788 ( .IN1(n4555), .IN2(n4554), .IN3(n4553), .IN4(n4552), .QN(
        n1850) );
  OA22X1 U4789 ( .IN1(n5156), .IN2(n4559), .IN3(n5155), .IN4(n4556), .Q(n4563)
         );
  NAND2X0 U4790 ( .IN1(n5158), .IN2(n4557), .QN(n4562) );
  NAND2X0 U4791 ( .IN1(Datai[7]), .IN2(n4558), .QN(n4561) );
  NAND2X0 U4792 ( .IN1(\InstQueue[1][7] ), .IN2(n4559), .QN(n4560) );
  NAND4X0 U4793 ( .IN1(n4563), .IN2(n4562), .IN3(n4561), .IN4(n4560), .QN(
        n1849) );
  NAND3X0 U4794 ( .IN1(n4605), .IN2(N4188), .IN3(n5199), .QN(n4688) );
  OA22X1 U4795 ( .IN1(n4972), .IN2(n4688), .IN3(n4973), .IN4(n4648), .Q(n4565)
         );
  NOR2X0 U4796 ( .IN1(n5020), .IN2(n4608), .QN(n4597) );
  INVX0 U4797 ( .INP(n4597), .ZN(n4606) );
  NAND3X0 U4798 ( .IN1(n4565), .IN2(n4564), .IN3(n4606), .QN(n4587) );
  INVX0 U4799 ( .INP(n4587), .ZN(n4599) );
  NAND2X0 U4800 ( .IN1(n5095), .IN2(n4587), .QN(n4596) );
  OA22X1 U4801 ( .IN1(n4599), .IN2(n5105), .IN3(n5100), .IN4(n4596), .Q(n4570)
         );
  AND4X1 U4802 ( .IN1(n4977), .IN2(n4566), .IN3(n4608), .IN4(n4587), .Q(n4598)
         );
  NAND2X0 U4803 ( .IN1(Datai[0]), .IN2(n4598), .QN(n4569) );
  NAND2X0 U4804 ( .IN1(\InstQueue[2][0] ), .IN2(n4599), .QN(n4568) );
  NAND2X0 U4805 ( .IN1(n4597), .IN2(n5108), .QN(n4567) );
  NAND4X0 U4806 ( .IN1(n4570), .IN2(n4569), .IN3(n4568), .IN4(n4567), .QN(
        n1848) );
  OA22X1 U4807 ( .IN1(n4599), .IN2(n5113), .IN3(n5112), .IN4(n4596), .Q(n4574)
         );
  NAND2X0 U4808 ( .IN1(Datai[1]), .IN2(n4598), .QN(n4573) );
  NAND2X0 U4809 ( .IN1(\InstQueue[2][1] ), .IN2(n4599), .QN(n4572) );
  NAND2X0 U4810 ( .IN1(n4597), .IN2(n5114), .QN(n4571) );
  NAND4X0 U4811 ( .IN1(n4574), .IN2(n4573), .IN3(n4572), .IN4(n4571), .QN(
        n1847) );
  OA22X1 U4812 ( .IN1(n4599), .IN2(n5120), .IN3(n5119), .IN4(n4596), .Q(n4578)
         );
  NAND2X0 U4813 ( .IN1(n4597), .IN2(n5121), .QN(n4577) );
  NAND2X0 U4814 ( .IN1(\InstQueue[2][2] ), .IN2(n4599), .QN(n4576) );
  NAND2X0 U4815 ( .IN1(Datai[2]), .IN2(n4598), .QN(n4575) );
  NAND4X0 U4816 ( .IN1(n4578), .IN2(n4577), .IN3(n4576), .IN4(n4575), .QN(
        n1846) );
  OA22X1 U4817 ( .IN1(n4599), .IN2(n5127), .IN3(n5126), .IN4(n4596), .Q(n4582)
         );
  NAND2X0 U4818 ( .IN1(n4597), .IN2(n5128), .QN(n4581) );
  NAND2X0 U4819 ( .IN1(\InstQueue[2][3] ), .IN2(n4599), .QN(n4580) );
  NAND2X0 U4820 ( .IN1(Datai[3]), .IN2(n4598), .QN(n4579) );
  NAND4X0 U4821 ( .IN1(n4582), .IN2(n4581), .IN3(n4580), .IN4(n4579), .QN(
        n1845) );
  OA22X1 U4822 ( .IN1(n4599), .IN2(n5134), .IN3(n5133), .IN4(n4596), .Q(n4586)
         );
  NAND2X0 U4823 ( .IN1(n4597), .IN2(n5135), .QN(n4585) );
  NAND2X0 U4824 ( .IN1(Datai[4]), .IN2(n4598), .QN(n4584) );
  NAND2X0 U4825 ( .IN1(\InstQueue[2][4] ), .IN2(n4599), .QN(n4583) );
  NAND4X0 U4826 ( .IN1(n4586), .IN2(n4585), .IN3(n4584), .IN4(n4583), .QN(
        n1844) );
  OA22X1 U4827 ( .IN1(n4606), .IN2(n5042), .IN3(n4596), .IN4(n5140), .Q(n4591)
         );
  NAND2X0 U4828 ( .IN1(n4587), .IN2(n5041), .QN(n4590) );
  NAND2X0 U4829 ( .IN1(Datai[5]), .IN2(n4598), .QN(n4589) );
  NAND2X0 U4830 ( .IN1(\InstQueue[2][5] ), .IN2(n4599), .QN(n4588) );
  NAND4X0 U4831 ( .IN1(n4591), .IN2(n4590), .IN3(n4589), .IN4(n4588), .QN(
        n1843) );
  OA22X1 U4832 ( .IN1(n4599), .IN2(n5148), .IN3(n5147), .IN4(n4596), .Q(n4595)
         );
  NAND2X0 U4833 ( .IN1(n4597), .IN2(n5149), .QN(n4594) );
  NAND2X0 U4834 ( .IN1(Datai[6]), .IN2(n4598), .QN(n4593) );
  NAND2X0 U4835 ( .IN1(\InstQueue[2][6] ), .IN2(n4599), .QN(n4592) );
  NAND4X0 U4836 ( .IN1(n4595), .IN2(n4594), .IN3(n4593), .IN4(n4592), .QN(
        n1842) );
  OA22X1 U4837 ( .IN1(n5156), .IN2(n4599), .IN3(n5155), .IN4(n4596), .Q(n4603)
         );
  NAND2X0 U4838 ( .IN1(n5158), .IN2(n4597), .QN(n4602) );
  NAND2X0 U4839 ( .IN1(Datai[7]), .IN2(n4598), .QN(n4601) );
  NAND2X0 U4840 ( .IN1(\InstQueue[2][7] ), .IN2(n4599), .QN(n4600) );
  NAND4X0 U4841 ( .IN1(n4603), .IN2(n4602), .IN3(n4601), .IN4(n4600), .QN(
        n1841) );
  NAND2X0 U4842 ( .IN1(n4605), .IN2(n4604), .QN(n4729) );
  OA22X1 U4843 ( .IN1(n4972), .IN2(n4729), .IN3(n4973), .IN4(n4688), .Q(n4607)
         );
  NOR2X0 U4844 ( .IN1(n5020), .IN2(n4648), .QN(n4639) );
  INVX0 U4845 ( .INP(n4639), .ZN(n4646) );
  NAND3X0 U4846 ( .IN1(n4607), .IN2(n4606), .IN3(n4646), .QN(n4629) );
  INVX0 U4847 ( .INP(n4629), .ZN(n4641) );
  OR2X1 U4848 ( .IN1(n4608), .IN2(n4641), .Q(n4638) );
  OA22X1 U4849 ( .IN1(n4641), .IN2(n5105), .IN3(n5100), .IN4(n4638), .Q(n4612)
         );
  AND4X1 U4850 ( .IN1(n4977), .IN2(n4648), .IN3(n4608), .IN4(n4629), .Q(n4640)
         );
  NAND2X0 U4851 ( .IN1(Datai[0]), .IN2(n4640), .QN(n4611) );
  NAND2X0 U4852 ( .IN1(\InstQueue[3][0] ), .IN2(n4641), .QN(n4610) );
  NAND2X0 U4853 ( .IN1(n4639), .IN2(n5108), .QN(n4609) );
  NAND4X0 U4854 ( .IN1(n4612), .IN2(n4611), .IN3(n4610), .IN4(n4609), .QN(
        n1840) );
  OA22X1 U4855 ( .IN1(n4641), .IN2(n5113), .IN3(n5112), .IN4(n4638), .Q(n4616)
         );
  NAND2X0 U4856 ( .IN1(Datai[1]), .IN2(n4640), .QN(n4615) );
  NAND2X0 U4857 ( .IN1(\InstQueue[3][1] ), .IN2(n4641), .QN(n4614) );
  NAND2X0 U4858 ( .IN1(n4639), .IN2(n5114), .QN(n4613) );
  NAND4X0 U4859 ( .IN1(n4616), .IN2(n4615), .IN3(n4614), .IN4(n4613), .QN(
        n1839) );
  OA22X1 U4860 ( .IN1(n4641), .IN2(n5120), .IN3(n5119), .IN4(n4638), .Q(n4620)
         );
  NAND2X0 U4861 ( .IN1(n4639), .IN2(n5121), .QN(n4619) );
  NAND2X0 U4862 ( .IN1(\InstQueue[3][2] ), .IN2(n4641), .QN(n4618) );
  NAND2X0 U4863 ( .IN1(Datai[2]), .IN2(n4640), .QN(n4617) );
  NAND4X0 U4864 ( .IN1(n4620), .IN2(n4619), .IN3(n4618), .IN4(n4617), .QN(
        n1838) );
  OA22X1 U4865 ( .IN1(n4641), .IN2(n5127), .IN3(n5126), .IN4(n4638), .Q(n4624)
         );
  NAND2X0 U4866 ( .IN1(n4639), .IN2(n5128), .QN(n4623) );
  NAND2X0 U4867 ( .IN1(\InstQueue[3][3] ), .IN2(n4641), .QN(n4622) );
  NAND2X0 U4868 ( .IN1(Datai[3]), .IN2(n4640), .QN(n4621) );
  NAND4X0 U4869 ( .IN1(n4624), .IN2(n4623), .IN3(n4622), .IN4(n4621), .QN(
        n1837) );
  OA22X1 U4870 ( .IN1(n4641), .IN2(n5134), .IN3(n5133), .IN4(n4638), .Q(n4628)
         );
  NAND2X0 U4871 ( .IN1(n4639), .IN2(n5135), .QN(n4627) );
  NAND2X0 U4872 ( .IN1(Datai[4]), .IN2(n4640), .QN(n4626) );
  NAND2X0 U4873 ( .IN1(\InstQueue[3][4] ), .IN2(n4641), .QN(n4625) );
  NAND4X0 U4874 ( .IN1(n4628), .IN2(n4627), .IN3(n4626), .IN4(n4625), .QN(
        n1836) );
  OA22X1 U4875 ( .IN1(n4646), .IN2(n5042), .IN3(n4638), .IN4(n5140), .Q(n4633)
         );
  NAND2X0 U4876 ( .IN1(n4629), .IN2(n5041), .QN(n4632) );
  NAND2X0 U4877 ( .IN1(Datai[5]), .IN2(n4640), .QN(n4631) );
  NAND2X0 U4878 ( .IN1(\InstQueue[3][5] ), .IN2(n4641), .QN(n4630) );
  NAND4X0 U4879 ( .IN1(n4633), .IN2(n4632), .IN3(n4631), .IN4(n4630), .QN(
        n1835) );
  OA22X1 U4880 ( .IN1(n4641), .IN2(n5148), .IN3(n5147), .IN4(n4638), .Q(n4637)
         );
  NAND2X0 U4881 ( .IN1(n4639), .IN2(n5149), .QN(n4636) );
  NAND2X0 U4882 ( .IN1(Datai[6]), .IN2(n4640), .QN(n4635) );
  NAND2X0 U4883 ( .IN1(\InstQueue[3][6] ), .IN2(n4641), .QN(n4634) );
  NAND4X0 U4884 ( .IN1(n4637), .IN2(n4636), .IN3(n4635), .IN4(n4634), .QN(
        n1834) );
  OA22X1 U4885 ( .IN1(n5156), .IN2(n4641), .IN3(n5155), .IN4(n4638), .Q(n4645)
         );
  NAND2X0 U4886 ( .IN1(n5158), .IN2(n4639), .QN(n4644) );
  NAND2X0 U4887 ( .IN1(Datai[7]), .IN2(n4640), .QN(n4643) );
  NAND2X0 U4888 ( .IN1(\InstQueue[3][7] ), .IN2(n4641), .QN(n4642) );
  NAND4X0 U4889 ( .IN1(n4645), .IN2(n4644), .IN3(n4643), .IN4(n4642), .QN(
        n1833) );
  NAND2X0 U4890 ( .IN1(n4807), .IN2(n4726), .QN(n4769) );
  OA22X1 U4891 ( .IN1(n4972), .IN2(n4769), .IN3(n4973), .IN4(n4729), .Q(n4647)
         );
  NOR2X0 U4892 ( .IN1(n5020), .IN2(n4688), .QN(n4679) );
  INVX0 U4893 ( .INP(n4679), .ZN(n4686) );
  NAND3X0 U4894 ( .IN1(n4647), .IN2(n4646), .IN3(n4686), .QN(n4669) );
  INVX0 U4895 ( .INP(n4669), .ZN(n4681) );
  OR2X1 U4896 ( .IN1(n4648), .IN2(n4681), .Q(n4678) );
  OA22X1 U4897 ( .IN1(n4681), .IN2(n5105), .IN3(n5100), .IN4(n4678), .Q(n4652)
         );
  AND4X1 U4898 ( .IN1(n4977), .IN2(n4688), .IN3(n4648), .IN4(n4669), .Q(n4680)
         );
  NAND2X0 U4899 ( .IN1(Datai[0]), .IN2(n4680), .QN(n4651) );
  NAND2X0 U4900 ( .IN1(\InstQueue[4][0] ), .IN2(n4681), .QN(n4650) );
  NAND2X0 U4901 ( .IN1(n4679), .IN2(n5108), .QN(n4649) );
  NAND4X0 U4902 ( .IN1(n4652), .IN2(n4651), .IN3(n4650), .IN4(n4649), .QN(
        n1832) );
  OA22X1 U4903 ( .IN1(n4681), .IN2(n5113), .IN3(n5112), .IN4(n4678), .Q(n4656)
         );
  NAND2X0 U4904 ( .IN1(Datai[1]), .IN2(n4680), .QN(n4655) );
  NAND2X0 U4905 ( .IN1(\InstQueue[4][1] ), .IN2(n4681), .QN(n4654) );
  NAND2X0 U4906 ( .IN1(n4679), .IN2(n5114), .QN(n4653) );
  NAND4X0 U4907 ( .IN1(n4656), .IN2(n4655), .IN3(n4654), .IN4(n4653), .QN(
        n1831) );
  OA22X1 U4908 ( .IN1(n4681), .IN2(n5120), .IN3(n5119), .IN4(n4678), .Q(n4660)
         );
  NAND2X0 U4909 ( .IN1(n4679), .IN2(n5121), .QN(n4659) );
  NAND2X0 U4910 ( .IN1(\InstQueue[4][2] ), .IN2(n4681), .QN(n4658) );
  NAND2X0 U4911 ( .IN1(Datai[2]), .IN2(n4680), .QN(n4657) );
  NAND4X0 U4912 ( .IN1(n4660), .IN2(n4659), .IN3(n4658), .IN4(n4657), .QN(
        n1830) );
  OA22X1 U4913 ( .IN1(n4681), .IN2(n5127), .IN3(n5126), .IN4(n4678), .Q(n4664)
         );
  NAND2X0 U4914 ( .IN1(n4679), .IN2(n5128), .QN(n4663) );
  NAND2X0 U4915 ( .IN1(\InstQueue[4][3] ), .IN2(n4681), .QN(n4662) );
  NAND2X0 U4916 ( .IN1(Datai[3]), .IN2(n4680), .QN(n4661) );
  NAND4X0 U4917 ( .IN1(n4664), .IN2(n4663), .IN3(n4662), .IN4(n4661), .QN(
        n1829) );
  OA22X1 U4918 ( .IN1(n4681), .IN2(n5134), .IN3(n5133), .IN4(n4678), .Q(n4668)
         );
  NAND2X0 U4919 ( .IN1(n4679), .IN2(n5135), .QN(n4667) );
  NAND2X0 U4920 ( .IN1(Datai[4]), .IN2(n4680), .QN(n4666) );
  NAND2X0 U4921 ( .IN1(\InstQueue[4][4] ), .IN2(n4681), .QN(n4665) );
  NAND4X0 U4922 ( .IN1(n4668), .IN2(n4667), .IN3(n4666), .IN4(n4665), .QN(
        n1828) );
  OA22X1 U4923 ( .IN1(n4686), .IN2(n5042), .IN3(n4678), .IN4(n5140), .Q(n4673)
         );
  NAND2X0 U4924 ( .IN1(n4669), .IN2(n5041), .QN(n4672) );
  NAND2X0 U4925 ( .IN1(Datai[5]), .IN2(n4680), .QN(n4671) );
  NAND2X0 U4926 ( .IN1(\InstQueue[4][5] ), .IN2(n4681), .QN(n4670) );
  NAND4X0 U4927 ( .IN1(n4673), .IN2(n4672), .IN3(n4671), .IN4(n4670), .QN(
        n1827) );
  OA22X1 U4928 ( .IN1(n4681), .IN2(n5148), .IN3(n5147), .IN4(n4678), .Q(n4677)
         );
  NAND2X0 U4929 ( .IN1(n4679), .IN2(n5149), .QN(n4676) );
  NAND2X0 U4930 ( .IN1(Datai[6]), .IN2(n4680), .QN(n4675) );
  NAND2X0 U4931 ( .IN1(\InstQueue[4][6] ), .IN2(n4681), .QN(n4674) );
  NAND4X0 U4932 ( .IN1(n4677), .IN2(n4676), .IN3(n4675), .IN4(n4674), .QN(
        n1826) );
  OA22X1 U4933 ( .IN1(n5156), .IN2(n4681), .IN3(n5155), .IN4(n4678), .Q(n4685)
         );
  NAND2X0 U4934 ( .IN1(n5158), .IN2(n4679), .QN(n4684) );
  NAND2X0 U4935 ( .IN1(Datai[7]), .IN2(n4680), .QN(n4683) );
  NAND2X0 U4936 ( .IN1(\InstQueue[4][7] ), .IN2(n4681), .QN(n4682) );
  NAND4X0 U4937 ( .IN1(n4685), .IN2(n4684), .IN3(n4683), .IN4(n4682), .QN(
        n1825) );
  NAND2X0 U4938 ( .IN1(n4848), .IN2(n4726), .QN(n4810) );
  OA22X1 U4939 ( .IN1(n4972), .IN2(n4810), .IN3(n4973), .IN4(n4769), .Q(n4687)
         );
  NOR2X0 U4940 ( .IN1(n5020), .IN2(n4729), .QN(n4719) );
  INVX0 U4941 ( .INP(n4719), .ZN(n4727) );
  NAND3X0 U4942 ( .IN1(n4687), .IN2(n4686), .IN3(n4727), .QN(n4709) );
  INVX0 U4943 ( .INP(n4709), .ZN(n4721) );
  OR2X1 U4944 ( .IN1(n4688), .IN2(n4721), .Q(n4718) );
  OA22X1 U4945 ( .IN1(n4721), .IN2(n5105), .IN3(n5100), .IN4(n4718), .Q(n4692)
         );
  AND4X1 U4946 ( .IN1(n4977), .IN2(n4729), .IN3(n4688), .IN4(n4709), .Q(n4720)
         );
  NAND2X0 U4947 ( .IN1(Datai[0]), .IN2(n4720), .QN(n4691) );
  NAND2X0 U4948 ( .IN1(\InstQueue[5][0] ), .IN2(n4721), .QN(n4690) );
  NAND2X0 U4949 ( .IN1(n4719), .IN2(n5108), .QN(n4689) );
  NAND4X0 U4950 ( .IN1(n4692), .IN2(n4691), .IN3(n4690), .IN4(n4689), .QN(
        n1824) );
  OA22X1 U4951 ( .IN1(n4721), .IN2(n5113), .IN3(n5112), .IN4(n4718), .Q(n4696)
         );
  NAND2X0 U4952 ( .IN1(Datai[1]), .IN2(n4720), .QN(n4695) );
  NAND2X0 U4953 ( .IN1(\InstQueue[5][1] ), .IN2(n4721), .QN(n4694) );
  NAND2X0 U4954 ( .IN1(n4719), .IN2(n5114), .QN(n4693) );
  NAND4X0 U4955 ( .IN1(n4696), .IN2(n4695), .IN3(n4694), .IN4(n4693), .QN(
        n1823) );
  OA22X1 U4956 ( .IN1(n4721), .IN2(n5120), .IN3(n5119), .IN4(n4718), .Q(n4700)
         );
  NAND2X0 U4957 ( .IN1(n4719), .IN2(n5121), .QN(n4699) );
  NAND2X0 U4958 ( .IN1(\InstQueue[5][2] ), .IN2(n4721), .QN(n4698) );
  NAND2X0 U4959 ( .IN1(Datai[2]), .IN2(n4720), .QN(n4697) );
  NAND4X0 U4960 ( .IN1(n4700), .IN2(n4699), .IN3(n4698), .IN4(n4697), .QN(
        n1822) );
  OA22X1 U4961 ( .IN1(n4721), .IN2(n5127), .IN3(n5126), .IN4(n4718), .Q(n4704)
         );
  NAND2X0 U4962 ( .IN1(n4719), .IN2(n5128), .QN(n4703) );
  NAND2X0 U4963 ( .IN1(\InstQueue[5][3] ), .IN2(n4721), .QN(n4702) );
  NAND2X0 U4964 ( .IN1(Datai[3]), .IN2(n4720), .QN(n4701) );
  NAND4X0 U4965 ( .IN1(n4704), .IN2(n4703), .IN3(n4702), .IN4(n4701), .QN(
        n1821) );
  OA22X1 U4966 ( .IN1(n4721), .IN2(n5134), .IN3(n5133), .IN4(n4718), .Q(n4708)
         );
  NAND2X0 U4967 ( .IN1(n4719), .IN2(n5135), .QN(n4707) );
  NAND2X0 U4968 ( .IN1(Datai[4]), .IN2(n4720), .QN(n4706) );
  NAND2X0 U4969 ( .IN1(\InstQueue[5][4] ), .IN2(n4721), .QN(n4705) );
  NAND4X0 U4970 ( .IN1(n4708), .IN2(n4707), .IN3(n4706), .IN4(n4705), .QN(
        n1820) );
  OA22X1 U4971 ( .IN1(n4727), .IN2(n5042), .IN3(n4718), .IN4(n5140), .Q(n4713)
         );
  NAND2X0 U4972 ( .IN1(n4709), .IN2(n5041), .QN(n4712) );
  NAND2X0 U4973 ( .IN1(Datai[5]), .IN2(n4720), .QN(n4711) );
  NAND2X0 U4974 ( .IN1(\InstQueue[5][5] ), .IN2(n4721), .QN(n4710) );
  NAND4X0 U4975 ( .IN1(n4713), .IN2(n4712), .IN3(n4711), .IN4(n4710), .QN(
        n1819) );
  OA22X1 U4976 ( .IN1(n4721), .IN2(n5148), .IN3(n5147), .IN4(n4718), .Q(n4717)
         );
  NAND2X0 U4977 ( .IN1(n4719), .IN2(n5149), .QN(n4716) );
  NAND2X0 U4978 ( .IN1(Datai[6]), .IN2(n4720), .QN(n4715) );
  NAND2X0 U4979 ( .IN1(\InstQueue[5][6] ), .IN2(n4721), .QN(n4714) );
  NAND4X0 U4980 ( .IN1(n4717), .IN2(n4716), .IN3(n4715), .IN4(n4714), .QN(
        n1818) );
  OA22X1 U4981 ( .IN1(n5156), .IN2(n4721), .IN3(n5155), .IN4(n4718), .Q(n4725)
         );
  NAND2X0 U4982 ( .IN1(n5158), .IN2(n4719), .QN(n4724) );
  NAND2X0 U4983 ( .IN1(Datai[7]), .IN2(n4720), .QN(n4723) );
  NAND2X0 U4984 ( .IN1(\InstQueue[5][7] ), .IN2(n4721), .QN(n4722) );
  NAND4X0 U4985 ( .IN1(n4725), .IN2(n4724), .IN3(n4723), .IN4(n4722), .QN(
        n1817) );
  NAND3X0 U4986 ( .IN1(N4188), .IN2(n4726), .IN3(n5199), .QN(n4852) );
  OA22X1 U4987 ( .IN1(n4972), .IN2(n4852), .IN3(n4973), .IN4(n4810), .Q(n4728)
         );
  NOR2X0 U4988 ( .IN1(n5020), .IN2(n4769), .QN(n4760) );
  INVX0 U4989 ( .INP(n4760), .ZN(n4767) );
  NAND3X0 U4990 ( .IN1(n4728), .IN2(n4727), .IN3(n4767), .QN(n4750) );
  INVX0 U4991 ( .INP(n4750), .ZN(n4762) );
  OR2X1 U4992 ( .IN1(n4729), .IN2(n4762), .Q(n4759) );
  OA22X1 U4993 ( .IN1(n4762), .IN2(n5105), .IN3(n5100), .IN4(n4759), .Q(n4733)
         );
  AND4X1 U4994 ( .IN1(n4977), .IN2(n4769), .IN3(n4729), .IN4(n4750), .Q(n4761)
         );
  NAND2X0 U4995 ( .IN1(Datai[0]), .IN2(n4761), .QN(n4732) );
  NAND2X0 U4996 ( .IN1(\InstQueue[6][0] ), .IN2(n4762), .QN(n4731) );
  NAND2X0 U4997 ( .IN1(n4760), .IN2(n5108), .QN(n4730) );
  NAND4X0 U4998 ( .IN1(n4733), .IN2(n4732), .IN3(n4731), .IN4(n4730), .QN(
        n1816) );
  OA22X1 U4999 ( .IN1(n4762), .IN2(n5113), .IN3(n5112), .IN4(n4759), .Q(n4737)
         );
  NAND2X0 U5000 ( .IN1(Datai[1]), .IN2(n4761), .QN(n4736) );
  NAND2X0 U5001 ( .IN1(\InstQueue[6][1] ), .IN2(n4762), .QN(n4735) );
  NAND2X0 U5002 ( .IN1(n4760), .IN2(n5114), .QN(n4734) );
  NAND4X0 U5003 ( .IN1(n4737), .IN2(n4736), .IN3(n4735), .IN4(n4734), .QN(
        n1815) );
  OA22X1 U5004 ( .IN1(n4762), .IN2(n5120), .IN3(n5119), .IN4(n4759), .Q(n4741)
         );
  NAND2X0 U5005 ( .IN1(n4760), .IN2(n5121), .QN(n4740) );
  NAND2X0 U5006 ( .IN1(\InstQueue[6][2] ), .IN2(n4762), .QN(n4739) );
  NAND2X0 U5007 ( .IN1(Datai[2]), .IN2(n4761), .QN(n4738) );
  NAND4X0 U5008 ( .IN1(n4741), .IN2(n4740), .IN3(n4739), .IN4(n4738), .QN(
        n1814) );
  OA22X1 U5009 ( .IN1(n4762), .IN2(n5127), .IN3(n5126), .IN4(n4759), .Q(n4745)
         );
  NAND2X0 U5010 ( .IN1(n4760), .IN2(n5128), .QN(n4744) );
  NAND2X0 U5011 ( .IN1(\InstQueue[6][3] ), .IN2(n4762), .QN(n4743) );
  NAND2X0 U5012 ( .IN1(Datai[3]), .IN2(n4761), .QN(n4742) );
  NAND4X0 U5013 ( .IN1(n4745), .IN2(n4744), .IN3(n4743), .IN4(n4742), .QN(
        n1813) );
  OA22X1 U5014 ( .IN1(n4762), .IN2(n5134), .IN3(n5133), .IN4(n4759), .Q(n4749)
         );
  NAND2X0 U5015 ( .IN1(n4760), .IN2(n5135), .QN(n4748) );
  NAND2X0 U5016 ( .IN1(Datai[4]), .IN2(n4761), .QN(n4747) );
  NAND2X0 U5017 ( .IN1(\InstQueue[6][4] ), .IN2(n4762), .QN(n4746) );
  NAND4X0 U5018 ( .IN1(n4749), .IN2(n4748), .IN3(n4747), .IN4(n4746), .QN(
        n1812) );
  OA22X1 U5019 ( .IN1(n4767), .IN2(n5042), .IN3(n4759), .IN4(n5140), .Q(n4754)
         );
  NAND2X0 U5020 ( .IN1(n4750), .IN2(n5041), .QN(n4753) );
  NAND2X0 U5021 ( .IN1(Datai[5]), .IN2(n4761), .QN(n4752) );
  NAND2X0 U5022 ( .IN1(\InstQueue[6][5] ), .IN2(n4762), .QN(n4751) );
  NAND4X0 U5023 ( .IN1(n4754), .IN2(n4753), .IN3(n4752), .IN4(n4751), .QN(
        n1811) );
  OA22X1 U5024 ( .IN1(n4762), .IN2(n5148), .IN3(n5147), .IN4(n4759), .Q(n4758)
         );
  NAND2X0 U5025 ( .IN1(n4760), .IN2(n5149), .QN(n4757) );
  NAND2X0 U5026 ( .IN1(Datai[6]), .IN2(n4761), .QN(n4756) );
  NAND2X0 U5027 ( .IN1(\InstQueue[6][6] ), .IN2(n4762), .QN(n4755) );
  NAND4X0 U5028 ( .IN1(n4758), .IN2(n4757), .IN3(n4756), .IN4(n4755), .QN(
        n1810) );
  OA22X1 U5029 ( .IN1(n5156), .IN2(n4762), .IN3(n5155), .IN4(n4759), .Q(n4766)
         );
  NAND2X0 U5030 ( .IN1(n5158), .IN2(n4760), .QN(n4765) );
  NAND2X0 U5031 ( .IN1(Datai[7]), .IN2(n4761), .QN(n4764) );
  NAND2X0 U5032 ( .IN1(\InstQueue[6][7] ), .IN2(n4762), .QN(n4763) );
  NAND4X0 U5033 ( .IN1(n4766), .IN2(n4765), .IN3(n4764), .IN4(n4763), .QN(
        n1809) );
  OA22X1 U5034 ( .IN1(n4972), .IN2(n4893), .IN3(n4973), .IN4(n4852), .Q(n4768)
         );
  NOR2X0 U5035 ( .IN1(n5020), .IN2(n4810), .QN(n4800) );
  INVX0 U5036 ( .INP(n4800), .ZN(n4808) );
  NAND3X0 U5037 ( .IN1(n4768), .IN2(n4767), .IN3(n4808), .QN(n4790) );
  INVX0 U5038 ( .INP(n4790), .ZN(n4802) );
  OR2X1 U5039 ( .IN1(n4769), .IN2(n4802), .Q(n4799) );
  OA22X1 U5040 ( .IN1(n4802), .IN2(n5105), .IN3(n5100), .IN4(n4799), .Q(n4773)
         );
  AND4X1 U5041 ( .IN1(n4977), .IN2(n4810), .IN3(n4769), .IN4(n4790), .Q(n4801)
         );
  NAND2X0 U5042 ( .IN1(Datai[0]), .IN2(n4801), .QN(n4772) );
  NAND2X0 U5043 ( .IN1(\InstQueue[7][0] ), .IN2(n4802), .QN(n4771) );
  NAND2X0 U5044 ( .IN1(n4800), .IN2(n5108), .QN(n4770) );
  NAND4X0 U5045 ( .IN1(n4773), .IN2(n4772), .IN3(n4771), .IN4(n4770), .QN(
        n1808) );
  OA22X1 U5046 ( .IN1(n4802), .IN2(n5113), .IN3(n5112), .IN4(n4799), .Q(n4777)
         );
  NAND2X0 U5047 ( .IN1(Datai[1]), .IN2(n4801), .QN(n4776) );
  NAND2X0 U5048 ( .IN1(\InstQueue[7][1] ), .IN2(n4802), .QN(n4775) );
  NAND2X0 U5049 ( .IN1(n4800), .IN2(n5114), .QN(n4774) );
  NAND4X0 U5050 ( .IN1(n4777), .IN2(n4776), .IN3(n4775), .IN4(n4774), .QN(
        n1807) );
  OA22X1 U5051 ( .IN1(n4802), .IN2(n5120), .IN3(n5119), .IN4(n4799), .Q(n4781)
         );
  NAND2X0 U5052 ( .IN1(n4800), .IN2(n5121), .QN(n4780) );
  NAND2X0 U5053 ( .IN1(\InstQueue[7][2] ), .IN2(n4802), .QN(n4779) );
  NAND2X0 U5054 ( .IN1(Datai[2]), .IN2(n4801), .QN(n4778) );
  NAND4X0 U5055 ( .IN1(n4781), .IN2(n4780), .IN3(n4779), .IN4(n4778), .QN(
        n1806) );
  OA22X1 U5056 ( .IN1(n4802), .IN2(n5127), .IN3(n5126), .IN4(n4799), .Q(n4785)
         );
  NAND2X0 U5057 ( .IN1(n4800), .IN2(n5128), .QN(n4784) );
  NAND2X0 U5058 ( .IN1(\InstQueue[7][3] ), .IN2(n4802), .QN(n4783) );
  NAND2X0 U5059 ( .IN1(Datai[3]), .IN2(n4801), .QN(n4782) );
  NAND4X0 U5060 ( .IN1(n4785), .IN2(n4784), .IN3(n4783), .IN4(n4782), .QN(
        n1805) );
  OA22X1 U5061 ( .IN1(n4802), .IN2(n5134), .IN3(n5133), .IN4(n4799), .Q(n4789)
         );
  NAND2X0 U5062 ( .IN1(n4800), .IN2(n5135), .QN(n4788) );
  NAND2X0 U5063 ( .IN1(Datai[4]), .IN2(n4801), .QN(n4787) );
  NAND2X0 U5064 ( .IN1(\InstQueue[7][4] ), .IN2(n4802), .QN(n4786) );
  NAND4X0 U5065 ( .IN1(n4789), .IN2(n4788), .IN3(n4787), .IN4(n4786), .QN(
        n1804) );
  OA22X1 U5066 ( .IN1(n4808), .IN2(n5042), .IN3(n4799), .IN4(n5140), .Q(n4794)
         );
  NAND2X0 U5067 ( .IN1(n4790), .IN2(n5041), .QN(n4793) );
  NAND2X0 U5068 ( .IN1(Datai[5]), .IN2(n4801), .QN(n4792) );
  NAND2X0 U5069 ( .IN1(\InstQueue[7][5] ), .IN2(n4802), .QN(n4791) );
  NAND4X0 U5070 ( .IN1(n4794), .IN2(n4793), .IN3(n4792), .IN4(n4791), .QN(
        n1803) );
  OA22X1 U5071 ( .IN1(n4802), .IN2(n5148), .IN3(n5147), .IN4(n4799), .Q(n4798)
         );
  NAND2X0 U5072 ( .IN1(n4800), .IN2(n5149), .QN(n4797) );
  NAND2X0 U5073 ( .IN1(Datai[6]), .IN2(n4801), .QN(n4796) );
  NAND2X0 U5074 ( .IN1(\InstQueue[7][6] ), .IN2(n4802), .QN(n4795) );
  NAND4X0 U5075 ( .IN1(n4798), .IN2(n4797), .IN3(n4796), .IN4(n4795), .QN(
        n1802) );
  OA22X1 U5076 ( .IN1(n5156), .IN2(n4802), .IN3(n5155), .IN4(n4799), .Q(n4806)
         );
  NAND2X0 U5077 ( .IN1(n5158), .IN2(n4800), .QN(n4805) );
  NAND2X0 U5078 ( .IN1(Datai[7]), .IN2(n4801), .QN(n4804) );
  NAND2X0 U5079 ( .IN1(\InstQueue[7][7] ), .IN2(n4802), .QN(n4803) );
  NAND4X0 U5080 ( .IN1(n4806), .IN2(n4805), .IN3(n4804), .IN4(n4803), .QN(
        n1801) );
  NAND2X0 U5081 ( .IN1(n4807), .IN2(n4849), .QN(n4933) );
  OA22X1 U5082 ( .IN1(n4972), .IN2(n4933), .IN3(n4973), .IN4(n4893), .Q(n4809)
         );
  NOR2X0 U5083 ( .IN1(n5020), .IN2(n4852), .QN(n4841) );
  INVX0 U5084 ( .INP(n4841), .ZN(n4850) );
  NAND3X0 U5085 ( .IN1(n4809), .IN2(n4808), .IN3(n4850), .QN(n4831) );
  INVX0 U5086 ( .INP(n4831), .ZN(n4843) );
  OR2X1 U5087 ( .IN1(n4810), .IN2(n4843), .Q(n4840) );
  OA22X1 U5088 ( .IN1(n4843), .IN2(n5105), .IN3(n5100), .IN4(n4840), .Q(n4814)
         );
  AND4X1 U5089 ( .IN1(n4977), .IN2(n4852), .IN3(n4810), .IN4(n4831), .Q(n4842)
         );
  NAND2X0 U5090 ( .IN1(Datai[0]), .IN2(n4842), .QN(n4813) );
  NAND2X0 U5091 ( .IN1(\InstQueue[8][0] ), .IN2(n4843), .QN(n4812) );
  NAND2X0 U5092 ( .IN1(n4841), .IN2(n5108), .QN(n4811) );
  NAND4X0 U5093 ( .IN1(n4814), .IN2(n4813), .IN3(n4812), .IN4(n4811), .QN(
        n1800) );
  OA22X1 U5094 ( .IN1(n4843), .IN2(n5113), .IN3(n5112), .IN4(n4840), .Q(n4818)
         );
  NAND2X0 U5095 ( .IN1(Datai[1]), .IN2(n4842), .QN(n4817) );
  NAND2X0 U5096 ( .IN1(\InstQueue[8][1] ), .IN2(n4843), .QN(n4816) );
  NAND2X0 U5097 ( .IN1(n4841), .IN2(n5114), .QN(n4815) );
  NAND4X0 U5098 ( .IN1(n4818), .IN2(n4817), .IN3(n4816), .IN4(n4815), .QN(
        n1799) );
  OA22X1 U5099 ( .IN1(n4843), .IN2(n5120), .IN3(n5119), .IN4(n4840), .Q(n4822)
         );
  NAND2X0 U5100 ( .IN1(n4841), .IN2(n5121), .QN(n4821) );
  NAND2X0 U5101 ( .IN1(\InstQueue[8][2] ), .IN2(n4843), .QN(n4820) );
  NAND2X0 U5102 ( .IN1(Datai[2]), .IN2(n4842), .QN(n4819) );
  NAND4X0 U5103 ( .IN1(n4822), .IN2(n4821), .IN3(n4820), .IN4(n4819), .QN(
        n1798) );
  OA22X1 U5104 ( .IN1(n4843), .IN2(n5127), .IN3(n5126), .IN4(n4840), .Q(n4826)
         );
  NAND2X0 U5105 ( .IN1(n4841), .IN2(n5128), .QN(n4825) );
  NAND2X0 U5106 ( .IN1(\InstQueue[8][3] ), .IN2(n4843), .QN(n4824) );
  NAND2X0 U5107 ( .IN1(Datai[3]), .IN2(n4842), .QN(n4823) );
  NAND4X0 U5108 ( .IN1(n4826), .IN2(n4825), .IN3(n4824), .IN4(n4823), .QN(
        n1797) );
  OA22X1 U5109 ( .IN1(n4843), .IN2(n5134), .IN3(n5133), .IN4(n4840), .Q(n4830)
         );
  NAND2X0 U5110 ( .IN1(n4841), .IN2(n5135), .QN(n4829) );
  NAND2X0 U5111 ( .IN1(Datai[4]), .IN2(n4842), .QN(n4828) );
  NAND2X0 U5112 ( .IN1(\InstQueue[8][4] ), .IN2(n4843), .QN(n4827) );
  NAND4X0 U5113 ( .IN1(n4830), .IN2(n4829), .IN3(n4828), .IN4(n4827), .QN(
        n1796) );
  OA22X1 U5114 ( .IN1(n4850), .IN2(n5042), .IN3(n4840), .IN4(n5140), .Q(n4835)
         );
  NAND2X0 U5115 ( .IN1(n4831), .IN2(n5041), .QN(n4834) );
  NAND2X0 U5116 ( .IN1(Datai[5]), .IN2(n4842), .QN(n4833) );
  NAND2X0 U5117 ( .IN1(\InstQueue[8][5] ), .IN2(n4843), .QN(n4832) );
  NAND4X0 U5118 ( .IN1(n4835), .IN2(n4834), .IN3(n4833), .IN4(n4832), .QN(
        n1795) );
  OA22X1 U5119 ( .IN1(n4843), .IN2(n5148), .IN3(n5147), .IN4(n4840), .Q(n4839)
         );
  NAND2X0 U5120 ( .IN1(n4841), .IN2(n5149), .QN(n4838) );
  NAND2X0 U5121 ( .IN1(Datai[6]), .IN2(n4842), .QN(n4837) );
  NAND2X0 U5122 ( .IN1(\InstQueue[8][6] ), .IN2(n4843), .QN(n4836) );
  NAND4X0 U5123 ( .IN1(n4839), .IN2(n4838), .IN3(n4837), .IN4(n4836), .QN(
        n1794) );
  OA22X1 U5124 ( .IN1(n5156), .IN2(n4843), .IN3(n5155), .IN4(n4840), .Q(n4847)
         );
  NAND2X0 U5125 ( .IN1(n5158), .IN2(n4841), .QN(n4846) );
  NAND2X0 U5126 ( .IN1(Datai[7]), .IN2(n4842), .QN(n4845) );
  NAND2X0 U5127 ( .IN1(\InstQueue[8][7] ), .IN2(n4843), .QN(n4844) );
  NAND4X0 U5128 ( .IN1(n4847), .IN2(n4846), .IN3(n4845), .IN4(n4844), .QN(
        n1793) );
  NAND2X0 U5129 ( .IN1(n4849), .IN2(n4848), .QN(n4976) );
  OA22X1 U5130 ( .IN1(n4972), .IN2(n4976), .IN3(n4973), .IN4(n4933), .Q(n4851)
         );
  NOR2X0 U5131 ( .IN1(n5020), .IN2(n4893), .QN(n4883) );
  INVX0 U5132 ( .INP(n4883), .ZN(n4891) );
  NAND3X0 U5133 ( .IN1(n4851), .IN2(n4850), .IN3(n4891), .QN(n4873) );
  INVX0 U5134 ( .INP(n4873), .ZN(n4885) );
  OR2X1 U5135 ( .IN1(n4852), .IN2(n4885), .Q(n4882) );
  OA22X1 U5136 ( .IN1(n4885), .IN2(n5105), .IN3(n5100), .IN4(n4882), .Q(n4856)
         );
  AND4X1 U5137 ( .IN1(n4977), .IN2(n4893), .IN3(n4852), .IN4(n4873), .Q(n4884)
         );
  NAND2X0 U5138 ( .IN1(Datai[0]), .IN2(n4884), .QN(n4855) );
  NAND2X0 U5139 ( .IN1(\InstQueue[9][0] ), .IN2(n4885), .QN(n4854) );
  NAND2X0 U5140 ( .IN1(n4883), .IN2(n5108), .QN(n4853) );
  NAND4X0 U5141 ( .IN1(n4856), .IN2(n4855), .IN3(n4854), .IN4(n4853), .QN(
        n1792) );
  OA22X1 U5142 ( .IN1(n4885), .IN2(n5113), .IN3(n5112), .IN4(n4882), .Q(n4860)
         );
  NAND2X0 U5143 ( .IN1(Datai[1]), .IN2(n4884), .QN(n4859) );
  NAND2X0 U5144 ( .IN1(\InstQueue[9][1] ), .IN2(n4885), .QN(n4858) );
  NAND2X0 U5145 ( .IN1(n4883), .IN2(n5114), .QN(n4857) );
  NAND4X0 U5146 ( .IN1(n4860), .IN2(n4859), .IN3(n4858), .IN4(n4857), .QN(
        n1791) );
  OA22X1 U5147 ( .IN1(n4885), .IN2(n5120), .IN3(n5119), .IN4(n4882), .Q(n4864)
         );
  NAND2X0 U5148 ( .IN1(n4883), .IN2(n5121), .QN(n4863) );
  NAND2X0 U5149 ( .IN1(\InstQueue[9][2] ), .IN2(n4885), .QN(n4862) );
  NAND2X0 U5150 ( .IN1(Datai[2]), .IN2(n4884), .QN(n4861) );
  NAND4X0 U5151 ( .IN1(n4864), .IN2(n4863), .IN3(n4862), .IN4(n4861), .QN(
        n1790) );
  OA22X1 U5152 ( .IN1(n4885), .IN2(n5127), .IN3(n5126), .IN4(n4882), .Q(n4868)
         );
  NAND2X0 U5153 ( .IN1(n4883), .IN2(n5128), .QN(n4867) );
  NAND2X0 U5154 ( .IN1(\InstQueue[9][3] ), .IN2(n4885), .QN(n4866) );
  NAND2X0 U5155 ( .IN1(Datai[3]), .IN2(n4884), .QN(n4865) );
  NAND4X0 U5156 ( .IN1(n4868), .IN2(n4867), .IN3(n4866), .IN4(n4865), .QN(
        n1789) );
  OA22X1 U5157 ( .IN1(n4885), .IN2(n5134), .IN3(n5133), .IN4(n4882), .Q(n4872)
         );
  NAND2X0 U5158 ( .IN1(n4883), .IN2(n5135), .QN(n4871) );
  NAND2X0 U5159 ( .IN1(Datai[4]), .IN2(n4884), .QN(n4870) );
  NAND2X0 U5160 ( .IN1(\InstQueue[9][4] ), .IN2(n4885), .QN(n4869) );
  NAND4X0 U5161 ( .IN1(n4872), .IN2(n4871), .IN3(n4870), .IN4(n4869), .QN(
        n1788) );
  OA22X1 U5162 ( .IN1(n4891), .IN2(n5042), .IN3(n4882), .IN4(n5140), .Q(n4877)
         );
  NAND2X0 U5163 ( .IN1(n4873), .IN2(n5041), .QN(n4876) );
  NAND2X0 U5164 ( .IN1(Datai[5]), .IN2(n4884), .QN(n4875) );
  NAND2X0 U5165 ( .IN1(\InstQueue[9][5] ), .IN2(n4885), .QN(n4874) );
  NAND4X0 U5166 ( .IN1(n4877), .IN2(n4876), .IN3(n4875), .IN4(n4874), .QN(
        n1787) );
  OA22X1 U5167 ( .IN1(n4885), .IN2(n5148), .IN3(n5147), .IN4(n4882), .Q(n4881)
         );
  NAND2X0 U5168 ( .IN1(n4883), .IN2(n5149), .QN(n4880) );
  NAND2X0 U5169 ( .IN1(Datai[6]), .IN2(n4884), .QN(n4879) );
  NAND2X0 U5170 ( .IN1(\InstQueue[9][6] ), .IN2(n4885), .QN(n4878) );
  NAND4X0 U5171 ( .IN1(n4881), .IN2(n4880), .IN3(n4879), .IN4(n4878), .QN(
        n1786) );
  OA22X1 U5172 ( .IN1(n5156), .IN2(n4885), .IN3(n5155), .IN4(n4882), .Q(n4889)
         );
  NAND2X0 U5173 ( .IN1(n5158), .IN2(n4883), .QN(n4888) );
  NAND2X0 U5174 ( .IN1(Datai[7]), .IN2(n4884), .QN(n4887) );
  NAND2X0 U5175 ( .IN1(\InstQueue[9][7] ), .IN2(n4885), .QN(n4886) );
  NAND4X0 U5176 ( .IN1(n4889), .IN2(n4888), .IN3(n4887), .IN4(n4886), .QN(
        n1785) );
  NOR2X0 U5177 ( .IN1(n5182), .IN2(n4890), .QN(n5018) );
  NAND2X0 U5178 ( .IN1(n5018), .IN2(n5199), .QN(n5017) );
  OA22X1 U5179 ( .IN1(n4972), .IN2(n5017), .IN3(n4973), .IN4(n4976), .Q(n4892)
         );
  NOR2X0 U5180 ( .IN1(n5020), .IN2(n4933), .QN(n4924) );
  INVX0 U5181 ( .INP(n4924), .ZN(n4931) );
  NAND3X0 U5182 ( .IN1(n4892), .IN2(n4891), .IN3(n4931), .QN(n4914) );
  INVX0 U5183 ( .INP(n4914), .ZN(n4926) );
  OR2X1 U5184 ( .IN1(n4893), .IN2(n4926), .Q(n4923) );
  OA22X1 U5185 ( .IN1(n4926), .IN2(n5105), .IN3(n5100), .IN4(n4923), .Q(n4897)
         );
  AND4X1 U5186 ( .IN1(n4977), .IN2(n4933), .IN3(n4893), .IN4(n4914), .Q(n4925)
         );
  NAND2X0 U5187 ( .IN1(Datai[0]), .IN2(n4925), .QN(n4896) );
  NAND2X0 U5188 ( .IN1(\InstQueue[10][0] ), .IN2(n4926), .QN(n4895) );
  NAND2X0 U5189 ( .IN1(n4924), .IN2(n5108), .QN(n4894) );
  NAND4X0 U5190 ( .IN1(n4897), .IN2(n4896), .IN3(n4895), .IN4(n4894), .QN(
        n1784) );
  OA22X1 U5191 ( .IN1(n4926), .IN2(n5113), .IN3(n5112), .IN4(n4923), .Q(n4901)
         );
  NAND2X0 U5192 ( .IN1(Datai[1]), .IN2(n4925), .QN(n4900) );
  NAND2X0 U5193 ( .IN1(\InstQueue[10][1] ), .IN2(n4926), .QN(n4899) );
  NAND2X0 U5194 ( .IN1(n4924), .IN2(n5114), .QN(n4898) );
  NAND4X0 U5195 ( .IN1(n4901), .IN2(n4900), .IN3(n4899), .IN4(n4898), .QN(
        n1783) );
  OA22X1 U5196 ( .IN1(n4926), .IN2(n5120), .IN3(n5119), .IN4(n4923), .Q(n4905)
         );
  NAND2X0 U5197 ( .IN1(n4924), .IN2(n5121), .QN(n4904) );
  NAND2X0 U5198 ( .IN1(\InstQueue[10][2] ), .IN2(n4926), .QN(n4903) );
  NAND2X0 U5199 ( .IN1(Datai[2]), .IN2(n4925), .QN(n4902) );
  NAND4X0 U5200 ( .IN1(n4905), .IN2(n4904), .IN3(n4903), .IN4(n4902), .QN(
        n1782) );
  OA22X1 U5201 ( .IN1(n4926), .IN2(n5127), .IN3(n5126), .IN4(n4923), .Q(n4909)
         );
  NAND2X0 U5202 ( .IN1(n4924), .IN2(n5128), .QN(n4908) );
  NAND2X0 U5203 ( .IN1(\InstQueue[10][3] ), .IN2(n4926), .QN(n4907) );
  NAND2X0 U5204 ( .IN1(Datai[3]), .IN2(n4925), .QN(n4906) );
  NAND4X0 U5205 ( .IN1(n4909), .IN2(n4908), .IN3(n4907), .IN4(n4906), .QN(
        n1781) );
  OA22X1 U5206 ( .IN1(n4926), .IN2(n5134), .IN3(n5133), .IN4(n4923), .Q(n4913)
         );
  NAND2X0 U5207 ( .IN1(n4924), .IN2(n5135), .QN(n4912) );
  NAND2X0 U5208 ( .IN1(Datai[4]), .IN2(n4925), .QN(n4911) );
  NAND2X0 U5209 ( .IN1(\InstQueue[10][4] ), .IN2(n4926), .QN(n4910) );
  NAND4X0 U5210 ( .IN1(n4913), .IN2(n4912), .IN3(n4911), .IN4(n4910), .QN(
        n1780) );
  OA22X1 U5211 ( .IN1(n4931), .IN2(n5042), .IN3(n4923), .IN4(n5140), .Q(n4918)
         );
  NAND2X0 U5212 ( .IN1(n4914), .IN2(n5041), .QN(n4917) );
  NAND2X0 U5213 ( .IN1(Datai[5]), .IN2(n4925), .QN(n4916) );
  NAND2X0 U5214 ( .IN1(\InstQueue[10][5] ), .IN2(n4926), .QN(n4915) );
  NAND4X0 U5215 ( .IN1(n4918), .IN2(n4917), .IN3(n4916), .IN4(n4915), .QN(
        n1779) );
  OA22X1 U5216 ( .IN1(n4926), .IN2(n5148), .IN3(n5147), .IN4(n4923), .Q(n4922)
         );
  NAND2X0 U5217 ( .IN1(n4924), .IN2(n5149), .QN(n4921) );
  NAND2X0 U5218 ( .IN1(Datai[6]), .IN2(n4925), .QN(n4920) );
  NAND2X0 U5219 ( .IN1(\InstQueue[10][6] ), .IN2(n4926), .QN(n4919) );
  NAND4X0 U5220 ( .IN1(n4922), .IN2(n4921), .IN3(n4920), .IN4(n4919), .QN(
        n1778) );
  OA22X1 U5221 ( .IN1(n5156), .IN2(n4926), .IN3(n5155), .IN4(n4923), .Q(n4930)
         );
  NAND2X0 U5222 ( .IN1(n5158), .IN2(n4924), .QN(n4929) );
  NAND2X0 U5223 ( .IN1(Datai[7]), .IN2(n4925), .QN(n4928) );
  NAND2X0 U5224 ( .IN1(\InstQueue[10][7] ), .IN2(n4926), .QN(n4927) );
  NAND4X0 U5225 ( .IN1(n4930), .IN2(n4929), .IN3(n4928), .IN4(n4927), .QN(
        n1777) );
  OA22X1 U5226 ( .IN1(n4973), .IN2(n5017), .IN3(n4972), .IN4(n5019), .Q(n4932)
         );
  NOR2X0 U5227 ( .IN1(n5020), .IN2(n4976), .QN(n4964) );
  INVX0 U5228 ( .INP(n4964), .ZN(n4974) );
  NAND3X0 U5229 ( .IN1(n4932), .IN2(n4931), .IN3(n4974), .QN(n4954) );
  INVX0 U5230 ( .INP(n4954), .ZN(n4966) );
  OR2X1 U5231 ( .IN1(n4933), .IN2(n4966), .Q(n4963) );
  OA22X1 U5232 ( .IN1(n4966), .IN2(n5105), .IN3(n5100), .IN4(n4963), .Q(n4937)
         );
  AND4X1 U5233 ( .IN1(n4977), .IN2(n4976), .IN3(n4933), .IN4(n4954), .Q(n4965)
         );
  NAND2X0 U5234 ( .IN1(Datai[0]), .IN2(n4965), .QN(n4936) );
  NAND2X0 U5235 ( .IN1(\InstQueue[11][0] ), .IN2(n4966), .QN(n4935) );
  NAND2X0 U5236 ( .IN1(n4964), .IN2(n5108), .QN(n4934) );
  NAND4X0 U5237 ( .IN1(n4937), .IN2(n4936), .IN3(n4935), .IN4(n4934), .QN(
        n1776) );
  OA22X1 U5238 ( .IN1(n4966), .IN2(n5113), .IN3(n5112), .IN4(n4963), .Q(n4941)
         );
  NAND2X0 U5239 ( .IN1(Datai[1]), .IN2(n4965), .QN(n4940) );
  NAND2X0 U5240 ( .IN1(\InstQueue[11][1] ), .IN2(n4966), .QN(n4939) );
  NAND2X0 U5241 ( .IN1(n4964), .IN2(n5114), .QN(n4938) );
  NAND4X0 U5242 ( .IN1(n4941), .IN2(n4940), .IN3(n4939), .IN4(n4938), .QN(
        n1775) );
  OA22X1 U5243 ( .IN1(n4966), .IN2(n5120), .IN3(n5119), .IN4(n4963), .Q(n4945)
         );
  NAND2X0 U5244 ( .IN1(n4964), .IN2(n5121), .QN(n4944) );
  NAND2X0 U5245 ( .IN1(\InstQueue[11][2] ), .IN2(n4966), .QN(n4943) );
  NAND2X0 U5246 ( .IN1(Datai[2]), .IN2(n4965), .QN(n4942) );
  NAND4X0 U5247 ( .IN1(n4945), .IN2(n4944), .IN3(n4943), .IN4(n4942), .QN(
        n1774) );
  OA22X1 U5248 ( .IN1(n4966), .IN2(n5127), .IN3(n5126), .IN4(n4963), .Q(n4949)
         );
  NAND2X0 U5249 ( .IN1(n4964), .IN2(n5128), .QN(n4948) );
  NAND2X0 U5250 ( .IN1(\InstQueue[11][3] ), .IN2(n4966), .QN(n4947) );
  NAND2X0 U5251 ( .IN1(Datai[3]), .IN2(n4965), .QN(n4946) );
  NAND4X0 U5252 ( .IN1(n4949), .IN2(n4948), .IN3(n4947), .IN4(n4946), .QN(
        n1773) );
  OA22X1 U5253 ( .IN1(n4966), .IN2(n5134), .IN3(n5133), .IN4(n4963), .Q(n4953)
         );
  NAND2X0 U5254 ( .IN1(n4964), .IN2(n5135), .QN(n4952) );
  NAND2X0 U5255 ( .IN1(Datai[4]), .IN2(n4965), .QN(n4951) );
  NAND2X0 U5256 ( .IN1(\InstQueue[11][4] ), .IN2(n4966), .QN(n4950) );
  NAND4X0 U5257 ( .IN1(n4953), .IN2(n4952), .IN3(n4951), .IN4(n4950), .QN(
        n1772) );
  OA22X1 U5258 ( .IN1(n4974), .IN2(n5042), .IN3(n4963), .IN4(n5140), .Q(n4958)
         );
  NAND2X0 U5259 ( .IN1(n4954), .IN2(n5041), .QN(n4957) );
  NAND2X0 U5260 ( .IN1(Datai[5]), .IN2(n4965), .QN(n4956) );
  NAND2X0 U5261 ( .IN1(\InstQueue[11][5] ), .IN2(n4966), .QN(n4955) );
  NAND4X0 U5262 ( .IN1(n4958), .IN2(n4957), .IN3(n4956), .IN4(n4955), .QN(
        n1771) );
  OA22X1 U5263 ( .IN1(n4966), .IN2(n5148), .IN3(n5147), .IN4(n4963), .Q(n4962)
         );
  NAND2X0 U5264 ( .IN1(n4964), .IN2(n5149), .QN(n4961) );
  NAND2X0 U5265 ( .IN1(Datai[6]), .IN2(n4965), .QN(n4960) );
  NAND2X0 U5266 ( .IN1(\InstQueue[11][6] ), .IN2(n4966), .QN(n4959) );
  NAND4X0 U5267 ( .IN1(n4962), .IN2(n4961), .IN3(n4960), .IN4(n4959), .QN(
        n1770) );
  OA22X1 U5268 ( .IN1(n5156), .IN2(n4966), .IN3(n5155), .IN4(n4963), .Q(n4970)
         );
  NAND2X0 U5269 ( .IN1(n5158), .IN2(n4964), .QN(n4969) );
  NAND2X0 U5270 ( .IN1(Datai[7]), .IN2(n4965), .QN(n4968) );
  NAND2X0 U5271 ( .IN1(\InstQueue[11][7] ), .IN2(n4966), .QN(n4967) );
  NAND4X0 U5272 ( .IN1(n4970), .IN2(n4969), .IN3(n4968), .IN4(n4967), .QN(
        n1769) );
  OA22X1 U5273 ( .IN1(n4973), .IN2(n5019), .IN3(n4972), .IN4(n4971), .Q(n4975)
         );
  NOR2X0 U5274 ( .IN1(n5020), .IN2(n5017), .QN(n5009) );
  INVX0 U5275 ( .INP(n5009), .ZN(n4998) );
  NAND3X0 U5276 ( .IN1(n4975), .IN2(n4974), .IN3(n4998), .QN(n4999) );
  INVX0 U5277 ( .INP(n4999), .ZN(n5011) );
  OR2X1 U5278 ( .IN1(n4976), .IN2(n5011), .Q(n5008) );
  OA22X1 U5279 ( .IN1(n5011), .IN2(n5105), .IN3(n5100), .IN4(n5008), .Q(n4981)
         );
  AND4X1 U5280 ( .IN1(n4977), .IN2(n5017), .IN3(n4976), .IN4(n4999), .Q(n5010)
         );
  NAND2X0 U5281 ( .IN1(Datai[0]), .IN2(n5010), .QN(n4980) );
  NAND2X0 U5282 ( .IN1(\InstQueue[12][0] ), .IN2(n5011), .QN(n4979) );
  NAND2X0 U5283 ( .IN1(n5009), .IN2(n5108), .QN(n4978) );
  NAND4X0 U5284 ( .IN1(n4981), .IN2(n4980), .IN3(n4979), .IN4(n4978), .QN(
        n1768) );
  OA22X1 U5285 ( .IN1(n5011), .IN2(n5113), .IN3(n5112), .IN4(n5008), .Q(n4985)
         );
  NAND2X0 U5286 ( .IN1(Datai[1]), .IN2(n5010), .QN(n4984) );
  NAND2X0 U5287 ( .IN1(\InstQueue[12][1] ), .IN2(n5011), .QN(n4983) );
  NAND2X0 U5288 ( .IN1(n5009), .IN2(n5114), .QN(n4982) );
  NAND4X0 U5289 ( .IN1(n4985), .IN2(n4984), .IN3(n4983), .IN4(n4982), .QN(
        n1767) );
  OA22X1 U5290 ( .IN1(n5011), .IN2(n5120), .IN3(n5119), .IN4(n5008), .Q(n4989)
         );
  NAND2X0 U5291 ( .IN1(n5009), .IN2(n5121), .QN(n4988) );
  NAND2X0 U5292 ( .IN1(\InstQueue[12][2] ), .IN2(n5011), .QN(n4987) );
  NAND2X0 U5293 ( .IN1(Datai[2]), .IN2(n5010), .QN(n4986) );
  NAND4X0 U5294 ( .IN1(n4989), .IN2(n4988), .IN3(n4987), .IN4(n4986), .QN(
        n1766) );
  OA22X1 U5295 ( .IN1(n5011), .IN2(n5127), .IN3(n5126), .IN4(n5008), .Q(n4993)
         );
  NAND2X0 U5296 ( .IN1(n5009), .IN2(n5128), .QN(n4992) );
  NAND2X0 U5297 ( .IN1(\InstQueue[12][3] ), .IN2(n5011), .QN(n4991) );
  NAND2X0 U5298 ( .IN1(Datai[3]), .IN2(n5010), .QN(n4990) );
  NAND4X0 U5299 ( .IN1(n4993), .IN2(n4992), .IN3(n4991), .IN4(n4990), .QN(
        n1765) );
  OA22X1 U5300 ( .IN1(n5011), .IN2(n5134), .IN3(n5133), .IN4(n5008), .Q(n4997)
         );
  NAND2X0 U5301 ( .IN1(n5009), .IN2(n5135), .QN(n4996) );
  NAND2X0 U5302 ( .IN1(Datai[4]), .IN2(n5010), .QN(n4995) );
  NAND2X0 U5303 ( .IN1(\InstQueue[12][4] ), .IN2(n5011), .QN(n4994) );
  NAND4X0 U5304 ( .IN1(n4997), .IN2(n4996), .IN3(n4995), .IN4(n4994), .QN(
        n1764) );
  OA22X1 U5305 ( .IN1(n4998), .IN2(n5042), .IN3(n5008), .IN4(n5140), .Q(n5003)
         );
  NAND2X0 U5306 ( .IN1(n4999), .IN2(n5041), .QN(n5002) );
  NAND2X0 U5307 ( .IN1(Datai[5]), .IN2(n5010), .QN(n5001) );
  NAND2X0 U5308 ( .IN1(\InstQueue[12][5] ), .IN2(n5011), .QN(n5000) );
  NAND4X0 U5309 ( .IN1(n5003), .IN2(n5002), .IN3(n5001), .IN4(n5000), .QN(
        n1763) );
  OA22X1 U5310 ( .IN1(n5011), .IN2(n5148), .IN3(n5147), .IN4(n5008), .Q(n5007)
         );
  NAND2X0 U5311 ( .IN1(n5009), .IN2(n5149), .QN(n5006) );
  NAND2X0 U5312 ( .IN1(Datai[6]), .IN2(n5010), .QN(n5005) );
  NAND2X0 U5313 ( .IN1(\InstQueue[12][6] ), .IN2(n5011), .QN(n5004) );
  NAND4X0 U5314 ( .IN1(n5007), .IN2(n5006), .IN3(n5005), .IN4(n5004), .QN(
        n1762) );
  OA22X1 U5315 ( .IN1(n5156), .IN2(n5011), .IN3(n5155), .IN4(n5008), .Q(n5015)
         );
  NAND2X0 U5316 ( .IN1(n5158), .IN2(n5009), .QN(n5014) );
  NAND2X0 U5317 ( .IN1(Datai[7]), .IN2(n5010), .QN(n5013) );
  NAND2X0 U5318 ( .IN1(\InstQueue[12][7] ), .IN2(n5011), .QN(n5012) );
  NAND4X0 U5319 ( .IN1(n5015), .IN2(n5014), .IN3(n5013), .IN4(n5012), .QN(
        n1761) );
  AOI222X1 U5320 ( .IN1(n5096), .IN2(n5102), .IN3(n5106), .IN4(n5016), .IN5(
        n5098), .IN6(n5018), .QN(n5054) );
  OR2X1 U5321 ( .IN1(n5017), .IN2(n5054), .Q(n5051) );
  OA22X1 U5322 ( .IN1(n5054), .IN2(n5105), .IN3(n5100), .IN4(n5051), .Q(n5024)
         );
  NOR3X0 U5323 ( .IN1(n5018), .IN2(n5054), .IN3(n5101), .QN(n5053) );
  NAND2X0 U5324 ( .IN1(Datai[0]), .IN2(n5053), .QN(n5023) );
  NAND2X0 U5325 ( .IN1(\InstQueue[13][0] ), .IN2(n5054), .QN(n5022) );
  NOR2X0 U5326 ( .IN1(n5020), .IN2(n5019), .QN(n5052) );
  NAND2X0 U5327 ( .IN1(n5052), .IN2(n5108), .QN(n5021) );
  NAND4X0 U5328 ( .IN1(n5024), .IN2(n5023), .IN3(n5022), .IN4(n5021), .QN(
        n1760) );
  OA22X1 U5329 ( .IN1(n5054), .IN2(n5113), .IN3(n5112), .IN4(n5051), .Q(n5028)
         );
  NAND2X0 U5330 ( .IN1(n5052), .IN2(n5114), .QN(n5027) );
  NAND2X0 U5331 ( .IN1(\InstQueue[13][1] ), .IN2(n5054), .QN(n5026) );
  NAND2X0 U5332 ( .IN1(Datai[1]), .IN2(n5053), .QN(n5025) );
  NAND4X0 U5333 ( .IN1(n5028), .IN2(n5027), .IN3(n5026), .IN4(n5025), .QN(
        n1759) );
  OA22X1 U5334 ( .IN1(n5054), .IN2(n5120), .IN3(n5119), .IN4(n5051), .Q(n5032)
         );
  NAND2X0 U5335 ( .IN1(n5052), .IN2(n5121), .QN(n5031) );
  NAND2X0 U5336 ( .IN1(\InstQueue[13][2] ), .IN2(n5054), .QN(n5030) );
  NAND2X0 U5337 ( .IN1(Datai[2]), .IN2(n5053), .QN(n5029) );
  NAND4X0 U5338 ( .IN1(n5032), .IN2(n5031), .IN3(n5030), .IN4(n5029), .QN(
        n1758) );
  OA22X1 U5339 ( .IN1(n5054), .IN2(n5127), .IN3(n5126), .IN4(n5051), .Q(n5036)
         );
  NAND2X0 U5340 ( .IN1(n5052), .IN2(n5128), .QN(n5035) );
  NAND2X0 U5341 ( .IN1(\InstQueue[13][3] ), .IN2(n5054), .QN(n5034) );
  NAND2X0 U5342 ( .IN1(Datai[3]), .IN2(n5053), .QN(n5033) );
  NAND4X0 U5343 ( .IN1(n5036), .IN2(n5035), .IN3(n5034), .IN4(n5033), .QN(
        n1757) );
  OA22X1 U5344 ( .IN1(n5054), .IN2(n5134), .IN3(n5133), .IN4(n5051), .Q(n5040)
         );
  NAND2X0 U5345 ( .IN1(n5052), .IN2(n5135), .QN(n5039) );
  NAND2X0 U5346 ( .IN1(Datai[4]), .IN2(n5053), .QN(n5038) );
  NAND2X0 U5347 ( .IN1(\InstQueue[13][4] ), .IN2(n5054), .QN(n5037) );
  NAND4X0 U5348 ( .IN1(n5040), .IN2(n5039), .IN3(n5038), .IN4(n5037), .QN(
        n1756) );
  INVX0 U5349 ( .INP(n5041), .ZN(n5141) );
  OA22X1 U5350 ( .IN1(n5054), .IN2(n5141), .IN3(n5140), .IN4(n5051), .Q(n5046)
         );
  INVX0 U5351 ( .INP(n5042), .ZN(n5142) );
  NAND2X0 U5352 ( .IN1(n5052), .IN2(n5142), .QN(n5045) );
  NAND2X0 U5353 ( .IN1(Datai[5]), .IN2(n5053), .QN(n5044) );
  NAND2X0 U5354 ( .IN1(\InstQueue[13][5] ), .IN2(n5054), .QN(n5043) );
  NAND4X0 U5355 ( .IN1(n5046), .IN2(n5045), .IN3(n5044), .IN4(n5043), .QN(
        n1755) );
  OA22X1 U5356 ( .IN1(n5054), .IN2(n5148), .IN3(n5147), .IN4(n5051), .Q(n5050)
         );
  NAND2X0 U5357 ( .IN1(n5052), .IN2(n5149), .QN(n5049) );
  NAND2X0 U5358 ( .IN1(Datai[6]), .IN2(n5053), .QN(n5048) );
  NAND2X0 U5359 ( .IN1(\InstQueue[13][6] ), .IN2(n5054), .QN(n5047) );
  NAND4X0 U5360 ( .IN1(n5050), .IN2(n5049), .IN3(n5048), .IN4(n5047), .QN(
        n1754) );
  OA22X1 U5361 ( .IN1(n5156), .IN2(n5054), .IN3(n5155), .IN4(n5051), .Q(n5058)
         );
  NAND2X0 U5362 ( .IN1(n5158), .IN2(n5052), .QN(n5057) );
  NAND2X0 U5363 ( .IN1(Datai[7]), .IN2(n5053), .QN(n5056) );
  NAND2X0 U5364 ( .IN1(\InstQueue[13][7] ), .IN2(n5054), .QN(n5055) );
  NAND4X0 U5365 ( .IN1(n5058), .IN2(n5057), .IN3(n5056), .IN4(n5055), .QN(
        n1753) );
  NAND2X0 U5366 ( .IN1(n5088), .IN2(Datai[0]), .QN(n5062) );
  INVX0 U5367 ( .INP(n5108), .ZN(n5059) );
  INVX0 U5368 ( .INP(n5087), .ZN(n5064) );
  OA22X1 U5369 ( .IN1(n5089), .IN2(n5105), .IN3(n5059), .IN4(n5064), .Q(n5061)
         );
  OA22X1 U5370 ( .IN1(n5249), .IN2(n5069), .IN3(n5086), .IN4(n5100), .Q(n5060)
         );
  NAND3X0 U5371 ( .IN1(n5062), .IN2(n5061), .IN3(n5060), .QN(n1752) );
  NAND2X0 U5372 ( .IN1(n5088), .IN2(Datai[1]), .QN(n5066) );
  OA22X1 U5373 ( .IN1(n5064), .IN2(n5063), .IN3(n5086), .IN4(n5112), .Q(n5065)
         );
  NAND2X0 U5374 ( .IN1(n5066), .IN2(n5065), .QN(n5067) );
  AO221X1 U5375 ( .IN1(n5089), .IN2(\InstQueue[14][1] ), .IN3(n5069), .IN4(
        n5068), .IN5(n5067), .Q(n1751) );
  OA22X1 U5376 ( .IN1(n5089), .IN2(n5120), .IN3(n5119), .IN4(n5086), .Q(n5073)
         );
  NAND2X0 U5377 ( .IN1(Datai[2]), .IN2(n5088), .QN(n5072) );
  NAND2X0 U5378 ( .IN1(n5087), .IN2(n5121), .QN(n5071) );
  NAND2X0 U5379 ( .IN1(\InstQueue[14][2] ), .IN2(n5089), .QN(n5070) );
  NAND4X0 U5380 ( .IN1(n5073), .IN2(n5072), .IN3(n5071), .IN4(n5070), .QN(
        n1750) );
  OA22X1 U5381 ( .IN1(n5089), .IN2(n5127), .IN3(n5126), .IN4(n5086), .Q(n5077)
         );
  NAND2X0 U5382 ( .IN1(n5087), .IN2(n5128), .QN(n5076) );
  NAND2X0 U5383 ( .IN1(Datai[3]), .IN2(n5088), .QN(n5075) );
  NAND2X0 U5384 ( .IN1(\InstQueue[14][3] ), .IN2(n5089), .QN(n5074) );
  NAND4X0 U5385 ( .IN1(n5077), .IN2(n5076), .IN3(n5075), .IN4(n5074), .QN(
        n1749) );
  OA22X1 U5386 ( .IN1(n5089), .IN2(n5134), .IN3(n5133), .IN4(n5086), .Q(n5081)
         );
  NAND2X0 U5387 ( .IN1(n5087), .IN2(n5135), .QN(n5080) );
  NAND2X0 U5388 ( .IN1(Datai[4]), .IN2(n5088), .QN(n5079) );
  NAND2X0 U5389 ( .IN1(\InstQueue[14][4] ), .IN2(n5089), .QN(n5078) );
  NAND4X0 U5390 ( .IN1(n5081), .IN2(n5080), .IN3(n5079), .IN4(n5078), .QN(
        n1748) );
  OA22X1 U5391 ( .IN1(n5089), .IN2(n5141), .IN3(n5140), .IN4(n5086), .Q(n5085)
         );
  NAND2X0 U5392 ( .IN1(n5087), .IN2(n5142), .QN(n5084) );
  NAND2X0 U5393 ( .IN1(Datai[5]), .IN2(n5088), .QN(n5083) );
  NAND2X0 U5394 ( .IN1(\InstQueue[14][5] ), .IN2(n5089), .QN(n5082) );
  NAND4X0 U5395 ( .IN1(n5085), .IN2(n5084), .IN3(n5083), .IN4(n5082), .QN(
        n1747) );
  OA22X1 U5396 ( .IN1(n5089), .IN2(n5148), .IN3(n5147), .IN4(n5086), .Q(n5093)
         );
  NAND2X0 U5397 ( .IN1(n5087), .IN2(n5149), .QN(n5092) );
  NAND2X0 U5398 ( .IN1(Datai[6]), .IN2(n5088), .QN(n5091) );
  NAND2X0 U5399 ( .IN1(\InstQueue[14][6] ), .IN2(n5089), .QN(n5090) );
  NAND4X0 U5400 ( .IN1(n5093), .IN2(n5092), .IN3(n5091), .IN4(n5090), .QN(
        n1746) );
  AO222X1 U5401 ( .IN1(n5098), .IN2(n5102), .IN3(n5097), .IN4(n5096), .IN5(
        n5095), .IN6(n5094), .Q(n5107) );
  NAND2X0 U5402 ( .IN1(n5099), .IN2(n5107), .QN(n5154) );
  OA22X1 U5403 ( .IN1(n5252), .IN2(n5107), .IN3(n5154), .IN4(n5100), .Q(n5111)
         );
  INVX0 U5404 ( .INP(n5107), .ZN(n5160) );
  NOR3X0 U5405 ( .IN1(n5102), .IN2(n5160), .IN3(n5101), .QN(n5159) );
  INVX0 U5406 ( .INP(n5159), .ZN(n5103) );
  OA22X1 U5407 ( .IN1(n5160), .IN2(n5105), .IN3(n5104), .IN4(n5103), .Q(n5110)
         );
  AND2X1 U5408 ( .IN1(n5107), .IN2(n5106), .Q(n5157) );
  NAND2X0 U5409 ( .IN1(n5157), .IN2(n5108), .QN(n5109) );
  NAND3X0 U5410 ( .IN1(n5111), .IN2(n5110), .IN3(n5109), .QN(n1744) );
  OA22X1 U5411 ( .IN1(n5160), .IN2(n5113), .IN3(n5112), .IN4(n5154), .Q(n5118)
         );
  NAND2X0 U5412 ( .IN1(Datai[1]), .IN2(n5159), .QN(n5117) );
  NAND2X0 U5413 ( .IN1(\InstQueue[15][1] ), .IN2(n5160), .QN(n5116) );
  NAND2X0 U5414 ( .IN1(n5157), .IN2(n5114), .QN(n5115) );
  NAND4X0 U5415 ( .IN1(n5118), .IN2(n5117), .IN3(n5116), .IN4(n5115), .QN(
        n1743) );
  OA22X1 U5416 ( .IN1(n5160), .IN2(n5120), .IN3(n5119), .IN4(n5154), .Q(n5125)
         );
  NAND2X0 U5417 ( .IN1(n5157), .IN2(n5121), .QN(n5124) );
  NAND2X0 U5418 ( .IN1(\InstQueue[15][2] ), .IN2(n5160), .QN(n5123) );
  NAND2X0 U5419 ( .IN1(Datai[2]), .IN2(n5159), .QN(n5122) );
  NAND4X0 U5420 ( .IN1(n5125), .IN2(n5124), .IN3(n5123), .IN4(n5122), .QN(
        n1742) );
  OA22X1 U5421 ( .IN1(n5160), .IN2(n5127), .IN3(n5126), .IN4(n5154), .Q(n5132)
         );
  NAND2X0 U5422 ( .IN1(n5157), .IN2(n5128), .QN(n5131) );
  NAND2X0 U5423 ( .IN1(\InstQueue[15][3] ), .IN2(n5160), .QN(n5130) );
  NAND2X0 U5424 ( .IN1(Datai[3]), .IN2(n5159), .QN(n5129) );
  NAND4X0 U5425 ( .IN1(n5132), .IN2(n5131), .IN3(n5130), .IN4(n5129), .QN(
        n1741) );
  OA22X1 U5426 ( .IN1(n5160), .IN2(n5134), .IN3(n5133), .IN4(n5154), .Q(n5139)
         );
  NAND2X0 U5427 ( .IN1(n5157), .IN2(n5135), .QN(n5138) );
  NAND2X0 U5428 ( .IN1(\InstQueue[15][4] ), .IN2(n5160), .QN(n5137) );
  NAND2X0 U5429 ( .IN1(Datai[4]), .IN2(n5159), .QN(n5136) );
  NAND4X0 U5430 ( .IN1(n5139), .IN2(n5138), .IN3(n5137), .IN4(n5136), .QN(
        n1740) );
  OA22X1 U5431 ( .IN1(n5160), .IN2(n5141), .IN3(n5140), .IN4(n5154), .Q(n5146)
         );
  NAND2X0 U5432 ( .IN1(n5157), .IN2(n5142), .QN(n5145) );
  NAND2X0 U5433 ( .IN1(Datai[5]), .IN2(n5159), .QN(n5144) );
  NAND2X0 U5434 ( .IN1(\InstQueue[15][5] ), .IN2(n5160), .QN(n5143) );
  NAND4X0 U5435 ( .IN1(n5146), .IN2(n5145), .IN3(n5144), .IN4(n5143), .QN(
        n1739) );
  OA22X1 U5436 ( .IN1(n5160), .IN2(n5148), .IN3(n5147), .IN4(n5154), .Q(n5153)
         );
  NAND2X0 U5437 ( .IN1(n5157), .IN2(n5149), .QN(n5152) );
  NAND2X0 U5438 ( .IN1(Datai[6]), .IN2(n5159), .QN(n5151) );
  NAND2X0 U5439 ( .IN1(\InstQueue[15][6] ), .IN2(n5160), .QN(n5150) );
  NAND4X0 U5440 ( .IN1(n5153), .IN2(n5152), .IN3(n5151), .IN4(n5150), .QN(
        n1738) );
  OA22X1 U5441 ( .IN1(n5156), .IN2(n5160), .IN3(n5155), .IN4(n5154), .Q(n5164)
         );
  NAND2X0 U5442 ( .IN1(n5158), .IN2(n5157), .QN(n5163) );
  NAND2X0 U5443 ( .IN1(Datai[7]), .IN2(n5159), .QN(n5162) );
  NAND2X0 U5444 ( .IN1(\InstQueue[15][7] ), .IN2(n5160), .QN(n5161) );
  NAND4X0 U5445 ( .IN1(n5164), .IN2(n5163), .IN3(n5162), .IN4(n5161), .QN(
        n1737) );
  OAI22X1 U5446 ( .IN1(BS16_n), .IN2(n5166), .IN3(n5169), .IN4(n5250), .QN(
        n1704) );
  AO21X1 U5447 ( .IN1(DataWidth[1]), .IN2(n5166), .IN3(n5165), .Q(n1703) );
  INVX0 U5448 ( .INP(n5168), .ZN(n5170) );
  MUX21X1 U5449 ( .IN1(MemoryFetch), .IN2(M_IO_n), .S(n5170), .Q(n1672) );
  MUX21X1 U5450 ( .IN1(n5251), .IN2(W_R_n), .S(n5170), .Q(n1671) );
  AO221X1 U5451 ( .IN1(n5168), .IN2(n5197), .IN3(n5170), .IN4(D_C_n), .IN5(
        n5167), .Q(n1670) );
  AO21X1 U5452 ( .IN1(State[0]), .IN2(ADS_n), .IN3(n5169), .Q(n1669) );
  MUX21X1 U5453 ( .IN1(ByteEnable[3]), .IN2(BE_n[3]), .S(n5170), .Q(n1668) );
  MUX21X1 U5454 ( .IN1(ByteEnable[2]), .IN2(BE_n[2]), .S(n5170), .Q(n1667) );
  MUX21X1 U5455 ( .IN1(ByteEnable[1]), .IN2(BE_n[1]), .S(n5170), .Q(n1666) );
  MUX21X1 U5456 ( .IN1(ByteEnable[0]), .IN2(BE_n[0]), .S(n5170), .Q(n1664) );
  NAND2X0 U5457 ( .IN1(rEIP[0]), .IN2(DataWidth[0]), .QN(n5172) );
  AO222X1 U5458 ( .IN1(n5172), .IN2(n5171), .IN3(n5175), .IN4(ByteEnable[2]), 
        .IN5(rEIP[0]), .IN6(n5173), .Q(n1662) );
  AO221X1 U5459 ( .IN1(n5175), .IN2(ByteEnable[0]), .IN3(n5174), .IN4(rEIP[0]), 
        .IN5(n5173), .Q(n1660) );
endmodule

