
module wb_conmax_top ( clock, rst_i, m0_data_i, m0_data_o, m0_addr_i, m0_sel_i, 
        m0_we_i, m0_cyc_i, m0_stb_i, m0_ack_o, m0_err_o, m0_rty_o, m1_data_i, 
        m1_data_o, m1_addr_i, m1_sel_i, m1_we_i, m1_cyc_i, m1_stb_i, m1_ack_o, 
        m1_err_o, m1_rty_o, m2_data_i, m2_data_o, m2_addr_i, m2_sel_i, m2_we_i, 
        m2_cyc_i, m2_stb_i, m2_ack_o, m2_err_o, m2_rty_o, m3_data_i, m3_data_o, 
        m3_addr_i, m3_sel_i, m3_we_i, m3_cyc_i, m3_stb_i, m3_ack_o, m3_err_o, 
        m3_rty_o, m4_data_i, m4_data_o, m4_addr_i, m4_sel_i, m4_we_i, m4_cyc_i, 
        m4_stb_i, m4_ack_o, m4_err_o, m4_rty_o, m5_data_i, m5_data_o, 
        m5_addr_i, m5_sel_i, m5_we_i, m5_cyc_i, m5_stb_i, m5_ack_o, m5_err_o, 
        m5_rty_o, m6_data_i, m6_data_o, m6_addr_i, m6_sel_i, m6_we_i, m6_cyc_i, 
        m6_stb_i, m6_ack_o, m6_err_o, m6_rty_o, m7_data_i, m7_data_o, 
        m7_addr_i, m7_sel_i, m7_we_i, m7_cyc_i, m7_stb_i, m7_ack_o, m7_err_o, 
        m7_rty_o, s0_data_i, s0_data_o, s0_addr_o, s0_sel_o, s0_we_o, s0_cyc_o, 
        s0_stb_o, s0_ack_i, s0_err_i, s0_rty_i, s1_data_i, s1_data_o, 
        s1_addr_o, s1_sel_o, s1_we_o, s1_cyc_o, s1_stb_o, s1_ack_i, s1_err_i, 
        s1_rty_i, s2_data_i, s2_data_o, s2_addr_o, s2_sel_o, s2_we_o, s2_cyc_o, 
        s2_stb_o, s2_ack_i, s2_err_i, s2_rty_i, s3_data_i, s3_data_o, 
        s3_addr_o, s3_sel_o, s3_we_o, s3_cyc_o, s3_stb_o, s3_ack_i, s3_err_i, 
        s3_rty_i, s4_data_i, s4_data_o, s4_addr_o, s4_sel_o, s4_we_o, s4_cyc_o, 
        s4_stb_o, s4_ack_i, s4_err_i, s4_rty_i, s5_data_i, s5_data_o, 
        s5_addr_o, s5_sel_o, s5_we_o, s5_cyc_o, s5_stb_o, s5_ack_i, s5_err_i, 
        s5_rty_i, s6_data_i, s6_data_o, s6_addr_o, s6_sel_o, s6_we_o, s6_cyc_o, 
        s6_stb_o, s6_ack_i, s6_err_i, s6_rty_i, s7_data_i, s7_data_o, 
        s7_addr_o, s7_sel_o, s7_we_o, s7_cyc_o, s7_stb_o, s7_ack_i, s7_err_i, 
        s7_rty_i, s8_data_i, s8_data_o, s8_addr_o, s8_sel_o, s8_we_o, s8_cyc_o, 
        s8_stb_o, s8_ack_i, s8_err_i, s8_rty_i, s9_data_i, s9_data_o, 
        s9_addr_o, s9_sel_o, s9_we_o, s9_cyc_o, s9_stb_o, s9_ack_i, s9_err_i, 
        s9_rty_i, s10_data_i, s10_data_o, s10_addr_o, s10_sel_o, s10_we_o, 
        s10_cyc_o, s10_stb_o, s10_ack_i, s10_err_i, s10_rty_i, s11_data_i, 
        s11_data_o, s11_addr_o, s11_sel_o, s11_we_o, s11_cyc_o, s11_stb_o, 
        s11_ack_i, s11_err_i, s11_rty_i, s12_data_i, s12_data_o, s12_addr_o, 
        s12_sel_o, s12_we_o, s12_cyc_o, s12_stb_o, s12_ack_i, s12_err_i, 
        s12_rty_i, s13_data_i, s13_data_o, s13_addr_o, s13_sel_o, s13_we_o, 
        s13_cyc_o, s13_stb_o, s13_ack_i, s13_err_i, s13_rty_i, s14_data_i, 
        s14_data_o, s14_addr_o, s14_sel_o, s14_we_o, s14_cyc_o, s14_stb_o, 
        s14_ack_i, s14_err_i, s14_rty_i, s15_data_i, s15_data_o, s15_addr_o, 
        s15_sel_o, s15_we_o, s15_cyc_o, s15_stb_o, s15_ack_i, s15_err_i, 
        s15_rty_i );
  input [31:0] m0_data_i;
  output [31:0] m0_data_o;
  input [31:0] m0_addr_i;
  input [3:0] m0_sel_i;
  input [31:0] m1_data_i;
  output [31:0] m1_data_o;
  input [31:0] m1_addr_i;
  input [3:0] m1_sel_i;
  input [31:0] m2_data_i;
  output [31:0] m2_data_o;
  input [31:0] m2_addr_i;
  input [3:0] m2_sel_i;
  input [31:0] m3_data_i;
  output [31:0] m3_data_o;
  input [31:0] m3_addr_i;
  input [3:0] m3_sel_i;
  input [31:0] m4_data_i;
  output [31:0] m4_data_o;
  input [31:0] m4_addr_i;
  input [3:0] m4_sel_i;
  input [31:0] m5_data_i;
  output [31:0] m5_data_o;
  input [31:0] m5_addr_i;
  input [3:0] m5_sel_i;
  input [31:0] m6_data_i;
  output [31:0] m6_data_o;
  input [31:0] m6_addr_i;
  input [3:0] m6_sel_i;
  input [31:0] m7_data_i;
  output [31:0] m7_data_o;
  input [31:0] m7_addr_i;
  input [3:0] m7_sel_i;
  input [31:0] s0_data_i;
  output [31:0] s0_data_o;
  output [31:0] s0_addr_o;
  output [3:0] s0_sel_o;
  input [31:0] s1_data_i;
  output [31:0] s1_data_o;
  output [31:0] s1_addr_o;
  output [3:0] s1_sel_o;
  input [31:0] s2_data_i;
  output [31:0] s2_data_o;
  output [31:0] s2_addr_o;
  output [3:0] s2_sel_o;
  input [31:0] s3_data_i;
  output [31:0] s3_data_o;
  output [31:0] s3_addr_o;
  output [3:0] s3_sel_o;
  input [31:0] s4_data_i;
  output [31:0] s4_data_o;
  output [31:0] s4_addr_o;
  output [3:0] s4_sel_o;
  input [31:0] s5_data_i;
  output [31:0] s5_data_o;
  output [31:0] s5_addr_o;
  output [3:0] s5_sel_o;
  input [31:0] s6_data_i;
  output [31:0] s6_data_o;
  output [31:0] s6_addr_o;
  output [3:0] s6_sel_o;
  input [31:0] s7_data_i;
  output [31:0] s7_data_o;
  output [31:0] s7_addr_o;
  output [3:0] s7_sel_o;
  input [31:0] s8_data_i;
  output [31:0] s8_data_o;
  output [31:0] s8_addr_o;
  output [3:0] s8_sel_o;
  input [31:0] s9_data_i;
  output [31:0] s9_data_o;
  output [31:0] s9_addr_o;
  output [3:0] s9_sel_o;
  input [31:0] s10_data_i;
  output [31:0] s10_data_o;
  output [31:0] s10_addr_o;
  output [3:0] s10_sel_o;
  input [31:0] s11_data_i;
  output [31:0] s11_data_o;
  output [31:0] s11_addr_o;
  output [3:0] s11_sel_o;
  input [31:0] s12_data_i;
  output [31:0] s12_data_o;
  output [31:0] s12_addr_o;
  output [3:0] s12_sel_o;
  input [31:0] s13_data_i;
  output [31:0] s13_data_o;
  output [31:0] s13_addr_o;
  output [3:0] s13_sel_o;
  input [31:0] s14_data_i;
  output [31:0] s14_data_o;
  output [31:0] s14_addr_o;
  output [3:0] s14_sel_o;
  input [31:0] s15_data_i;
  output [31:0] s15_data_o;
  output [31:0] s15_addr_o;
  output [3:0] s15_sel_o;
  input clock, rst_i, m0_we_i, m0_cyc_i, m0_stb_i, m1_we_i, m1_cyc_i, m1_stb_i,
         m2_we_i, m2_cyc_i, m2_stb_i, m3_we_i, m3_cyc_i, m3_stb_i, m4_we_i,
         m4_cyc_i, m4_stb_i, m5_we_i, m5_cyc_i, m5_stb_i, m6_we_i, m6_cyc_i,
         m6_stb_i, m7_we_i, m7_cyc_i, m7_stb_i, s0_ack_i, s0_err_i, s0_rty_i,
         s1_ack_i, s1_err_i, s1_rty_i, s2_ack_i, s2_err_i, s2_rty_i, s3_ack_i,
         s3_err_i, s3_rty_i, s4_ack_i, s4_err_i, s4_rty_i, s5_ack_i, s5_err_i,
         s5_rty_i, s6_ack_i, s6_err_i, s6_rty_i, s7_ack_i, s7_err_i, s7_rty_i,
         s8_ack_i, s8_err_i, s8_rty_i, s9_ack_i, s9_err_i, s9_rty_i, s10_ack_i,
         s10_err_i, s10_rty_i, s11_ack_i, s11_err_i, s11_rty_i, s12_ack_i,
         s12_err_i, s12_rty_i, s13_ack_i, s13_err_i, s13_rty_i, s14_ack_i,
         s14_err_i, s14_rty_i, s15_ack_i, s15_err_i, s15_rty_i;
  output m0_ack_o, m0_err_o, m0_rty_o, m1_ack_o, m1_err_o, m1_rty_o, m2_ack_o,
         m2_err_o, m2_rty_o, m3_ack_o, m3_err_o, m3_rty_o, m4_ack_o, m4_err_o,
         m4_rty_o, m5_ack_o, m5_err_o, m5_rty_o, m6_ack_o, m6_err_o, m6_rty_o,
         m7_ack_o, m7_err_o, m7_rty_o, s0_we_o, s0_cyc_o, s0_stb_o, s1_we_o,
         s1_cyc_o, s1_stb_o, s2_we_o, s2_cyc_o, s2_stb_o, s3_we_o, s3_cyc_o,
         s3_stb_o, s4_we_o, s4_cyc_o, s4_stb_o, s5_we_o, s5_cyc_o, s5_stb_o,
         s6_we_o, s6_cyc_o, s6_stb_o, s7_we_o, s7_cyc_o, s7_stb_o, s8_we_o,
         s8_cyc_o, s8_stb_o, s9_we_o, s9_cyc_o, s9_stb_o, s10_we_o, s10_cyc_o,
         s10_stb_o, s11_we_o, s11_cyc_o, s11_stb_o, s12_we_o, s12_cyc_o,
         s12_stb_o, s13_we_o, s13_cyc_o, s13_stb_o, s14_we_o, s14_cyc_o,
         s14_stb_o, s15_we_o, s15_cyc_o, s15_stb_o;
  wire   m0s0_we, m0s0_cyc, m0s1_cyc, m0s2_cyc, m0s3_cyc, m0s4_cyc, m0s5_cyc,
         m0s6_cyc, m0s7_cyc, m0s8_cyc, m0s9_cyc, m0s10_cyc, m0s11_cyc,
         m0s12_cyc, m0s13_cyc, m0s14_cyc, m0s15_cyc, m1s0_we, m1s0_cyc,
         m1s1_cyc, m1s2_cyc, m1s3_cyc, m1s4_cyc, m1s5_cyc, m1s6_cyc, m1s7_cyc,
         m1s8_cyc, m1s9_cyc, m1s10_cyc, m1s11_cyc, m1s12_cyc, m1s13_cyc,
         m1s14_cyc, m1s15_cyc, m2s0_we, m2s0_cyc, m2s1_cyc, m2s2_cyc, m2s3_cyc,
         m2s4_cyc, m2s5_cyc, m2s6_cyc, m2s7_cyc, m2s8_cyc, m2s9_cyc, m2s10_cyc,
         m2s11_cyc, m2s12_cyc, m2s13_cyc, m2s14_cyc, m2s15_cyc, m3s0_we,
         m3s0_cyc, m3s1_cyc, m3s2_cyc, m3s3_cyc, m3s4_cyc, m3s5_cyc, m3s6_cyc,
         m3s7_cyc, m3s8_cyc, m3s9_cyc, m3s10_cyc, m3s11_cyc, m3s12_cyc,
         m3s13_cyc, m3s14_cyc, m3s15_cyc, m4s0_we, m4s0_cyc, m4s1_cyc,
         m4s2_cyc, m4s3_cyc, m4s4_cyc, m4s5_cyc, m4s6_cyc, m4s7_cyc, m4s8_cyc,
         m4s9_cyc, m4s10_cyc, m4s11_cyc, m4s12_cyc, m4s13_cyc, m4s14_cyc,
         m4s15_cyc, m5s0_we, m5s0_cyc, m5s1_cyc, m5s2_cyc, m5s3_cyc, m5s4_cyc,
         m5s5_cyc, m5s6_cyc, m5s7_cyc, m5s8_cyc, m5s9_cyc, m5s10_cyc,
         m5s11_cyc, m5s12_cyc, m5s13_cyc, m5s14_cyc, m5s15_cyc, m6s0_we,
         m6s0_cyc, m6s1_cyc, m6s2_cyc, m6s3_cyc, m6s4_cyc, m6s5_cyc, m6s6_cyc,
         m6s7_cyc, m6s8_cyc, m6s9_cyc, m6s10_cyc, m6s11_cyc, m6s12_cyc,
         m6s13_cyc, m6s14_cyc, m6s15_cyc, m7s0_we, m7s0_cyc, m7s1_cyc,
         m7s2_cyc, m7s3_cyc, m7s4_cyc, m7s5_cyc, m7s6_cyc, m7s7_cyc, m7s8_cyc,
         m7s9_cyc, m7s10_cyc, m7s11_cyc, m7s12_cyc, m7s13_cyc, m7s14_cyc,
         m7s15_cyc, \s0/m7_cyc_r , \s0/m6_cyc_r , \s0/m5_cyc_r , \s0/m4_cyc_r ,
         \s0/m3_cyc_r , \s0/m2_cyc_r , \s0/m1_cyc_r , \s0/m0_cyc_r , \s0/next ,
         \s1/m7_cyc_r , \s1/m6_cyc_r , \s1/m5_cyc_r , \s1/m4_cyc_r ,
         \s1/m3_cyc_r , \s1/m2_cyc_r , \s1/m1_cyc_r , \s1/m0_cyc_r , \s1/next ,
         \s2/m7_cyc_r , \s2/m6_cyc_r , \s2/m5_cyc_r , \s2/m4_cyc_r ,
         \s2/m3_cyc_r , \s2/m2_cyc_r , \s2/m1_cyc_r , \s2/m0_cyc_r , \s2/next ,
         \s3/m7_cyc_r , \s3/m6_cyc_r , \s3/m5_cyc_r , \s3/m4_cyc_r ,
         \s3/m3_cyc_r , \s3/m2_cyc_r , \s3/m1_cyc_r , \s3/m0_cyc_r , \s3/next ,
         \s4/m7_cyc_r , \s4/m6_cyc_r , \s4/m5_cyc_r , \s4/m4_cyc_r ,
         \s4/m3_cyc_r , \s4/m2_cyc_r , \s4/m1_cyc_r , \s4/m0_cyc_r , \s4/next ,
         \s5/m7_cyc_r , \s5/m6_cyc_r , \s5/m5_cyc_r , \s5/m4_cyc_r ,
         \s5/m3_cyc_r , \s5/m2_cyc_r , \s5/m1_cyc_r , \s5/m0_cyc_r , \s5/next ,
         \s6/m7_cyc_r , \s6/m6_cyc_r , \s6/m5_cyc_r , \s6/m4_cyc_r ,
         \s6/m3_cyc_r , \s6/m2_cyc_r , \s6/m1_cyc_r , \s6/m0_cyc_r , \s6/next ,
         \s7/m7_cyc_r , \s7/m6_cyc_r , \s7/m5_cyc_r , \s7/m4_cyc_r ,
         \s7/m3_cyc_r , \s7/m2_cyc_r , \s7/m1_cyc_r , \s7/m0_cyc_r , \s7/next ,
         \s8/m7_cyc_r , \s8/m6_cyc_r , \s8/m5_cyc_r , \s8/m4_cyc_r ,
         \s8/m3_cyc_r , \s8/m2_cyc_r , \s8/m1_cyc_r , \s8/m0_cyc_r , \s8/next ,
         \s9/m7_cyc_r , \s9/m6_cyc_r , \s9/m5_cyc_r , \s9/m4_cyc_r ,
         \s9/m3_cyc_r , \s9/m2_cyc_r , \s9/m1_cyc_r , \s9/m0_cyc_r , \s9/next ,
         \s10/m7_cyc_r , \s10/m6_cyc_r , \s10/m5_cyc_r , \s10/m4_cyc_r ,
         \s10/m3_cyc_r , \s10/m2_cyc_r , \s10/m1_cyc_r , \s10/m0_cyc_r ,
         \s10/next , \s11/m7_cyc_r , \s11/m6_cyc_r , \s11/m5_cyc_r ,
         \s11/m4_cyc_r , \s11/m3_cyc_r , \s11/m2_cyc_r , \s11/m1_cyc_r ,
         \s11/m0_cyc_r , \s11/next , \s12/m7_cyc_r , \s12/m6_cyc_r ,
         \s12/m5_cyc_r , \s12/m4_cyc_r , \s12/m3_cyc_r , \s12/m2_cyc_r ,
         \s12/m1_cyc_r , \s12/m0_cyc_r , \s12/next , \s13/m7_cyc_r ,
         \s13/m6_cyc_r , \s13/m5_cyc_r , \s13/m4_cyc_r , \s13/m3_cyc_r ,
         \s13/m2_cyc_r , \s13/m1_cyc_r , \s13/m0_cyc_r , \s13/next ,
         \s14/m7_cyc_r , \s14/m6_cyc_r , \s14/m5_cyc_r , \s14/m4_cyc_r ,
         \s14/m3_cyc_r , \s14/m2_cyc_r , \s14/m1_cyc_r , \s14/m0_cyc_r ,
         \s14/next , \s15/m7_cyc_r , \s15/m6_cyc_r , \s15/m5_cyc_r ,
         \s15/m4_cyc_r , \s15/m3_cyc_r , \s15/m2_cyc_r , \s15/m1_cyc_r ,
         \s15/m0_cyc_r , \s15/next , \rf/N130 , \rf/N129 , \rf/N128 ,
         \rf/N127 , \rf/N126 , \rf/N125 , \rf/N124 , \rf/N123 , \rf/N122 ,
         \rf/N121 , \rf/N120 , \rf/N119 , \rf/N118 , \rf/N117 , \rf/N116 ,
         \rf/N115 , \rf/N19 , \rf/rf_ack , \rf/N18 , n13464, n13465, n13469,
         n13470, n13471, n13472, n13474, n13475, n13481, n13482, n13484,
         n13485, n13489, n13490, n13494, n13495, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13888, n13890, n13892,
         n13894, n13896, n13898, n13900, n13902, n13908, n13910, n13912,
         n13914, n13916, n13918, n13920, n13922, n17568, n17569, n17570,
         n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578,
         n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586,
         n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594,
         n17595, n17596, n17597, n17598, n17599, n17601, n17603, n17604,
         n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612,
         n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620,
         n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628,
         n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636,
         n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644,
         n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652,
         n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660,
         n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668,
         n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676,
         n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684,
         n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692,
         n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700,
         n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708,
         n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716,
         n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724,
         n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732,
         n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740,
         n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748,
         n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756,
         n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764,
         n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772,
         n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780,
         n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788,
         n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796,
         n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804,
         n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812,
         n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820,
         n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828,
         n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836,
         n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844,
         n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852,
         n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860,
         n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868,
         n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876,
         n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884,
         n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892,
         n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900,
         n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908,
         n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916,
         n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924,
         n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932,
         n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940,
         n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948,
         n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956,
         n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964,
         n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972,
         n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980,
         n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988,
         n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996,
         n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004,
         n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012,
         n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020,
         n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028,
         n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036,
         n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044,
         n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052,
         n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060,
         n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068,
         n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076,
         n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084,
         n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092,
         n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100,
         n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108,
         n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116,
         n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124,
         n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132,
         n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140,
         n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148,
         n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156,
         n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164,
         n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172,
         n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180,
         n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188,
         n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196,
         n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204,
         n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212,
         n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220,
         n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228,
         n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236,
         n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244,
         n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252,
         n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260,
         n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268,
         n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276,
         n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284,
         n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292,
         n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300,
         n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308,
         n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316,
         n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324,
         n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332,
         n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340,
         n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348,
         n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356,
         n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364,
         n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372,
         n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380,
         n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388,
         n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396,
         n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404,
         n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412,
         n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420,
         n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428,
         n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436,
         n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444,
         n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452,
         n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460,
         n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468,
         n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476,
         n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484,
         n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492,
         n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500,
         n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508,
         n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516,
         n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524,
         n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532,
         n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540,
         n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548,
         n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556,
         n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564,
         n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572,
         n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580,
         n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588,
         n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596,
         n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604,
         n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612,
         n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620,
         n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628,
         n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636,
         n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644,
         n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652,
         n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660,
         n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668,
         n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676,
         n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684,
         n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692,
         n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700,
         n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708,
         n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716,
         n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724,
         n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732,
         n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740,
         n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748,
         n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756,
         n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764,
         n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772,
         n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780,
         n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788,
         n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796,
         n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804,
         n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812,
         n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820,
         n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828,
         n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836,
         n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844,
         n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852,
         n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860,
         n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868,
         n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876,
         n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884,
         n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892,
         n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900,
         n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908,
         n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916,
         n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924,
         n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932,
         n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940,
         n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948,
         n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956,
         n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964,
         n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972,
         n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980,
         n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988,
         n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996,
         n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004,
         n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012,
         n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020,
         n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028,
         n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036,
         n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044,
         n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052,
         n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060,
         n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068,
         n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076,
         n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084,
         n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092,
         n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100,
         n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108,
         n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116,
         n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124,
         n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132,
         n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140,
         n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148,
         n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156,
         n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164,
         n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172,
         n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180,
         n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188,
         n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196,
         n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204,
         n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212,
         n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220,
         n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228,
         n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236,
         n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244,
         n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252,
         n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260,
         n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268,
         n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276,
         n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284,
         n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292,
         n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300,
         n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308,
         n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316,
         n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324,
         n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332,
         n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340,
         n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348,
         n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356,
         n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364,
         n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372,
         n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380,
         n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388,
         n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396,
         n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404,
         n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412,
         n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420,
         n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428,
         n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436,
         n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444,
         n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452,
         n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460,
         n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468,
         n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476,
         n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484,
         n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492,
         n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500,
         n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508,
         n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516,
         n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524,
         n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532,
         n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540,
         n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548,
         n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556,
         n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564,
         n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572,
         n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580,
         n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588,
         n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596,
         n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604,
         n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612,
         n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620,
         n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628,
         n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636,
         n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644,
         n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652,
         n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660,
         n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668,
         n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676,
         n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684,
         n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692,
         n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700,
         n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708,
         n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716,
         n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724,
         n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732,
         n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740,
         n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748,
         n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756,
         n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764,
         n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772,
         n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780,
         n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788,
         n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796,
         n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804,
         n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812,
         n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820,
         n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828,
         n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836,
         n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844,
         n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852,
         n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860,
         n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868,
         n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876,
         n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884,
         n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892,
         n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900,
         n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908,
         n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916,
         n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924,
         n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932,
         n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940,
         n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948,
         n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956,
         n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964,
         n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972,
         n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980,
         n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988,
         n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996,
         n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004,
         n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012,
         n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020,
         n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028,
         n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036,
         n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044,
         n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052,
         n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060,
         n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068,
         n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076,
         n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084,
         n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092,
         n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100,
         n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108,
         n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116,
         n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124,
         n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132,
         n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140,
         n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148,
         n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156,
         n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164,
         n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172,
         n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180,
         n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188,
         n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196,
         n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204,
         n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212,
         n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220,
         n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228,
         n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236,
         n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244,
         n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252,
         n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260,
         n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268,
         n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276,
         n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284,
         n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292,
         n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300,
         n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308,
         n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316,
         n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324,
         n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332,
         n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340,
         n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348,
         n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356,
         n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364,
         n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372,
         n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380,
         n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388,
         n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396,
         n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404,
         n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412,
         n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420,
         n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428,
         n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436,
         n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444,
         n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452,
         n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460,
         n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468,
         n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476,
         n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484,
         n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492,
         n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500,
         n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508,
         n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516,
         n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524,
         n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532,
         n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540,
         n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548,
         n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556,
         n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564,
         n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572,
         n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580,
         n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588,
         n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596,
         n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604,
         n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612,
         n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620,
         n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628,
         n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636,
         n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644,
         n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652,
         n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660,
         n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668,
         n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676,
         n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684,
         n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692,
         n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700,
         n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708,
         n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716,
         n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724,
         n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732,
         n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740,
         n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748,
         n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756,
         n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764,
         n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772,
         n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780,
         n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788,
         n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796,
         n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804,
         n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812,
         n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820,
         n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828,
         n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836,
         n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844,
         n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852,
         n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860,
         n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868,
         n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876,
         n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884,
         n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892,
         n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900,
         n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908,
         n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916,
         n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924,
         n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932,
         n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940,
         n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948,
         n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956,
         n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964,
         n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972,
         n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980,
         n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988,
         n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996,
         n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004,
         n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012,
         n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020,
         n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028,
         n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036,
         n21037, n21038, n21039, n21040, n21041, n21042, n21043, n21044,
         n21045, n21046, n21047, n21048, n21049, n21050, n21051, n21052,
         n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060,
         n21061, n21062, n21063, n21064, n21065, n21066, n21067, n21068,
         n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076,
         n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084,
         n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092,
         n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100,
         n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108,
         n21109, n21110, n21111, n21112, n21113, n21114, n21115, n21116,
         n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124,
         n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132,
         n21133, n21134, n21135, n21136, n21137, n21138, n21139, n21140,
         n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148,
         n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156,
         n21157, n21158, n21159, n21160, n21161, n21162, n21163, n21164,
         n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172,
         n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180,
         n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188,
         n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196,
         n21197, n21198, n21199, n21200, n21201, n21202, n21203, n21204,
         n21205, n21206, n21207, n21208, n21209, n21210, n21211, n21212,
         n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220,
         n21221, n21222, n21223, n21224, n21225, n21226, n21227, n21228,
         n21229, n21230, n21231, n21232, n21233, n21234, n21235, n21236,
         n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244,
         n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252,
         n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260,
         n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268,
         n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21276,
         n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284,
         n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292,
         n21293, n21294, n21295, n21296, n21297, n21298, n21299, n21300,
         n21301, n21302, n21303, n21304, n21305, n21306, n21307, n21308,
         n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316,
         n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324,
         n21325, n21326, n21327, n21328, n21329, n21330, n21331, n21332,
         n21333, n21334, n21335, n21336, n21337, n21338, n21339, n21340,
         n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348,
         n21349, n21350, n21351, n21352, n21353, n21354, n21355, n21356,
         n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364,
         n21365, n21366, n21367, n21368, n21369, n21370, n21371, n21372,
         n21373, n21374, n21375, n21376, n21377, n21378, n21379, n21380,
         n21381, n21382, n21383, n21384, n21385, n21386, n21387, n21388,
         n21389, n21390, n21391, n21392, n21393, n21394, n21395, n21396,
         n21397, n21398, n21399, n21400, n21401, n21402, n21403, n21404,
         n21405, n21406, n21407, n21408, n21409, n21410, n21411, n21412,
         n21413, n21414, n21415, n21416, n21417, n21418, n21419, n21420,
         n21421, n21422, n21423, n21424, n21425, n21426, n21427, n21428,
         n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436,
         n21437, n21438, n21439, n21440, n21441, n21442, n21443, n21444,
         n21445, n21446, n21447, n21448, n21449, n21450, n21451, n21452,
         n21453, n21454, n21455, n21456, n21457, n21458, n21459, n21460,
         n21461, n21462, n21463, n21464, n21465, n21466, n21467, n21468,
         n21469, n21470, n21471, n21472, n21473, n21474, n21475, n21476,
         n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484,
         n21485, n21486, n21487, n21488, n21489, n21490, n21491, n21492,
         n21493, n21494, n21495, n21496, n21497, n21498, n21499, n21500,
         n21501, n21502, n21503, n21504, n21505, n21506, n21507, n21508,
         n21509, n21510, n21511, n21512, n21513, n21514, n21515, n21516,
         n21517, n21518, n21519, n21520, n21521, n21522, n21523, n21524,
         n21525, n21526, n21527, n21528, n21529, n21530, n21531, n21532,
         n21533, n21534, n21535, n21536, n21537, n21538, n21539, n21540,
         n21541, n21542, n21543, n21544, n21545, n21546, n21547, n21548,
         n21549, n21550, n21551, n21552, n21553, n21554, n21555, n21556,
         n21557, n21558, n21559, n21560, n21561, n21562, n21563, n21564,
         n21565, n21566, n21567, n21568, n21569, n21570, n21571, n21572,
         n21573, n21574, n21575, n21576, n21577, n21578, n21579, n21580,
         n21581, n21582, n21583, n21584, n21585, n21586, n21587, n21588,
         n21589, n21590, n21591, n21592, n21593, n21594, n21595, n21596,
         n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604,
         n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612,
         n21613, n21614, n21615, n21616, n21617, n21618, n21619, n21620,
         n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628,
         n21629, n21630, n21631, n21632, n21633, n21634, n21635, n21636,
         n21637, n21638, n21639, n21640, n21641, n21642, n21643, n21644,
         n21645, n21646, n21647, n21648, n21649, n21650, n21651, n21652,
         n21653, n21654, n21655, n21656, n21657, n21658, n21659, n21660,
         n21661, n21662, n21663, n21664, n21665, n21666, n21667, n21668,
         n21669, n21670, n21671, n21672, n21673, n21674, n21675, n21676,
         n21677, n21678, n21679, n21680, n21681, n21682, n21683, n21684,
         n21685, n21686, n21687, n21688, n21689, n21690, n21691, n21692,
         n21693, n21694, n21695, n21696, n21697, n21698, n21699, n21700,
         n21701, n21702, n21703, n21704, n21705, n21706, n21707, n21708,
         n21709, n21710, n21711, n21712, n21713, n21714, n21715, n21716,
         n21717, n21718, n21719, n21720, n21721, n21722, n21723, n21724,
         n21725, n21726, n21727, n21728, n21729, n21730, n21731, n21732,
         n21733, n21734, n21735, n21736, n21737, n21738, n21739, n21740,
         n21741, n21742, n21743, n21744, n21745, n21746, n21747, n21748,
         n21749, n21750, n21751, n21752, n21753, n21754, n21755, n21756,
         n21757, n21758, n21759, n21760, n21761, n21762, n21763, n21764,
         n21765, n21766, n21767, n21768, n21769, n21770, n21771, n21772,
         n21773, n21774, n21775, n21776, n21777, n21778, n21779, n21780,
         n21781, n21782, n21783, n21784, n21785, n21786, n21787, n21788,
         n21789, n21790, n21791, n21792, n21793, n21794, n21795, n21796,
         n21797, n21798, n21799, n21800, n21801, n21802, n21803, n21804,
         n21805, n21806, n21807, n21808, n21809, n21810, n21811, n21812,
         n21813, n21814, n21815, n21816, n21817, n21818, n21819, n21820,
         n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828,
         n21829, n21830, n21831, n21832, n21833, n21834, n21835, n21836,
         n21837, n21838, n21839, n21840, n21841, n21842, n21843, n21844,
         n21845, n21846, n21847, n21848, n21849, n21850, n21851, n21852,
         n21853, n21854, n21855, n21856, n21857, n21858, n21859, n21860,
         n21861, n21862, n21863, n21864, n21865, n21866, n21867, n21868,
         n21869, n21870, n21871, n21872, n21873, n21874, n21875, n21876,
         n21877, n21878, n21879, n21880, n21881, n21882, n21883, n21884,
         n21885, n21886, n21887, n21888, n21889, n21890, n21891, n21892,
         n21893, n21894, n21895, n21896, n21897, n21898, n21899, n21900,
         n21901, n21902, n21903, n21904, n21905, n21906, n21907, n21908,
         n21909, n21910, n21911, n21912, n21913, n21914, n21915, n21916,
         n21917, n21918, n21919, n21920, n21921, n21922, n21923, n21924,
         n21925, n21926, n21927, n21928, n21929, n21930, n21931, n21932,
         n21933, n21934, n21935, n21936, n21937, n21938, n21939, n21940,
         n21941, n21942, n21943, n21944, n21945, n21946, n21947, n21948,
         n21949, n21950, n21951, n21952, n21953, n21954, n21955, n21956,
         n21957, n21958, n21959, n21960, n21961, n21962, n21963, n21964,
         n21965, n21966, n21967, n21968, n21969, n21970, n21971, n21972,
         n21973, n21974, n21975, n21976, n21977, n21978, n21979, n21980,
         n21981, n21982, n21983, n21984, n21985, n21986, n21987, n21988,
         n21989, n21990, n21991, n21992, n21993, n21994, n21995, n21996,
         n21997, n21998, n21999, n22000, n22001, n22002, n22003, n22004,
         n22005, n22006, n22007, n22008, n22009, n22010, n22011, n22012,
         n22013, n22014, n22015, n22016, n22017, n22018, n22019, n22020,
         n22021, n22022, n22023, n22024, n22025, n22026, n22027, n22028,
         n22029, n22030, n22031, n22032, n22033, n22034, n22035, n22036,
         n22037, n22038, n22039, n22040, n22041, n22042, n22043, n22044,
         n22045, n22046, n22047, n22048, n22049, n22050, n22051, n22052,
         n22053, n22054, n22055, n22056, n22057, n22058, n22059, n22060,
         n22061, n22062, n22063, n22064, n22065, n22066, n22067, n22068,
         n22069, n22070, n22071, n22072, n22073, n22074, n22075, n22076,
         n22077, n22078, n22079, n22080, n22081, n22082, n22083, n22084,
         n22085, n22086, n22087, n22088, n22089, n22090, n22091, n22092,
         n22093, n22094, n22095, n22096, n22097, n22098, n22099, n22100,
         n22101, n22102, n22103, n22104, n22105, n22106, n22107, n22108,
         n22109, n22110, n22111, n22112, n22113, n22114, n22115, n22116,
         n22117, n22118, n22119, n22120, n22121, n22122, n22123, n22124,
         n22125, n22126, n22127, n22128, n22129, n22130, n22131, n22132,
         n22133, n22134, n22135, n22136, n22137, n22138, n22139, n22140,
         n22141, n22142, n22143, n22144, n22145, n22146, n22147, n22148,
         n22149, n22150, n22151, n22152, n22153, n22154, n22155, n22156,
         n22157, n22158, n22159, n22160, n22161, n22162, n22163, n22164,
         n22165, n22166, n22167, n22168, n22169, n22170, n22171, n22172,
         n22173, n22174, n22175, n22176, n22177, n22178, n22179, n22180,
         n22181, n22182, n22183, n22184, n22185, n22186, n22187, n22188,
         n22189, n22190, n22191, n22192, n22193, n22194, n22195, n22196,
         n22197, n22198, n22199, n22200, n22201, n22202, n22203, n22204,
         n22205, n22206, n22207, n22208, n22209, n22210, n22211, n22212,
         n22213, n22214, n22215, n22216, n22217, n22218, n22219, n22220,
         n22221, n22222, n22223, n22224, n22225, n22226, n22227, n22228,
         n22229, n22230, n22231, n22232, n22233, n22234, n22235, n22236,
         n22237, n22238, n22239, n22240, n22241, n22242, n22243, n22244,
         n22245, n22246, n22247, n22248, n22249, n22250, n22251, n22252,
         n22253, n22254, n22255, n22256, n22257, n22258, n22259, n22260,
         n22261, n22262, n22263, n22264, n22265, n22266, n22267, n22268,
         n22269, n22270, n22271, n22272, n22273, n22274, n22275, n22276,
         n22277, n22278, n22279, n22280, n22281, n22282, n22283, n22284,
         n22285, n22286, n22287, n22288, n22289, n22290, n22291, n22292,
         n22293, n22294, n22295, n22296, n22297, n22298, n22299, n22300,
         n22301, n22302, n22303, n22304, n22305, n22306, n22307, n22308,
         n22309, n22310, n22311, n22312, n22313, n22314, n22315, n22316,
         n22317, n22318, n22319, n22320, n22321, n22322, n22323, n22324,
         n22325, n22326, n22327, n22328, n22329, n22330, n22331, n22332,
         n22333, n22334, n22335, n22336, n22337, n22338, n22339, n22340,
         n22341, n22342, n22343, n22344, n22345, n22346, n22347, n22348,
         n22349, n22350, n22351, n22352, n22353, n22354, n22355, n22356,
         n22357, n22358, n22359, n22360, n22361, n22362, n22363, n22364,
         n22365, n22366, n22367, n22368, n22369, n22370, n22371, n22372,
         n22373, n22374, n22375, n22376, n22377, n22378, n22379, n22380,
         n22381, n22382, n22383, n22384, n22385, n22386, n22387, n22388,
         n22389, n22390, n22391, n22392, n22393, n22394, n22395, n22396,
         n22397, n22398, n22399, n22400, n22401, n22402, n22403, n22404,
         n22405, n22406, n22407, n22408, n22409, n22410, n22411, n22412,
         n22413, n22414, n22415, n22416, n22417, n22418, n22419, n22420,
         n22421, n22422, n22423, n22424, n22425, n22426, n22427, n22428,
         n22429, n22430, n22431, n22432, n22433, n22434, n22435, n22436,
         n22437, n22438, n22439, n22440, n22441, n22442, n22443, n22444,
         n22445, n22446, n22447, n22448, n22449, n22450, n22451, n22452,
         n22453, n22454, n22455, n22456, n22457, n22458, n22459, n22460,
         n22461, n22462, n22463, n22464, n22465, n22466, n22467, n22468,
         n22469, n22470, n22471, n22472, n22473, n22474, n22475, n22476,
         n22477, n22478, n22479, n22480, n22481, n22482, n22483, n22484,
         n22485, n22486, n22487, n22488, n22489, n22490, n22491, n22492,
         n22493, n22494, n22495, n22496, n22497, n22498, n22499, n22500,
         n22501, n22502, n22503, n22504, n22505, n22506, n22507, n22508,
         n22509, n22510, n22511, n22512, n22513, n22514, n22515, n22516,
         n22517, n22518, n22519, n22520, n22521, n22522, n22523, n22524,
         n22525, n22526, n22527, n22528, n22529, n22530, n22531, n22532,
         n22533, n22534, n22535, n22536, n22537, n22538, n22539, n22540,
         n22541, n22542, n22543, n22544, n22545, n22546, n22547, n22548,
         n22549, n22550, n22551, n22552, n22553, n22554, n22555, n22556,
         n22557, n22558, n22559, n22560, n22561, n22562, n22563, n22564,
         n22565, n22566, n22567, n22568, n22569, n22570, n22571, n22572,
         n22573, n22574, n22575, n22576, n22577, n22578, n22579, n22580,
         n22581, n22582, n22583, n22584, n22585, n22586, n22587, n22588,
         n22589, n22590, n22591, n22592, n22593, n22594, n22595, n22596,
         n22597, n22598, n22599, n22600, n22601, n22602, n22603, n22604,
         n22605, n22606, n22607, n22608, n22609, n22610, n22611, n22612,
         n22613, n22614, n22615, n22616, n22617, n22618, n22619, n22620,
         n22621, n22622, n22623, n22624, n22625, n22626, n22627, n22628,
         n22629, n22630, n22631, n22632, n22633, n22634, n22635, n22636,
         n22637, n22638, n22639, n22640, n22641, n22642, n22643, n22644,
         n22645, n22646, n22647, n22648, n22649, n22650, n22651, n22652,
         n22653, n22654, n22655, n22656, n22657, n22658, n22659, n22660,
         n22661, n22662, n22663, n22664, n22665, n22666, n22667, n22668,
         n22669, n22670, n22671, n22672, n22673, n22674, n22675, n22676,
         n22677, n22678, n22679, n22680, n22681, n22682, n22683, n22684,
         n22685, n22686, n22687, n22688, n22689, n22690, n22691, n22692,
         n22693, n22694, n22695, n22696, n22697, n22698, n22699, n22700,
         n22701, n22702, n22703, n22704, n22705, n22706, n22707, n22708,
         n22709, n22710, n22711, n22712, n22713, n22714, n22715, n22716,
         n22717, n22718, n22719, n22720, n22721, n22722, n22723, n22724,
         n22725, n22726, n22727, n22728, n22729, n22730, n22731, n22732,
         n22733, n22734, n22735, n22736, n22737, n22738, n22739, n22740,
         n22741, n22742, n22743, n22744, n22745, n22746, n22747, n22748,
         n22749, n22750, n22751, n22752, n22753, n22754, n22755, n22756,
         n22757, n22758, n22759, n22760, n22761, n22762, n22763, n22764,
         n22765, n22766, n22767, n22768, n22769, n22770, n22771, n22772,
         n22773, n22774, n22775, n22776, n22777, n22778, n22779, n22780,
         n22781, n22782, n22783, n22784, n22785, n22786, n22787, n22788,
         n22789, n22790, n22791, n22792, n22793, n22794, n22795, n22796,
         n22797, n22798, n22799, n22800, n22801, n22802, n22803, n22804,
         n22805, n22806, n22807, n22808, n22809, n22810, n22811, n22812,
         n22813, n22814, n22815, n22816, n22817, n22818, n22819, n22820,
         n22821, n22822, n22823, n22824, n22825, n22826, n22827, n22828,
         n22829, n22830, n22831, n22832, n22833, n22834, n22835, n22836,
         n22837, n22838, n22839, n22840, n22841, n22842, n22843, n22844,
         n22845, n22846, n22847, n22848, n22849, n22850, n22851, n22852,
         n22853, n22854, n22855, n22856, n22857, n22858, n22859, n22860,
         n22861, n22862, n22863, n22864, n22865, n22866, n22867, n22868,
         n22869, n22870, n22871, n22872, n22873, n22874, n22875, n22876,
         n22877, n22878, n22879, n22880, n22881, n22882, n22883, n22884,
         n22885, n22886, n22887, n22888, n22889, n22890, n22891, n22892,
         n22893, n22894, n22895, n22896, n22897, n22898, n22899, n22900,
         n22901, n22902, n22903, n22904, n22905, n22906, n22907, n22908,
         n22909, n22910, n22911, n22912, n22913, n22914, n22915, n22916,
         n22917, n22918, n22919, n22920, n22921, n22922, n22923, n22924,
         n22925, n22926, n22927, n22928, n22929, n22930, n22931, n22932,
         n22933, n22934, n22935, n22936, n22937, n22938, n22939, n22940,
         n22941, n22942, n22943, n22944, n22945, n22946, n22947, n22948,
         n22949, n22950, n22951, n22952, n22953, n22954, n22955, n22956,
         n22957, n22958, n22959, n22960, n22961, n22962, n22963, n22964,
         n22965, n22966, n22967, n22968, n22969, n22970, n22971, n22972,
         n22973, n22974, n22975, n22976, n22977, n22978, n22979, n22980,
         n22981, n22982, n22983, n22984, n22985, n22986, n22987, n22988,
         n22989, n22990, n22991, n22992, n22993, n22994, n22995, n22996,
         n22997, n22998, n22999, n23000, n23001, n23002, n23003, n23004,
         n23005, n23006, n23007, n23008, n23009, n23010, n23011, n23012,
         n23013, n23014, n23015, n23016, n23017, n23018, n23019, n23020,
         n23021, n23022, n23023, n23024, n23025, n23026, n23027, n23028,
         n23029, n23030, n23031, n23032, n23033, n23034, n23035, n23036,
         n23037, n23038, n23039, n23040, n23041, n23042, n23043, n23044,
         n23045, n23046, n23047, n23048, n23049, n23050, n23051, n23052,
         n23053, n23054, n23055, n23056, n23057, n23058, n23059, n23060,
         n23061, n23062, n23063, n23064, n23065, n23066, n23067, n23068,
         n23069, n23070, n23071, n23072, n23073, n23074, n23075, n23076,
         n23077, n23078, n23079, n23080, n23081, n23082, n23083, n23084,
         n23085, n23086, n23087, n23088, n23089, n23090, n23091, n23092,
         n23093, n23094, n23095, n23096, n23097, n23098, n23099, n23100,
         n23101, n23102, n23103, n23104, n23105, n23106, n23107, n23108,
         n23109, n23110, n23111, n23112, n23113, n23114, n23115, n23116,
         n23117, n23118, n23119, n23120, n23121, n23122, n23123, n23124,
         n23125, n23126, n23127, n23128, n23129, n23130, n23131, n23132,
         n23133, n23134, n23135, n23136, n23137, n23138, n23139, n23140,
         n23141, n23142, n23143, n23144, n23145, n23146, n23147, n23148,
         n23149, n23150, n23151, n23152, n23153, n23154, n23155, n23156,
         n23157, n23158, n23159, n23160, n23161, n23162, n23163, n23164,
         n23165, n23166, n23167, n23168, n23169, n23170, n23171, n23172,
         n23173, n23174, n23175, n23176, n23177, n23178, n23179, n23180,
         n23181, n23182, n23183, n23184, n23185, n23186, n23187, n23188,
         n23189, n23190, n23191, n23192, n23193, n23194, n23195, n23196,
         n23197, n23198, n23199, n23200, n23201, n23202, n23203, n23204,
         n23205, n23206, n23207, n23208, n23209, n23210, n23211, n23212,
         n23213, n23214, n23215, n23216, n23217, n23218, n23219, n23220,
         n23221, n23222, n23223, n23224, n23225, n23226, n23227, n23228,
         n23229, n23230, n23231, n23232, n23233, n23234, n23235, n23236,
         n23237, n23238, n23239, n23240, n23241, n23242, n23243, n23244,
         n23245, n23246, n23247, n23248, n23249, n23250, n23251, n23252,
         n23253, n23254, n23255, n23256, n23257, n23258, n23259, n23260,
         n23261, n23262, n23263, n23264, n23265, n23266, n23267, n23268,
         n23269, n23270, n23271, n23272, n23273, n23274, n23275, n23276,
         n23277, n23278, n23279, n23280, n23281, n23282, n23283, n23284,
         n23285, n23286, n23287, n23288, n23289, n23290, n23291, n23292,
         n23293, n23294, n23295, n23296, n23297, n23298, n23299, n23300,
         n23301, n23302, n23303, n23304, n23305, n23306, n23307, n23308,
         n23309, n23310, n23311, n23312, n23313, n23314, n23315, n23316,
         n23317, n23318, n23319, n23320, n23321, n23322, n23323, n23324,
         n23325, n23326, n23327, n23328, n23329, n23330, n23331, n23332,
         n23333, n23334, n23335, n23336, n23337, n23338, n23339, n23340,
         n23341, n23342, n23343, n23344, n23345, n23346, n23347, n23348,
         n23349, n23350, n23351, n23352, n23353, n23354, n23355, n23356,
         n23357, n23358, n23359, n23360, n23361, n23362, n23363, n23364,
         n23365, n23366, n23367, n23368, n23369, n23370, n23371, n23372,
         n23373, n23374, n23375, n23376, n23377, n23378, n23379, n23380,
         n23381, n23382, n23383, n23384, n23385, n23386, n23387, n23388,
         n23389, n23390, n23391, n23392, n23393, n23394, n23395, n23396,
         n23397, n23398, n23399, n23400, n23401, n23402, n23403, n23404,
         n23405, n23406, n23407, n23408, n23409, n23410, n23411, n23412,
         n23413, n23414, n23415, n23416, n23417, n23418, n23419, n23420,
         n23421, n23422, n23423, n23424, n23425, n23426, n23427, n23428,
         n23429, n23430, n23431, n23432, n23433, n23434, n23435, n23436,
         n23437, n23438, n23439, n23440, n23441, n23442, n23443, n23444,
         n23445, n23446, n23447, n23448, n23449, n23450, n23451, n23452,
         n23453, n23454, n23455, n23456, n23457, n23458, n23459, n23460,
         n23461, n23462, n23463, n23464, n23465, n23466, n23467, n23468,
         n23469, n23470, n23471, n23472, n23473, n23474, n23475, n23476,
         n23477, n23478, n23479, n23480, n23481, n23482, n23483, n23484,
         n23485, n23486, n23487, n23488, n23489, n23490, n23491, n23492,
         n23493, n23494, n23495, n23496, n23497, n23498, n23499, n23500,
         n23501, n23502, n23503, n23504, n23505, n23506, n23507, n23508,
         n23509, n23510, n23511, n23512, n23513, n23514, n23515, n23516,
         n23517, n23518, n23519, n23520, n23521, n23522, n23523, n23524,
         n23525, n23526, n23527, n23528, n23529, n23530, n23531, n23532,
         n23533, n23534, n23535, n23536, n23537, n23538, n23539, n23540,
         n23541, n23542, n23543, n23544, n23545, n23546, n23547, n23548,
         n23549, n23550, n23551, n23552, n23553, n23554, n23555, n23556,
         n23557, n23558, n23559, n23560, n23561, n23562, n23563, n23564,
         n23565, n23566, n23567, n23568, n23569, n23570, n23571, n23572,
         n23573, n23574, n23575, n23576, n23577, n23578, n23579, n23580,
         n23581, n23582, n23583, n23584, n23585, n23586, n23587, n23588,
         n23589, n23590, n23591, n23592, n23593, n23594, n23595, n23596,
         n23597, n23598, n23599, n23600, n23601, n23602, n23603, n23604,
         n23605, n23606, n23607, n23608, n23609, n23610, n23611, n23612,
         n23613, n23614, n23615, n23616, n23617, n23618, n23619, n23620,
         n23621, n23622, n23623, n23624, n23625, n23626, n23627, n23628,
         n23629, n23630, n23631, n23632, n23633, n23634, n23635, n23636,
         n23637, n23638, n23639, n23640, n23641, n23642, n23643, n23644,
         n23645, n23646, n23647, n23648, n23649, n23650, n23651, n23652,
         n23653, n23654, n23655, n23656, n23657, n23658, n23659, n23660,
         n23661, n23662, n23663, n23664, n23665, n23666, n23667, n23668,
         n23669, n23670, n23671, n23672, n23673, n23674, n23675, n23676,
         n23677, n23678, n23679, n23680, n23681, n23682, n23683, n23684,
         n23685, n23686, n23687, n23688, n23689, n23690, n23691, n23692,
         n23693, n23694, n23695, n23696, n23697, n23698, n23699, n23700,
         n23701, n23702, n23703, n23704, n23705, n23706, n23707, n23708,
         n23709, n23710, n23711, n23712, n23713, n23714, n23715, n23716,
         n23717, n23718, n23719, n23720, n23721, n23722, n23723, n23724,
         n23725, n23726, n23727, n23728, n23729, n23730, n23731, n23732,
         n23733, n23734, n23735, n23736, n23737, n23738, n23739, n23740,
         n23741, n23742, n23743, n23744, n23745, n23746, n23747, n23748,
         n23749, n23750, n23751, n23752, n23753, n23754, n23755, n23756,
         n23757, n23758, n23759, n23760, n23761, n23762, n23763, n23764,
         n23765, n23766, n23767, n23768, n23769, n23770, n23771, n23772,
         n23773, n23774, n23775, n23776, n23777, n23778, n23779, n23780,
         n23781, n23782, n23783, n23784, n23785, n23786, n23787, n23788,
         n23789, n23790, n23791, n23792, n23793, n23794, n23795, n23796,
         n23797, n23798, n23799, n23800, n23801, n23802, n23803, n23804,
         n23805, n23806, n23807, n23808, n23809, n23810, n23811, n23812,
         n23813, n23814, n23815, n23816, n23817, n23818, n23819, n23820,
         n23821, n23822, n23823, n23824, n23825, n23826, n23827, n23828,
         n23829, n23830, n23831, n23832, n23833, n23834, n23835, n23836,
         n23837, n23838, n23839, n23840, n23841, n23842, n23843, n23844,
         n23845, n23846, n23847, n23848, n23849, n23850, n23851, n23852,
         n23853, n23854, n23855, n23856, n23857, n23858, n23859, n23860,
         n23861, n23862, n23863, n23864, n23865, n23866, n23867, n23868,
         n23869, n23870, n23871, n23872, n23873, n23874, n23875, n23876,
         n23877, n23878, n23879, n23880, n23881, n23882, n23883, n23884,
         n23885, n23886, n23887, n23888, n23889, n23890, n23891, n23892,
         n23893, n23894, n23895, n23896, n23897, n23898, n23899, n23900,
         n23901, n23902, n23903, n23904, n23905, n23906, n23907, n23908,
         n23909, n23910, n23911, n23912, n23913, n23914, n23915, n23916,
         n23917, n23918, n23919, n23920, n23921, n23922, n23923, n23924,
         n23925, n23926, n23927, n23928, n23929, n23930, n23931, n23932,
         n23933, n23934, n23935, n23936, n23937, n23938, n23939, n23940,
         n23941, n23942, n23943, n23944, n23945, n23946, n23947, n23948,
         n23949, n23950, n23951, n23952, n23953, n23954, n23955, n23956,
         n23957, n23958, n23959, n23960, n23961, n23962, n23963, n23964,
         n23965, n23966, n23967, n23968, n23969, n23970, n23971, n23972,
         n23973, n23974, n23975, n23976, n23977, n23978, n23979, n23980,
         n23981, n23982, n23983, n23984, n23985, n23986, n23987, n23988,
         n23989, n23990, n23991, n23992, n23993, n23994, n23995, n23996,
         n23997, n23998, n23999, n24000, n24001, n24002, n24003, n24004,
         n24005, n24006, n24007, n24008, n24009, n24010, n24011, n24012,
         n24013, n24014, n24015, n24016, n24017, n24018, n24019, n24020,
         n24021, n24022, n24023, n24024, n24025, n24026, n24027, n24028,
         n24029, n24030, n24031, n24032, n24033, n24034, n24035, n24036,
         n24037, n24038, n24039, n24040, n24041, n24042, n24043, n24044,
         n24045, n24046, n24047, n24048, n24049, n24050, n24051, n24052,
         n24053, n24054, n24055, n24056, n24057, n24058, n24059, n24060,
         n24061, n24062, n24063, n24064, n24065, n24066, n24067, n24068,
         n24069, n24070, n24071, n24072, n24073, n24074, n24075, n24076,
         n24077, n24078, n24079, n24080, n24081, n24082, n24083, n24084,
         n24085, n24086, n24087, n24088, n24089, n24090, n24091, n24092,
         n24093, n24094, n24095, n24096, n24097, n24098, n24099, n24100,
         n24101, n24102, n24103, n24104, n24105, n24106, n24107, n24108,
         n24109, n24110, n24111, n24112, n24113, n24114, n24115, n24116,
         n24117, n24118, n24119, n24120, n24121, n24122, n24123, n24124,
         n24125, n24126, n24127, n24128, n24129, n24130, n24131, n24132,
         n24133, n24134, n24135, n24136, n24137, n24138, n24139, n24140,
         n24141, n24142, n24143, n24144, n24145, n24146, n24147, n24148,
         n24149, n24150, n24151, n24152, n24153, n24154, n24155, n24156,
         n24157, n24158, n24159, n24160, n24161, n24162, n24163, n24164,
         n24165, n24166, n24167, n24168, n24169, n24170, n24171, n24172,
         n24173, n24174, n24175, n24176, n24177, n24178, n24179, n24180,
         n24181, n24182, n24183, n24184, n24185, n24186, n24187, n24188,
         n24189, n24190, n24191, n24192, n24193, n24194, n24195, n24196,
         n24197, n24198, n24199, n24200, n24201, n24202, n24203, n24204,
         n24205, n24206, n24207, n24208, n24209, n24210, n24211, n24212,
         n24213, n24214, n24215, n24216, n24217, n24218, n24219, n24220,
         n24221, n24222, n24223, n24224, n24225, n24226, n24227, n24228,
         n24229, n24230, n24231, n24232, n24233, n24234, n24235, n24236,
         n24237, n24238, n24239, n24240, n24241, n24242, n24243, n24244,
         n24245, n24246, n24247, n24248, n24249, n24250, n24251, n24252,
         n24253, n24254, n24255, n24256, n24257, n24258, n24259, n24260,
         n24261, n24262, n24263, n24264, n24265, n24266, n24267, n24268,
         n24269, n24270, n24271, n24272, n24273, n24274, n24275, n24276,
         n24277, n24278, n24279, n24280, n24281, n24282, n24283, n24284,
         n24285, n24286, n24287, n24288, n24289, n24290, n24291, n24292,
         n24293, n24294, n24295, n24296, n24297, n24298, n24299, n24300,
         n24301, n24302, n24303, n24304, n24305, n24306, n24307, n24308,
         n24309, n24310, n24311, n24312, n24313, n24314, n24315, n24316,
         n24317, n24318, n24319, n24320, n24321, n24322, n24323, n24324,
         n24325, n24326, n24327, n24328, n24329, n24330, n24331, n24332,
         n24333, n24334, n24335, n24336, n24337, n24338, n24339, n24340,
         n24341, n24342, n24343, n24344, n24345, n24346, n24347, n24348,
         n24349, n24350, n24351, n24352, n24353, n24354, n24355, n24356,
         n24357, n24358, n24359, n24360, n24361, n24362, n24363, n24364,
         n24365, n24366, n24367, n24368, n24369, n24370, n24371, n24372,
         n24373, n24374, n24375, n24376, n24377, n24378, n24379, n24380,
         n24381, n24382, n24383, n24384, n24385, n24386, n24387, n24388,
         n24389, n24390, n24391, n24392, n24393, n24394, n24395, n24396,
         n24397, n24398, n24399, n24400, n24401, n24402, n24403, n24404,
         n24405, n24406, n24407, n24408, n24409, n24410, n24411, n24412,
         n24413, n24414, n24415, n24416, n24417, n24418, n24419, n24420,
         n24421, n24422, n24423, n24424, n24425, n24426, n24427, n24428,
         n24429, n24430, n24431, n24432, n24433, n24434, n24435, n24436,
         n24437, n24438, n24439, n24440, n24441, n24442, n24443, n24444,
         n24445, n24446, n24447, n24448, n24449, n24450, n24451, n24452,
         n24453, n24454, n24455, n24456, n24457, n24458, n24459, n24460,
         n24461, n24462, n24463, n24464, n24465, n24466, n24467, n24468,
         n24469, n24470, n24471, n24472, n24473, n24474, n24475, n24476,
         n24477, n24478, n24479, n24480, n24481, n24482, n24483, n24484,
         n24485, n24486, n24487, n24488, n24489, n24490, n24491, n24492,
         n24493, n24494, n24495, n24496, n24497, n24498, n24499, n24500,
         n24501, n24502, n24503, n24504, n24505, n24506, n24507, n24508,
         n24509, n24510, n24511, n24512, n24513, n24514, n24515, n24516,
         n24517, n24518, n24519, n24520, n24521, n24522, n24523, n24524,
         n24525, n24526, n24527, n24528, n24529, n24530, n24531, n24532,
         n24533, n24534, n24535, n24536, n24537, n24538, n24539, n24540,
         n24541, n24542, n24543, n24544, n24545, n24546, n24547, n24548,
         n24549, n24550, n24551, n24552, n24553, n24554, n24555, n24556,
         n24557, n24558, n24559, n24560, n24561, n24562, n24563, n24564,
         n24565, n24566, n24567, n24568, n24569, n24570, n24571, n24572,
         n24573, n24574, n24575, n24576, n24577, n24578, n24579, n24580,
         n24581, n24582, n24583, n24584, n24585, n24586, n24587, n24588,
         n24589, n24590, n24591, n24592, n24593, n24594, n24595, n24596,
         n24597, n24598, n24599, n24600, n24601, n24602, n24603, n24604,
         n24605, n24606, n24607, n24608, n24609, n24610, n24611, n24612,
         n24613, n24614, n24615, n24616, n24617, n24618, n24619, n24620,
         n24621, n24622, n24623, n24624, n24625, n24626, n24627, n24628,
         n24629, n24630, n24631, n24632, n24633, n24634, n24635, n24636,
         n24637, n24638, n24639, n24640, n24641, n24642, n24643, n24644,
         n24645, n24646, n24647, n24648, n24649, n24650, n24651, n24652,
         n24653, n24654, n24655, n24656, n24657, n24658, n24659, n24660,
         n24661, n24662, n24663, n24664, n24665, n24666, n24667, n24668,
         n24669, n24670, n24671, n24672, n24673, n24674, n24675, n24676,
         n24677, n24678, n24679, n24680, n24681, n24682, n24683, n24684,
         n24685, n24686, n24687, n24688, n24689, n24690, n24691, n24692,
         n24693, n24694, n24695, n24696, n24697, n24698, n24699, n24700,
         n24701, n24702, n24703, n24704, n24705, n24706, n24707, n24708,
         n24709, n24710, n24711, n24712, n24713, n24714, n24715, n24716,
         n24717, n24718, n24719, n24720, n24721, n24722, n24723, n24724,
         n24725, n24726, n24727, n24728, n24729, n24730, n24731, n24732,
         n24733, n24734, n24735, n24736, n24737, n24738, n24739, n24740,
         n24741, n24742, n24743, n24744, n24745, n24746, n24747, n24748,
         n24749, n24750, n24751, n24752, n24753, n24754, n24755, n24756,
         n24757, n24758, n24759, n24760, n24761, n24762, n24763, n24764,
         n24765, n24766, n24767, n24768, n24769, n24770, n24771, n24772,
         n24773, n24774, n24775, n24776, n24777, n24778, n24779, n24780,
         n24781, n24782, n24783, n24784, n24785, n24786, n24787, n24788,
         n24789, n24790, n24791, n24792, n24793, n24794, n24795, n24796,
         n24797, n24798, n24799, n24800, n24801, n24802, n24803, n24804,
         n24805, n24806, n24807, n24808, n24809, n24810, n24811, n24812,
         n24813, n24814, n24815, n24816, n24817, n24818, n24819, n24820,
         n24821, n24822, n24823, n24824, n24825, n24826, n24827, n24828,
         n24829, n24830, n24831, n24832, n24833, n24834, n24835, n24836,
         n24837, n24838, n24839, n24840, n24841, n24842, n24843, n24844,
         n24845, n24846, n24847, n24848, n24849, n24850, n24851, n24852,
         n24853, n24854, n24855, n24856, n24857, n24858, n24859, n24860,
         n24861, n24862, n24863, n24864, n24865, n24866, n24867, n24868,
         n24869, n24870, n24871, n24872, n24873, n24874, n24875, n24876,
         n24877, n24878, n24879, n24880, n24881, n24882, n24883, n24884,
         n24885, n24886, n24887, n24888, n24889, n24890, n24891, n24892,
         n24893, n24894, n24895, n24896, n24897, n24898, n24899, n24900,
         n24901, n24902, n24903, n24904, n24905, n24906, n24907, n24908,
         n24909, n24910, n24911, n24912, n24913, n24914, n24915, n24916,
         n24917, n24918, n24919, n24920, n24921, n24922, n24923, n24924,
         n24925, n24926, n24927, n24928, n24929, n24930, n24931, n24932,
         n24933, n24934, n24935, n24936, n24937, n24938, n24939, n24940,
         n24941, n24942, n24943, n24944, n24945, n24946, n24947, n24948,
         n24949, n24950, n24951, n24952, n24953, n24954, n24955, n24956,
         n24957, n24958, n24959, n24960, n24961, n24962, n24963, n24964,
         n24965, n24966, n24967, n24968, n24969, n24970, n24971, n24972,
         n24973, n24974, n24975, n24976, n24977, n24978, n24979, n24980,
         n24981, n24982, n24983, n24984, n24985, n24986, n24987, n24988,
         n24989, n24990, n24991, n24992, n24993, n24994, n24995, n24996,
         n24997, n24998, n24999, n25000, n25001, n25002, n25003, n25004,
         n25005, n25006, n25007, n25008, n25009, n25010, n25011, n25012,
         n25013, n25014, n25015, n25016, n25017, n25018, n25019, n25020,
         n25021, n25022, n25023, n25024, n25025, n25026, n25027, n25028,
         n25029, n25030, n25031, n25032, n25033, n25034, n25035, n25036,
         n25037, n25038, n25039, n25040, n25041, n25042, n25043, n25044,
         n25045, n25046, n25047, n25048, n25049, n25050, n25051, n25052,
         n25053, n25054, n25055, n25056, n25057, n25058, n25059, n25060,
         n25061, n25062, n25063, n25064, n25065, n25066, n25067, n25068,
         n25069, n25070, n25071, n25072, n25073, n25074, n25075, n25076,
         n25077, n25078, n25079, n25080, n25081, n25082, n25083, n25084,
         n25085, n25086, n25087, n25088, n25089, n25090, n25091, n25092,
         n25093, n25094, n25095, n25096, n25097, n25098, n25099, n25100,
         n25101, n25102, n25103, n25104, n25105, n25106, n25107, n25108,
         n25109, n25110, n25111, n25112, n25113, n25114, n25115, n25116,
         n25117, n25118, n25119, n25120, n25121, n25122, n25123, n25124,
         n25125, n25126, n25127, n25128, n25129, n25130, n25131, n25132,
         n25133, n25134, n25135, n25136, n25137, n25138, n25139, n25140,
         n25141, n25142, n25143, n25144, n25145, n25146, n25147, n25148,
         n25149, n25150, n25151, n25152, n25153, n25154, n25155, n25156,
         n25157, n25158, n25159, n25160, n25161, n25162, n25163, n25164,
         n25165, n25166, n25167, n25168, n25169, n25170, n25171, n25172,
         n25173, n25174, n25175, n25176, n25177, n25178, n25179, n25180,
         n25181, n25182, n25183, n25184, n25185, n25186, n25187, n25188,
         n25189, n25190, n25191, n25192, n25193, n25194, n25195, n25196,
         n25197, n25198, n25199, n25200, n25201, n25202, n25203, n25204,
         n25205, n25206, n25207, n25208, n25209, n25210, n25211, n25212,
         n25213, n25214, n25215, n25216, n25217, n25218, n25219, n25220,
         n25221, n25222, n25223, n25224, n25225, n25226, n25227, n25228,
         n25229, n25230, n25231, n25232, n25233, n25234, n25235, n25236,
         n25237, n25238, n25239, n25240, n25241, n25242, n25243, n25244,
         n25245, n25246, n25247, n25248, n25249, n25250, n25251, n25252,
         n25253, n25254, n25255, n25256, n25257, n25258, n25259, n25260,
         n25261, n25262, n25263, n25264, n25265, n25266, n25267, n25268,
         n25269, n25270, n25271, n25272, n25273, n25274, n25275, n25276,
         n25277, n25278, n25279, n25280, n25281, n25282, n25283, n25284,
         n25285, n25286, n25287, n25288, n25289, n25290, n25291, n25292,
         n25293, n25294, n25295, n25296, n25297, n25298, n25299, n25300,
         n25301, n25302, n25303, n25304, n25305, n25306, n25307, n25308,
         n25309, n25310, n25311, n25312, n25313, n25314, n25315, n25316,
         n25317, n25318, n25319, n25320, n25321, n25322, n25323, n25324,
         n25325, n25326, n25327, n25328, n25329, n25330, n25331, n25332,
         n25333, n25334, n25335, n25336, n25337, n25338, n25339, n25340,
         n25341, n25342, n25343, n25344, n25345, n25346, n25347, n25348,
         n25349, n25350, n25351, n25352, n25353, n25354, n25355, n25356,
         n25357, n25358, n25359, n25360, n25361, n25362, n25363, n25364,
         n25365, n25366, n25367, n25368, n25369, n25370, n25371, n25372,
         n25373, n25374, n25375, n25376, n25377, n25378, n25379, n25380,
         n25381, n25382, n25383, n25384, n25385, n25386, n25387, n25388,
         n25389, n25390, n25391, n25392, n25393, n25394, n25395, n25396,
         n25397, n25398, n25399, n25400, n25401, n25402, n25403, n25404,
         n25405, n25406, n25407, n25408, n25409, n25410, n25411, n25412,
         n25413, n25414, n25415, n25416, n25417, n25418, n25419, n25420,
         n25421, n25422, n25423, n25424, n25425, n25426, n25427, n25428,
         n25429, n25430, n25431, n25432, n25433, n25434, n25435, n25436,
         n25437, n25438, n25439, n25440, n25441, n25442, n25443, n25444,
         n25445, n25446, n25447, n25448, n25449, n25450, n25451, n25452,
         n25453, n25454, n25455, n25456, n25457, n25458, n25459, n25460,
         n25461, n25462, n25463, n25464, n25465, n25466, n25467, n25468,
         n25469, n25470, n25471, n25472, n25473, n25474, n25475, n25476,
         n25477, n25478, n25479, n25480, n25481, n25482, n25483, n25484,
         n25485, n25486, n25487, n25488, n25489, n25490, n25491, n25492,
         n25493, n25494, n25495, n25496, n25497, n25498, n25499, n25500,
         n25501, n25502, n25503, n25504, n25505, n25506, n25507, n25508,
         n25509, n25510, n25511, n25512, n25513, n25514, n25515, n25516,
         n25517, n25518, n25519, n25520, n25521, n25522, n25523, n25524,
         n25525, n25526, n25527, n25528, n25529, n25530, n25531, n25532,
         n25533, n25534, n25535, n25536, n25537, n25538, n25539, n25540,
         n25541, n25542, n25543, n25544, n25545, n25546, n25547, n25548,
         n25549, n25550, n25551, n25552, n25553, n25554, n25555, n25556,
         n25557, n25558, n25559, n25560, n25561, n25562, n25563, n25564,
         n25565, n25566, n25567, n25568, n25569, n25570, n25571, n25572,
         n25573, n25574, n25575, n25576, n25577, n25578, n25579, n25580,
         n25581, n25582, n25583, n25584, n25585, n25586, n25587, n25588,
         n25589, n25590, n25591, n25592, n25593, n25594, n25595, n25596,
         n25597, n25598, n25599, n25600, n25601, n25602, n25603, n25604,
         n25605, n25606, n25607, n25608, n25609, n25610, n25611, n25612,
         n25613, n25614, n25615, n25616, n25617, n25618, n25619, n25620,
         n25621, n25622, n25623, n25624, n25625, n25626, n25627, n25628,
         n25629, n25630, n25631, n25632, n25633, n25634, n25635, n25636,
         n25637, n25638, n25639, n25640, n25641, n25642, n25643, n25644,
         n25645, n25646, n25647, n25648, n25649, n25650, n25651, n25652,
         n25653, n25654, n25655, n25656, n25657, n25658, n25659, n25660,
         n25661, n25662, n25663, n25664, n25665, n25666, n25667, n25668,
         n25669, n25670, n25671, n25672, n25673, n25674, n25675, n25676,
         n25677, n25678, n25679, n25680, n25681, n25682, n25683, n25684,
         n25685, n25686, n25687, n25688, n25689, n25690, n25691, n25692,
         n25693, n25694, n25695, n25696, n25697, n25698, n25699, n25700,
         n25701, n25702, n25703, n25704, n25705, n25706, n25707, n25708,
         n25709, n25710, n25711, n25712, n25713, n25714, n25715, n25716,
         n25717, n25718, n25719, n25720, n25721, n25722, n25723, n25724,
         n25725, n25726, n25727, n25728, n25729, n25730, n25731, n25732,
         n25733, n25734, n25735, n25736, n25737, n25738, n25739, n25740,
         n25741, n25742, n25743, n25744, n25745, n25746, n25747, n25748,
         n25749, n25750, n25751, n25752, n25753, n25754, n25755, n25756,
         n25757, n25758, n25759, n25760, n25761, n25762, n25763, n25764,
         n25765, n25766, n25767, n25768, n25769, n25770, n25771, n25772,
         n25773, n25774, n25775, n25776, n25777, n25778, n25779, n25780,
         n25781, n25782, n25783, n25784, n25785, n25786, n25787, n25788,
         n25789, n25790, n25791, n25792, n25793, n25794, n25795, n25796,
         n25797, n25798, n25799, n25800, n25801, n25802, n25803, n25804,
         n25805, n25806, n25807, n25808, n25809, n25810, n25811, n25812,
         n25813, n25814, n25815, n25816, n25817, n25818, n25819, n25820,
         n25821, n25822, n25823, n25824, n25825, n25826, n25827, n25828,
         n25829, n25830, n25831, n25832, n25833, n25834, n25835, n25836,
         n25837, n25838, n25839, n25840, n25841, n25842, n25843, n25844,
         n25845, n25846, n25847, n25848, n25849, n25850, n25851, n25852,
         n25853, n25854, n25855, n25856, n25857, n25858, n25859, n25860,
         n25861, n25862, n25863, n25864, n25865, n25866, n25867, n25868,
         n25869, n25870, n25871, n25872, n25873, n25874, n25875, n25876,
         n25877, n25878, n25879, n25880, n25881, n25882, n25883, n25884,
         n25885, n25886, n25887, n25888, n25889, n25890, n25891, n25892,
         n25893, n25894, n25895, n25896, n25897, n25898, n25899, n25900,
         n25901, n25902, n25903, n25904, n25905, n25906, n25907, n25908,
         n25909, n25910, n25911, n25912, n25913, n25914, n25915, n25916,
         n25917, n25918, n25919, n25920, n25921, n25922, n25923, n25924,
         n25925, n25926, n25927, n25928, n25929, n25930, n25931, n25932,
         n25933, n25934, n25935, n25936, n25937, n25938, n25939, n25940,
         n25941, n25942, n25943, n25944, n25945, n25946, n25947, n25948,
         n25949, n25950, n25951, n25952, n25953, n25954, n25955, n25956,
         n25957, n25958, n25959, n25960, n25961, n25962, n25963, n25964,
         n25965, n25966, n25967, n25968, n25969, n25970, n25971, n25972,
         n25973, n25974, n25975, n25976, n25977, n25978, n25979, n25980,
         n25981, n25982, n25983, n25984, n25985, n25986, n25987, n25988,
         n25989, n25990, n25991, n25992, n25993, n25994, n25995, n25996,
         n25997, n25998, n25999, n26000, n26001, n26002, n26003, n26004,
         n26005, n26006, n26007, n26008, n26009, n26010, n26011, n26012,
         n26013, n26014, n26015, n26016, n26017, n26018, n26019, n26020,
         n26021, n26022, n26023, n26024, n26025, n26026, n26027, n26028,
         n26029, n26030, n26031, n26032, n26033, n26034, n26035, n26036,
         n26037, n26038, n26039, n26040, n26041, n26042, n26043, n26044,
         n26045, n26046, n26047, n26048, n26049, n26050, n26051, n26052,
         n26053, n26054, n26055, n26056, n26057, n26058, n26059, n26060,
         n26061, n26062, n26063, n26064, n26065, n26066, n26067, n26068,
         n26069, n26070, n26071, n26072, n26073, n26074, n26075, n26076,
         n26077, n26078, n26079, n26080, n26081, n26082, n26083, n26084,
         n26085, n26086, n26087, n26088, n26089, n26090, n26091, n26092,
         n26093, n26094, n26095, n26096, n26097, n26098, n26099, n26100,
         n26101, n26102, n26103, n26104, n26105, n26106, n26107, n26108,
         n26109, n26110, n26111, n26112, n26113, n26114, n26115, n26116,
         n26117, n26118, n26119, n26120, n26121, n26122, n26123, n26124,
         n26125, n26126, n26127, n26128, n26129, n26130, n26131, n26132,
         n26133, n26134, n26135, n26136, n26137, n26138, n26139, n26140,
         n26141, n26142, n26143, n26144, n26145, n26146, n26147, n26148,
         n26149, n26150, n26151, n26152, n26153, n26154, n26155, n26156,
         n26157, n26158, n26159, n26160, n26161, n26162, n26163, n26164,
         n26165, n26166, n26167, n26168, n26169, n26170, n26171, n26172,
         n26173, n26174, n26175, n26176, n26177, n26178, n26179, n26180,
         n26181, n26182, n26183, n26184, n26185, n26186, n26187, n26188,
         n26189, n26190, n26191, n26192, n26193, n26194, n26195, n26196,
         n26197, n26198, n26199, n26200, n26201, n26202, n26203, n26204,
         n26205, n26206, n26207, n26208, n26209, n26210, n26211, n26212,
         n26213, n26214, n26215, n26216, n26217, n26218, n26219, n26220,
         n26221, n26222, n26223, n26224, n26225, n26226, n26227, n26228,
         n26229, n26230, n26231, n26232, n26233, n26234, n26235, n26236,
         n26237, n26238, n26239, n26240, n26241, n26242, n26243, n26244,
         n26245, n26246, n26247, n26248, n26249, n26250, n26251, n26252,
         n26253, n26254, n26255, n26256, n26257, n26258, n26259, n26260,
         n26261, n26262, n26263, n26264, n26265, n26266, n26267, n26268,
         n26269, n26270, n26271, n26272, n26273, n26274, n26275, n26276,
         n26277, n26278, n26279, n26280, n26281, n26282, n26283, n26284,
         n26285, n26286, n26287, n26288, n26289, n26290, n26291, n26292,
         n26293, n26294, n26295, n26296, n26297, n26298, n26299, n26300,
         n26301, n26302, n26303, n26304, n26305, n26306, n26307, n26308,
         n26309, n26310, n26311, n26312, n26313, n26314, n26315, n26316,
         n26317, n26318, n26319, n26320, n26321, n26322, n26323, n26324,
         n26325, n26326, n26327, n26328, n26329, n26330, n26331, n26332,
         n26333, n26334, n26335, n26336, n26337, n26338, n26339, n26340,
         n26341, n26342, n26343, n26344, n26345, n26346, n26347, n26348,
         n26349, n26350, n26351, n26352, n26353, n26354, n26355, n26356,
         n26357, n26358, n26359, n26360, n26361, n26362, n26363, n26364,
         n26365, n26366, n26367, n26368, n26369, n26370, n26371, n26372,
         n26373, n26374, n26375, n26376, n26377, n26378, n26379, n26380,
         n26381, n26382, n26383, n26384, n26385, n26386, n26387, n26388,
         n26389, n26390, n26391, n26392, n26393, n26394, n26395, n26396,
         n26397, n26398, n26399, n26400, n26401, n26402, n26403, n26404,
         n26405, n26406, n26407, n26408, n26409, n26410, n26411, n26412,
         n26413, n26414, n26415, n26416, n26417, n26418, n26419, n26420,
         n26421, n26422, n26423, n26424, n26425, n26426, n26427, n26428,
         n26429, n26430, n26431, n26432, n26433, n26434, n26435, n26436,
         n26437, n26438, n26439, n26440, n26441, n26442, n26443, n26444,
         n26445, n26446, n26447, n26448, n26449, n26450, n26451, n26452,
         n26453, n26454, n26455, n26456, n26457, n26458, n26459, n26460,
         n26461, n26462, n26463, n26464, n26465, n26466, n26467, n26468,
         n26469, n26470, n26471, n26472, n26473, n26474, n26475, n26476,
         n26477, n26478, n26479, n26480, n26481, n26482, n26483, n26484,
         n26485, n26486, n26487, n26488, n26489, n26490, n26491, n26492,
         n26493, n26494, n26495, n26496, n26497, n26498, n26499, n26500,
         n26501, n26502, n26503, n26504, n26505, n26506, n26507, n26508,
         n26509, n26510, n26511, n26512, n26513, n26514, n26515, n26516,
         n26517, n26518, n26519, n26520, n26521, n26522, n26523, n26524,
         n26525, n26526, n26527, n26528, n26529, n26530, n26531, n26532,
         n26533, n26534, n26535, n26536, n26537, n26538, n26539, n26540,
         n26541, n26542, n26543, n26544, n26545, n26546, n26547, n26548,
         n26549, n26550, n26551, n26552, n26553, n26554, n26555, n26556,
         n26557, n26558, n26559, n26560, n26561, n26562, n26563, n26564,
         n26565, n26566, n26567, n26568, n26569, n26570, n26571, n26572,
         n26573, n26574, n26575, n26576, n26577, n26578, n26579, n26580,
         n26581, n26582, n26583, n26584, n26585, n26586, n26587, n26588,
         n26589, n26590, n26591, n26592, n26593, n26594, n26595, n26596,
         n26597, n26598, n26599, n26600, n26601, n26602, n26603, n26604,
         n26605, n26606, n26607, n26608, n26609, n26610, n26611, n26612,
         n26613, n26614, n26615, n26616, n26617, n26618, n26619, n26620,
         n26621, n26622, n26623, n26624, n26625, n26626, n26627, n26628,
         n26629, n26630, n26631, n26632, n26633, n26634, n26635, n26636,
         n26637, n26638, n26639, n26640, n26641, n26642, n26643, n26644,
         n26645, n26646, n26647, n26648, n26649, n26650, n26651, n26652,
         n26653, n26654, n26655, n26656, n26657, n26658, n26659, n26660,
         n26661, n26662, n26663, n26664, n26665, n26666, n26667, n26668,
         n26669, n26670, n26671, n26672, n26673, n26674, n26675, n26676,
         n26677, n26678, n26679, n26680, n26681, n26682, n26683, n26684,
         n26685, n26686, n26687, n26688, n26689, n26690, n26691, n26692,
         n26693, n26694, n26695, n26696, n26697, n26698, n26699, n26700,
         n26701, n26702, n26703, n26704, n26705, n26706, n26707, n26708,
         n26709, n26710, n26711, n26712, n26713, n26714, n26715, n26716,
         n26717, n26718, n26719, n26720, n26721, n26722, n26723, n26724,
         n26725, n26726, n26727, n26728, n26729, n26730, n26731, n26732,
         n26733, n26734, n26735, n26736, n26737, n26738, n26739, n26740,
         n26741, n26742, n26743, n26744, n26745, n26746, n26747, n26748,
         n26749, n26750, n26751, n26752, n26753, n26754, n26755, n26756,
         n26757, n26758, n26759, n26760, n26761, n26762, n26763, n26764,
         n26765, n26766, n26767, n26768, n26769, n26770, n26771, n26772,
         n26773, n26774, n26775, n26776, n26777, n26778, n26779, n26780,
         n26781, n26782, n26783, n26784, n26785, n26786, n26787, n26788,
         n26789, n26790, n26791, n26792, n26793, n26794, n26795, n26796,
         n26797, n26798, n26799, n26800, n26801, n26802, n26803, n26804,
         n26805, n26806, n26807, n26808, n26809, n26810, n26811, n26812,
         n26813, n26814, n26815, n26816, n26817, n26818, n26819, n26820,
         n26821, n26822, n26823, n26824, n26825, n26826, n26827, n26828,
         n26829, n26830, n26831, n26832, n26833, n26834, n26835, n26836,
         n26837, n26838, n26839, n26840, n26841, n26842, n26843, n26844,
         n26845, n26846, n26847, n26848, n26849, n26850, n26851, n26852,
         n26853, n26854, n26855, n26856, n26857, n26858, n26859, n26860,
         n26861, n26862, n26863, n26864, n26865, n26866, n26867, n26868,
         n26869, n26870, n26871, n26872, n26873, n26874, n26875, n26876,
         n26877, n26878, n26879, n26880, n26881, n26882, n26883, n26884,
         n26885, n26886, n26887, n26888, n26889, n26890, n26891, n26892,
         n26893, n26894, n26895, n26896, n26897, n26898, n26899, n26900,
         n26901, n26902, n26903, n26904, n26905, n26906, n26907, n26908,
         n26909, n26910, n26911, n26912, n26913, n26914, n26915, n26916,
         n26917, n26918, n26919, n26920, n26921, n26922, n26923, n26924,
         n26925, n26926, n26927, n26928, n26929, n26930, n26931, n26932,
         n26933, n26934, n26935, n26936, n26937, n26938, n26939, n26940,
         n26941, n26942, n26943, n26944, n26945, n26946, n26947, n26948,
         n26949, n26950, n26951, n26952, n26953, n26954, n26955, n26956,
         n26957, n26958, n26959, n26960, n26961, n26962, n26963, n26964,
         n26965, n26966, n26967, n26968, n26969, n26970, n26971, n26972,
         n26973, n26974, n26975, n26976, n26977, n26978, n26979, n26980,
         n26981, n26982, n26983, n26984, n26985, n26986, n26987, n26988,
         n26989, n26990, n26991, n26992, n26993, n26994, n26995, n26996,
         n26997, n26998, n26999, n27000, n27001, n27002, n27003, n27004,
         n27005, n27006, n27007, n27008, n27009, n27010, n27011, n27012,
         n27013, n27014, n27015, n27016, n27017, n27018, n27019, n27020,
         n27021, n27022, n27023, n27024, n27025, n27026, n27027, n27028,
         n27029, n27030, n27031, n27032, n27033, n27034, n27035, n27036,
         n27037, n27038, n27039, n27040, n27041, n27042, n27043, n27044,
         n27045, n27046, n27047, n27048, n27049, n27050, n27051, n27052,
         n27053, n27054, n27055, n27056, n27057, n27058, n27059, n27060,
         n27061, n27062, n27063, n27064, n27065, n27066, n27067, n27068,
         n27069, n27070, n27071, n27072, n27073, n27074, n27075, n27076,
         n27077, n27078, n27079, n27080, n27081, n27082, n27083, n27084,
         n27085, n27086, n27087, n27088, n27089, n27090, n27091, n27092,
         n27093, n27094, n27095, n27096, n27097, n27098, n27099, n27100,
         n27101, n27102, n27103, n27104, n27105, n27106, n27107, n27108,
         n27109, n27110, n27111, n27112, n27113, n27114, n27115, n27116,
         n27117, n27118, n27119, n27120, n27121, n27122, n27123, n27124,
         n27125, n27126, n27127, n27128, n27129, n27130, n27131, n27132,
         n27133, n27134, n27135, n27136, n27137, n27138, n27139, n27140,
         n27141, n27142, n27143, n27144, n27145, n27146, n27147, n27148,
         n27149, n27150, n27151, n27152, n27153, n27154, n27155, n27156,
         n27157, n27158, n27159, n27160, n27161, n27162, n27163, n27164,
         n27165, n27166, n27167, n27168, n27169, n27170, n27171, n27172,
         n27173, n27174, n27175, n27176, n27177, n27178, n27179, n27180,
         n27181, n27182, n27183, n27184, n27185, n27186, n27187, n27188,
         n27189, n27190, n27191, n27192, n27193, n27194, n27195, n27196,
         n27197, n27198, n27199, n27200, n27201, n27202, n27203, n27204,
         n27205, n27206, n27207, n27208, n27209, n27210, n27211, n27212,
         n27213, n27214, n27215, n27216, n27217, n27218, n27219, n27220,
         n27221, n27222, n27223, n27224, n27225, n27226, n27227, n27228,
         n27229, n27230, n27231, n27232, n27233, n27234, n27235, n27236,
         n27237, n27238, n27239, n27240, n27241, n27242, n27243, n27244,
         n27245, n27246, n27247, n27248, n27249, n27250, n27251, n27252,
         n27253, n27254, n27255, n27256, n27257, n27258, n27259, n27260,
         n27261, n27262, n27263, n27264, n27265, n27266, n27267, n27268,
         n27269, n27270, n27271, n27272, n27273, n27274, n27275, n27276,
         n27277, n27278, n27279, n27280, n27281, n27282, n27283, n27284,
         n27285, n27286, n27287, n27288, n27289, n27290, n27291, n27292,
         n27293, n27294, n27295, n27296, n27297, n27298, n27299, n27300,
         n27301, n27302, n27303, n27304, n27305, n27306, n27307, n27308,
         n27309, n27310, n27311, n27312, n27313, n27314, n27315, n27316,
         n27317, n27318, n27319, n27320, n27321, n27322, n27323, n27324,
         n27325, n27326, n27327, n27328, n27329, n27330, n27331, n27332,
         n27333, n27334, n27335, n27336, n27337, n27338, n27339, n27340,
         n27341, n27342, n27343, n27344, n27345, n27346, n27347, n27348,
         n27349, n27350, n27351, n27352, n27353, n27354, n27355, n27356,
         n27357, n27358, n27359, n27360, n27361, n27362, n27363, n27364,
         n27365, n27366, n27367, n27368, n27369, n27370, n27371, n27372,
         n27373, n27374, n27375, n27376, n27377, n27378, n27379, n27380,
         n27381, n27382, n27383, n27384, n27385, n27386, n27387, n27388,
         n27389, n27390, n27391, n27392, n27393, n27394, n27395, n27396,
         n27397, n27398, n27399, n27400, n27401, n27402, n27403, n27404,
         n27405, n27406, n27407, n27408, n27409, n27410, n27411, n27412,
         n27413, n27414, n27415, n27416, n27417, n27418, n27419, n27420,
         n27421, n27422, n27423, n27424, n27425, n27426, n27427, n27428,
         n27429, n27430, n27431, n27432, n27433, n27434, n27435, n27436,
         n27437, n27438, n27439, n27440, n27441, n27442, n27443, n27444,
         n27445, n27446, n27447, n27448, n27449, n27450, n27451, n27452,
         n27453, n27454, n27455, n27456, n27457, n27458, n27459, n27460,
         n27461, n27462, n27463, n27464, n27465, n27466, n27467, n27468,
         n27469, n27470, n27471, n27472, n27473, n27474, n27475, n27476,
         n27477, n27478, n27479, n27480, n27481, n27482, n27483, n27484,
         n27485, n27486, n27487, n27488, n27489, n27490, n27491, n27492,
         n27493, n27494, n27495, n27496, n27497, n27498, n27499, n27500,
         n27501, n27502, n27503, n27504, n27505, n27506, n27507, n27508,
         n27509, n27510, n27511, n27512, n27513, n27514, n27515, n27516,
         n27517, n27518, n27519, n27520, n27521, n27522, n27523, n27524,
         n27525, n27526, n27527, n27528, n27529, n27530, n27531, n27532,
         n27533, n27534, n27535, n27536, n27537, n27538, n27539, n27540,
         n27541, n27542, n27543, n27544, n27545, n27546, n27547, n27548,
         n27549, n27550, n27551, n27552, n27553, n27554, n27555, n27556,
         n27557, n27558, n27559, n27560, n27561, n27562, n27563, n27564,
         n27565, n27566, n27567, n27568, n27569, n27570, n27571, n27572,
         n27573, n27574, n27575, n27576, n27577, n27578, n27579, n27580,
         n27581, n27582, n27583, n27584, n27585, n27586, n27587, n27588,
         n27589, n27590, n27591, n27592, n27593, n27594, n27595, n27596,
         n27597, n27598, n27599, n27600, n27601, n27602, n27603, n27604,
         n27605, n27606, n27607, n27608, n27609, n27610, n27611, n27612,
         n27613, n27614, n27615, n27616, n27617, n27618, n27619, n27620,
         n27621, n27622, n27623, n27624, n27625, n27626, n27627, n27628,
         n27629, n27630, n27631, n27632, n27633, n27634, n27635, n27636,
         n27637, n27638, n27639, n27640, n27641, n27642, n27643, n27644,
         n27645, n27646, n27647, n27648, n27649, n27650, n27651, n27652,
         n27653, n27654, n27655, n27656, n27657, n27658, n27659, n27660,
         n27661, n27662, n27663, n27664, n27665, n27666, n27667, n27668,
         n27669, n27670, n27671, n27672, n27673, n27674, n27675, n27676,
         n27677, n27678, n27679, n27680, n27681, n27682, n27683, n27684,
         n27685, n27686, n27687, n27688, n27689, n27690, n27691, n27692,
         n27693, n27694, n27695, n27696, n27697, n27698, n27699, n27700,
         n27701, n27702, n27703, n27704, n27705, n27706, n27707, n27708,
         n27709, n27710, n27711, n27712, n27713, n27714, n27715, n27716,
         n27717, n27718, n27719, n27720, n27721, n27722, n27723, n27724,
         n27725, n27726, n27727, n27728, n27729, n27730, n27731, n27732,
         n27733, n27734, n27735, n27736, n27737, n27738, n27739, n27740,
         n27741, n27742, n27743, n27744, n27745, n27746, n27747, n27748,
         n27749, n27750, n27751, n27752, n27753, n27754, n27755, n27756,
         n27757, n27758, n27759, n27760, n27761, n27762, n27763, n27764,
         n27765, n27766, n27767, n27768, n27769, n27770, n27771, n27772,
         n27773, n27774, n27775, n27776, n27777, n27778, n27779, n27780,
         n27781, n27782, n27783, n27784, n27785, n27786, n27787, n27788,
         n27789, n27790, n27791, n27792, n27793, n27794, n27795, n27796,
         n27797, n27798, n27799, n27800, n27801, n27802, n27803, n27804,
         n27805, n27806, n27807, n27808, n27809, n27810, n27811, n27812,
         n27813, n27814, n27815, n27816, n27817, n27818, n27819, n27820,
         n27821, n27822, n27823, n27824, n27825, n27826, n27827, n27828,
         n27829, n27830, n27831, n27832, n27833, n27834, n27835, n27836,
         n27837, n27838, n27839, n27840, n27841, n27842, n27843, n27844,
         n27845, n27846, n27847, n27848, n27849, n27850, n27851, n27852,
         n27853, n27854, n27855, n27856, n27857, n27858, n27859, n27860,
         n27861, n27862, n27863, n27864, n27865, n27866, n27867, n27868,
         n27869, n27870, n27871, n27872, n27873, n27874, n27875, n27876,
         n27877, n27878, n27879, n27880, n27881, n27882, n27883, n27884,
         n27885, n27886, n27887, n27888, n27889, n27890, n27891, n27892,
         n27893, n27894, n27895, n27896, n27897, n27898, n27899, n27900,
         n27901, n27902, n27903, n27904, n27905, n27906, n27907, n27908,
         n27909, n27910, n27911, n27912, n27913, n27914, n27915, n27916,
         n27917, n27918, n27919, n27920, n27921, n27922, n27923, n27924,
         n27925, n27926, n27927, n27928, n27929, n27930, n27931, n27932,
         n27933, n27934, n27935, n27936, n27937, n27938, n27939, n27940,
         n27941, n27942, n27943, n27944, n27945, n27946, n27947, n27948,
         n27949, n27950, n27951, n27952, n27953, n27954, n27955, n27956,
         n27957, n27958, n27959, n27960, n27961, n27962, n27963, n27964,
         n27965, n27966, n27967, n27968, n27969, n27970, n27971, n27972,
         n27973, n27974, n27975, n27976, n27977, n27978, n27979, n27980,
         n27981, n27982, n27983, n27984, n27985, n27986, n27987, n27988,
         n27989, n27990, n27991, n27992, n27993, n27994, n27995, n27996,
         n27997, n27998, n27999, n28000, n28001, n28002, n28003, n28004,
         n28005, n28006, n28007, n28008, n28009, n28010, n28011, n28012,
         n28013, n28014, n28015, n28016, n28017, n28018, n28019, n28020,
         n28021, n28022, n28023, n28024, n28025, n28026, n28027, n28028,
         n28029, n28030, n28031, n28032, n28033, n28034, n28035, n28036,
         n28037, n28038, n28039, n28040, n28041, n28042, n28043, n28044,
         n28045, n28046, n28047, n28048, n28049, n28050, n28051, n28052,
         n28053, n28054, n28055, n28056, n28057, n28058, n28059, n28060,
         n28061, n28062, n28063, n28064, n28065, n28066, n28067, n28068,
         n28069, n28070, n28071, n28072, n28073, n28074, n28075, n28076,
         n28077, n28078, n28079, n28080, n28081, n28082, n28083, n28084,
         n28085, n28086, n28087, n28088, n28089, n28090, n28091, n28092,
         n28093, n28094, n28095, n28096, n28097, n28098, n28099, n28100,
         n28101, n28102, n28103, n28104, n28105, n28106, n28107, n28108,
         n28109, n28110, n28111, n28112, n28113, n28114, n28115, n28116,
         n28117, n28118, n28119, n28120, n28121, n28122, n28123, n28124,
         n28125, n28126, n28127, n28128, n28129, n28130, n28131, n28132,
         n28133, n28134, n28135, n28136, n28137, n28138, n28139, n28140,
         n28141, n28142, n28143, n28144, n28145, n28146, n28147, n28148,
         n28149, n28150, n28151, n28152, n28153, n28154, n28155, n28156,
         n28157, n28158, n28159, n28160, n28161, n28162, n28163, n28164,
         n28165, n28166, n28167, n28168, n28169, n28170, n28171, n28172,
         n28173, n28174, n28175, n28176, n28177, n28178, n28179, n28180,
         n28181, n28182, n28183, n28184, n28185, n28186, n28187, n28188,
         n28189, n28190, n28191, n28192, n28193, n28194, n28195, n28196,
         n28197, n28198, n28199, n28200, n28201, n28202, n28203, n28204,
         n28205, n28206, n28207, n28208, n28209, n28210, n28211, n28212,
         n28213, n28214, n28215, n28216, n28217, n28218, n28219, n28220,
         n28221, n28222, n28223, n28224, n28225, n28226, n28227, n28228,
         n28229, n28230, n28231, n28232, n28233, n28234, n28235, n28236,
         n28237, n28238, n28239, n28240, n28241, n28242, n28243, n28244,
         n28245, n28246, n28247, n28248, n28249, n28250, n28251, n28252,
         n28253, n28254, n28255, n28256, n28257, n28258, n28259, n28260,
         n28261, n28262, n28263, n28264, n28265, n28266, n28267, n28268,
         n28269, n28270, n28271, n28272, n28273, n28274, n28275, n28276,
         n28277, n28278, n28279, n28280, n28281, n28282, n28283, n28284,
         n28285, n28286, n28287, n28288, n28289, n28290, n28291, n28292,
         n28293, n28294, n28295, n28296, n28297, n28298, n28299, n28300,
         n28301, n28302, n28303, n28304, n28305, n28306, n28307, n28308,
         n28309, n28310, n28311, n28312, n28313, n28314, n28315, n28316,
         n28317, n28318, n28319, n28320, n28321, n28322, n28323, n28324,
         n28325, n28326, n28327, n28328, n28329, n28330, n28331, n28332,
         n28333, n28334, n28335, n28336, n28337, n28338, n28339, n28340,
         n28341, n28342, n28343, n28344, n28345, n28346, n28347, n28348,
         n28349, n28350, n28351, n28352, n28353, n28354, n28355, n28356,
         n28357, n28358, n28359, n28360, n28361, n28362, n28363, n28364,
         n28365, n28366, n28367, n28368, n28369, n28370, n28371, n28372,
         n28373, n28374, n28375, n28376, n28377, n28378, n28379, n28380,
         n28381, n28382, n28383, n28384, n28385, n28386, n28387, n28388,
         n28389, n28390, n28391, n28392, n28393, n28394, n28395, n28396,
         n28397, n28398, n28399, n28400, n28401, n28402, n28403, n28404,
         n28405, n28406, n28407, n28408, n28409, n28410, n28411, n28412,
         n28413, n28414, n28415, n28416, n28417, n28418, n28419, n28420,
         n28421, n28422, n28423, n28424, n28425, n28426, n28427, n28428,
         n28429, n28430, n28431, n28432, n28433, n28434, n28435, n28436,
         n28437, n28438, n28439, n28440, n28441, n28442, n28443, n28444,
         n28445, n28446, n28447, n28448, n28449, n28450, n28451, n28452,
         n28453, n28454, n28455, n28456, n28457, n28458, n28459, n28460,
         n28461, n28462, n28463, n28464, n28465, n28466, n28467, n28468,
         n28469, n28470, n28471, n28472, n28473, n28474, n28475, n28476,
         n28477, n28478, n28479, n28480, n28481, n28482, n28483, n28484,
         n28485, n28486, n28487, n28488, n28489, n28490, n28491, n28492,
         n28493, n28494, n28495, n28496, n28497, n28498, n28499, n28500,
         n28501, n28502, n28503, n28504, n28505, n28506, n28507, n28508,
         n28509, n28510, n28511, n28512, n28513, n28514, n28515, n28516,
         n28517, n28518, n28519, n28520, n28521, n28522, n28523, n28524,
         n28525, n28526, n28527, n28528, n28529, n28530, n28531, n28532,
         n28533, n28534, n28535, n28536, n28537, n28538, n28539, n28540,
         n28541, n28542, n28543, n28544, n28545, n28546, n28547, n28548,
         n28549, n28550, n28551, n28552, n28553, n28554, n28555, n28556,
         n28557, n28558, n28559, n28560, n28561, n28562, n28563, n28564,
         n28565, n28566, n28567, n28568, n28569, n28570, n28571, n28572,
         n28573, n28574, n28575, n28576, n28577, n28578, n28579, n28580,
         n28581, n28582, n28583, n28584, n28585, n28586, n28587, n28588,
         n28589, n28590, n28591, n28592, n28593, n28594, n28595, n28596,
         n28597, n28598, n28599, n28600, n28601, n28602, n28603, n28604,
         n28605, n28606, n28607, n28608, n28609, n28610, n28611, n28612,
         n28613, n28614, n28615, n28616, n28617, n28618, n28619, n28620,
         n28621, n28622, n28623, n28624, n28625, n28626, n28627, n28628,
         n28629, n28630, n28631, n28632, n28633, n28634, n28635, n28636,
         n28637, n28638, n28639, n28640, n28641, n28642, n28643, n28644,
         n28645, n28646, n28647, n28648, n28649, n28650, n28651, n28652,
         n28653, n28654, n28655, n28656, n28657, n28658, n28659, n28660,
         n28661, n28662, n28663, n28664, n28665, n28666, n28667, n28668,
         n28669, n28670, n28671, n28672, n28673, n28674, n28675, n28676,
         n28677, n28678, n28679, n28680, n28681, n28682, n28683, n28684,
         n28685, n28686, n28687, n28688, n28689, n28690, n28691, n28692,
         n28693, n28694, n28695, n28696, n28697, n28698, n28699, n28700,
         n28701, n28702, n28703, n28704, n28705, n28706, n28707, n28708,
         n28709, n28710, n28711, n28712, n28713, n28714, n28715, n28716,
         n28717, n28718, n28719, n28720, n28721, n28722, n28723, n28724,
         n28725, n28726, n28727, n28728, n28729, n28730, n28731, n28732,
         n28733, n28734, n28735, n28736, n28737, n28738, n28739, n28740,
         n28741, n28742, n28743, n28744, n28745, n28746, n28747, n28748,
         n28749, n28750, n28751, n28752, n28753, n28754, n28755, n28756,
         n28757, n28758, n28759, n28760, n28761, n28762, n28763, n28764,
         n28765, n28766, n28767, n28768, n28769, n28770, n28771, n28772,
         n28773, n28774, n28775, n28776, n28777, n28778, n28779, n28780,
         n28781, n28782, n28783, n28784, n28785, n28786, n28787, n28788,
         n28789, n28790, n28791, n28792, n28793, n28794, n28795, n28796,
         n28797, n28798, n28799, n28800, n28801, n28802, n28803, n28804,
         n28805, n28806, n28807, n28808, n28809, n28810, n28811, n28812,
         n28813, n28814, n28815, n28816, n28817, n28818, n28819, n28820,
         n28821, n28822, n28823, n28824, n28825, n28826, n28827, n28828,
         n28829, n28830, n28831, n28832, n28833, n28834, n28835, n28836,
         n28837, n28838, n28839, n28840, n28841, n28842, n28843, n28844,
         n28845, n28846, n28847, n28848, n28849, n28850, n28851, n28852,
         n28853, n28854, n28855, n28856, n28857, n28858, n28859, n28860,
         n28861, n28862, n28863, n28864, n28865, n28866, n28867, n28868,
         n28869, n28870, n28871, n28872, n28873, n28874, n28875, n28876,
         n28877, n28878, n28879, n28880, n28881, n28882, n28883, n28884,
         n28885, n28886, n28887, n28888, n28889, n28890, n28891, n28892,
         n28893, n28894, n28895, n28896, n28897, n28898, n28899, n28900,
         n28901, n28902, n28903, n28904, n28905, n28906, n28907, n28908,
         n28909, n28910, n28911, n28912, n28913, n28914, n28915, n28916,
         n28917, n28918, n28919, n28920, n28921, n28922, n28923, n28924,
         n28925, n28926, n28927, n28928, n28929, n28930, n28931, n28932,
         n28933, n28934, n28935, n28936, n28937, n28938, n28939, n28940,
         n28941, n28942, n28943, n28944, n28945, n28946, n28947, n28948,
         n28949, n28950, n28951, n28952, n28953, n28954, n28955, n28956,
         n28957, n28958, n28959, n28960, n28961, n28962, n28963, n28964,
         n28965, n28966, n28967, n28968, n28969, n28970, n28971, n28972,
         n28973, n28974, n28975, n28976, n28977, n28978, n28979, n28980,
         n28981, n28982, n28983, n28984, n28985, n28986, n28987, n28988,
         n28989, n28990, n28991, n28992, n28993, n28994, n28995, n28996,
         n28997, n28998, n28999, n29000, n29001, n29002, n29003, n29004,
         n29005, n29006, n29007, n29008, n29009, n29010, n29011, n29012,
         n29013, n29014, n29015, n29016, n29017, n29018, n29019, n29020,
         n29021, n29022, n29023, n29024, n29025, n29026, n29027, n29028,
         n29029, n29030, n29031, n29032, n29033, n29034, n29035, n29036,
         n29037, n29038, n29039, n29040, n29041, n29042, n29043, n29044,
         n29045, n29046, n29047, n29048, n29049, n29050, n29051, n29052,
         n29053, n29054, n29055, n29056, n29057, n29058, n29059, n29060,
         n29061, n29062, n29063, n29064, n29065, n29066, n29067, n29068,
         n29069, n29070, n29071, n29072, n29073, n29074, n29075, n29076,
         n29077, n29078, n29079, n29080, n29081, n29082, n29083, n29084,
         n29085, n29086, n29087, n29088, n29089, n29090, n29091, n29092,
         n29093, n29094, n29095, n29096, n29097, n29098, n29099, n29100,
         n29101, n29102, n29103, n29104, n29105, n29106, n29107, n29108,
         n29109, n29110, n29111, n29112, n29113, n29114, n29115, n29116,
         n29117, n29118, n29119, n29120, n29121, n29122, n29123, n29124,
         n29125, n29126, n29127, n29128, n29129, n29130, n29131, n29132,
         n29133, n29134, n29135, n29136, n29137, n29138, n29139, n29140,
         n29141, n29142, n29143, n29144, n29145, n29146, n29147, n29148,
         n29149, n29150, n29151, n29152, n29153, n29154, n29155, n29156,
         n29157, n29158, n29159, n29160, n29161, n29162, n29163, n29164,
         n29165, n29166, n29167, n29168, n29169, n29170, n29171, n29172,
         n29173, n29174, n29175, n29176, n29177, n29178, n29179, n29180,
         n29181, n29182, n29183, n29184, n29185, n29186, n29187, n29188,
         n29189, n29190, n29191, n29192, n29193, n29194, n29195, n29196,
         n29197, n29198, n29199, n29200, n29201, n29202, n29203, n29204,
         n29205, n29206, n29207, n29208, n29209, n29210, n29211, n29212,
         n29213, n29214, n29215, n29216, n29217, n29218, n29219, n29220,
         n29221, n29222, n29223, n29224, n29225, n29226, n29227, n29228,
         n29229, n29230, n29231, n29232, n29233, n29234, n29235, n29236,
         n29237, n29238, n29239, n29240, n29241, n29242, n29243, n29244,
         n29245, n29246, n29247, n29248, n29249, n29250, n29251, n29252,
         n29253, n29254, n29255, n29256, n29257, n29258, n29259, n29260,
         n29261, n29262, n29263, n29264, n29265, n29266, n29267, n29268,
         n29269, n29270, n29271, n29272, n29273, n29274, n29275, n29276,
         n29277, n29278, n29279, n29280, n29281, n29282, n29283, n29284,
         n29285, n29286, n29287, n29288, n29289, n29290, n29291, n29292,
         n29293, n29294, n29295, n29296, n29297, n29298, n29299, n29300,
         n29301, n29302, n29303, n29304, n29305, n29306, n29307, n29308,
         n29309, n29310, n29311, n29312, n29313, n29314, n29315, n29316,
         n29317, n29318, n29319, n29320, n29321, n29322, n29323, n29324,
         n29325, n29326, n29327, n29328, n29329, n29330, n29331, n29332,
         n29333, n29334, n29335, n29336, n29337, n29338, n29339, n29340,
         n29341, n29342, n29343, n29344, n29345, n29346, n29347, n29348,
         n29349, n29350, n29351, n29352, n29353, n29354, n29355, n29356,
         n29357, n29358, n29359, n29360, n29361, n29362, n29363, n29364,
         n29365, n29366, n29367, n29368, n29369, n29370, n29371, n29372,
         n29373, n29374, n29375, n29376, n29377, n29378, n29379, n29380,
         n29381, n29382, n29383, n29384, n29385, n29386, n29387, n29388,
         n29389, n29390, n29391, n29392, n29393, n29394, n29395, n29396,
         n29397, n29398, n29399, n29400, n29401, n29402, n29403, n29404,
         n29405, n29406, n29407, n29408, n29409, n29410, n29411, n29412,
         n29413, n29414, n29415, n29416, n29417, n29418, n29419, n29420,
         n29421, n29422, n29423, n29424, n29425, n29426, n29427, n29428,
         n29429, n29430, n29431, n29432, n29433, n29434, n29435, n29436,
         n29437, n29438, n29439, n29440, n29441, n29442, n29443, n29444,
         n29445, n29446, n29447, n29448, n29449, n29450, n29451, n29452,
         n29453, n29454, n29455, n29456, n29457, n29458, n29459, n29460,
         n29461, n29462, n29463, n29464, n29465, n29466, n29467, n29468,
         n29469, n29470, n29471, n29472, n29473, n29474, n29475, n29476,
         n29477, n29478, n29479, n29480, n29481, n29482, n29483, n29484,
         n29485, n29486, n29487, n29488, n29489, n29490, n29491, n29492,
         n29493, n29494, n29495, n29496, n29497, n29498, n29499, n29500,
         n29501, n29502, n29503, n29504, n29505, n29506, n29507, n29508,
         n29509, n29510, n29511, n29512, n29513, n29514, n29515, n29516,
         n29517, n29518, n29519, n29520, n29521, n29522, n29523, n29524,
         n29525, n29526, n29527, n29528, n29529, n29530, n29531, n29532,
         n29533, n29534, n29535, n29536, n29537, n29538, n29539, n29540,
         n29541, n29542, n29543, n29544, n29545, n29546, n29547, n29548,
         n29549, n29550, n29551, n29552, n29553, n29554, n29555, n29556,
         n29557, n29558, n29559, n29560, n29561, n29562, n29563, n29564,
         n29565, n29566, n29567, n29568, n29569, n29570, n29571, n29572,
         n29573, n29574, n29575, n29576, n29577, n29578, n29579, n29580,
         n29581, n29582, n29583, n29584, n29585, n29586, n29587, n29588,
         n29589, n29590, n29591, n29592, n29593, n29594, n29595, n29596,
         n29597, n29598, n29599, n29600, n29601, n29602, n29603, n29604,
         n29605, n29606, n29607, n29608, n29609, n29610, n29611, n29612,
         n29613, n29614, n29615, n29616, n29617, n29618, n29619, n29620,
         n29621, n29622, n29623, n29624, n29625, n29626, n29627, n29628,
         n29629, n29630, n29631, n29632, n29633, n29634, n29635, n29636,
         n29637, n29638, n29639, n29640, n29641, n29642, n29643, n29644,
         n29645, n29646, n29647, n29648, n29649, n29650, n29651, n29652,
         n29653, n29654, n29655, n29656, n29657, n29658, n29659, n29660,
         n29661, n29662, n29663, n29664, n29665, n29666, n29667, n29668,
         n29669, n29670, n29671, n29672, n29673, n29674, n29675, n29676,
         n29677, n29678, n29679, n29680, n29681, n29682, n29683, n29684,
         n29685, n29686, n29687, n29688, n29689, n29690, n29691, n29692,
         n29693, n29694, n29695, n29696, n29697, n29698, n29699, n29700,
         n29701, n29702, n29703, n29704, n29705, n29706, n29707, n29708,
         n29709, n29710, n29711, n29712, n29713, n29714, n29715, n29716,
         n29717, n29718, n29719, n29720, n29721, n29722, n29723, n29724,
         n29725, n29726, n29727, n29728, n29729, n29730, n29731, n29732,
         n29733, n29734, n29735, n29736, n29737, n29738, n29739, n29740,
         n29741, n29742, n29743, n29744, n29745, n29746, n29747, n29748,
         n29749, n29750, n29751, n29752, n29753, n29754, n29755, n29756,
         n29757, n29758, n29759, n29760, n29761, n29762, n29763, n29764,
         n29765, n29766, n29767, n29768, n29769, n29770, n29771, n29772,
         n29773, n29774, n29775, n29776, n29777, n29778, n29779, n29780,
         n29781, n29782, n29783, n29784, n29785, n29786, n29787, n29788,
         n29789, n29790, n29791, n29792, n29793, n29794, n29795, n29796,
         n29797, n29798, n29799, n29800, n29801, n29802, n29803, n29804,
         n29805, n29806, n29807, n29808, n29809, n29810, n29811, n29812,
         n29813, n29814, n29815, n29816, n29817, n29818, n29819, n29820,
         n29821, n29822, n29823, n29824, n29825, n29826, n29827, n29828,
         n29829, n29830, n29831, n29832, n29833, n29834, n29835, n29836,
         n29837, n29838, n29839, n29840, n29841, n29842, n29843, n29844,
         n29845, n29846, n29847, n29848, n29849, n29850, n29851, n29852,
         n29853, n29854, n29855, n29856, n29857, n29858, n29859, n29860,
         n29861, n29862, n29863, n29864, n29865, n29866, n29867, n29868,
         n29869, n29870, n29871, n29872, n29873, n29874, n29875, n29876,
         n29877, n29878, n29879, n29880, n29881, n29882, n29883, n29884,
         n29885, n29886, n29887, n29888, n29889, n29890, n29891, n29892,
         n29893, n29894, n29895, n29896, n29897, n29898, n29899, n29900,
         n29901, n29902, n29903, n29904, n29905, n29906, n29907, n29908,
         n29909, n29910, n29911, n29912, n29913, n29914, n29915, n29916,
         n29917, n29918, n29919, n29920, n29921, n29922, n29923, n29924,
         n29925, n29926, n29927, n29928, n29929, n29930, n29931, n29932,
         n29933, n29934, n29935, n29936, n29937, n29938, n29939, n29940,
         n29941, n29942, n29943, n29944, n29945, n29946, n29947, n29948,
         n29949, n29950, n29951, n29952, n29953, n29954, n29955, n29956,
         n29957, n29958, n29959, n29960, n29961, n29962, n29963, n29964,
         n29965, n29966, n29967, n29968, n29969, n29970, n29971, n29972,
         n29973, n29974, n29975, n29976, n29977, n29978, n29979, n29980,
         n29981, n29982, n29983, n29984, n29985, n29986, n29987, n29988,
         n29989, n29990, n29991, n29992, n29993, n29994, n29995, n29996,
         n29997, n29998, n29999, n30000, n30001, n30002, n30003, n30004,
         n30005, n30006, n30007, n30008, n30009, n30010, n30011, n30012,
         n30013, n30014, n30015, n30016, n30017, n30018, n30019, n30020,
         n30021, n30022, n30023, n30024, n30025, n30026, n30027, n30028,
         n30029, n30030, n30031, n30032, n30033, n30034, n30035, n30036,
         n30037, n30038, n30039, n30040, n30041, n30042, n30043, n30044,
         n30045, n30046, n30047, n30048, n30049, n30050, n30051, n30052,
         n30053, n30054, n30055, n30056, n30057, n30058, n30059, n30060,
         n30061, n30062, n30063, n30064, n30065, n30066, n30067, n30068,
         n30069, n30070, n30071, n30072, n30073, n30074, n30075, n30076,
         n30077, n30078, n30079, n30080, n30081, n30082, n30083, n30084,
         n30085, n30086, n30087, n30088, n30089, n30090, n30091, n30092,
         n30093, n30094, n30095, n30096, n30097, n30098, n30099, n30100,
         n30101, n30102, n30103, n30104, n30105, n30106, n30107, n30108,
         n30109, n30110, n30111, n30112, n30113, n30114, n30115, n30116,
         n30117, n30118, n30119, n30120, n30121, n30122, n30123, n30124,
         n30125, n30126, n30127, n30128, n30129, n30130, n30131, n30132,
         n30133, n30134, n30135, n30136, n30137, n30138, n30139, n30140,
         n30141, n30142, n30143, n30144, n30145, n30146, n30147, n30148,
         n30149, n30150, n30151, n30152, n30153, n30154, n30155, n30156,
         n30157, n30158, n30159, n30160, n30161, n30162, n30163, n30164,
         n30165, n30166, n30167, n30168, n30169, n30170, n30171, n30172,
         n30173, n30174, n30175, n30176, n30177, n30178, n30179, n30180,
         n30181, n30182, n30183, n30184, n30185, n30186, n30187, n30188,
         n30189, n30190, n30191, n30192, n30193, n30194, n30195, n30196,
         n30197, n30198, n30199, n30200, n30201, n30202, n30203, n30204,
         n30205, n30206, n30207, n30208, n30209, n30210, n30211, n30212,
         n30213, n30214, n30215, n30216, n30217, n30218, n30219, n30220,
         n30221, n30222, n30223, n30224, n30225, n30226, n30227, n30228,
         n30229, n30230, n30231, n30232, n30233, n30234, n30235, n30236,
         n30237, n30238, n30239, n30240, n30241, n30242, n30243, n30244,
         n30245, n30246, n30247, n30248, n30249, n30250, n30251, n30252,
         n30253, n30254, n30255, n30256, n30257, n30258, n30259, n30260,
         n30261, n30262, n30263, n30264, n30265, n30266, n30267, n30268,
         n30269, n30270, n30271, n30272, n30273, n30274, n30275, n30276,
         n30277, n30278, n30279, n30280, n30281, n30282, n30283, n30284,
         n30285, n30286, n30287, n30288, n30289, n30290, n30291, n30292,
         n30293, n30294, n30295, n30296, n30297, n30298, n30299, n30300,
         n30301, n30302, n30303, n30304, n30305, n30306, n30307, n30308,
         n30309, n30310, n30311, n30312, n30313, n30314, n30315, n30316,
         n30317, n30318, n30319, n30320, n30321, n30322, n30323, n30324,
         n30325, n30326, n30327, n30328, n30329, n30330, n30331, n30332,
         n30333, n30334, n30335, n30336, n30337, n30338, n30339, n30340,
         n30341, n30342, n30343, n30344, n30345, n30346, n30347, n30348,
         n30349, n30350, n30351, n30352, n30353, n30354, n30355, n30356,
         n30357, n30358, n30359, n30360, n30361, n30362, n30363, n30364,
         n30365, n30366, n30367, n30368, n30369, n30370, n30371, n30372,
         n30373, n30374, n30375, n30376, n30377, n30378, n30379, n30380,
         n30381, n30382, n30383, n30384, n30385, n30386, n30387, n30388,
         n30389, n30390, n30391, n30392, n30393, n30394, n30395, n30396,
         n30397, n30398, n30399, n30400, n30401, n30402, n30403, n30404,
         n30405, n30406, n30407, n30408, n30409, n30410, n30411, n30412,
         n30413, n30414, n30415, n30416, n30417, n30418, n30419, n30420,
         n30421, n30422, n30423, n30424, n30425, n30426, n30427, n30428,
         n30429, n30430, n30431, n30432, n30433, n30434, n30435, n30436,
         n30437, n30438, n30439, n30440, n30441, n30442, n30443, n30444,
         n30445, n30446, n30447, n30448, n30449, n30450, n30451, n30452,
         n30453, n30454, n30455, n30456, n30457, n30458, n30459, n30460,
         n30461, n30462, n30463, n30464, n30465, n30466, n30467, n30468,
         n30469, n30470, n30471, n30472, n30473, n30474, n30475, n30476,
         n30477, n30478, n30479, n30480, n30481, n30482, n30483, n30484,
         n30485, n30486, n30487, n30488, n30489, n30490, n30491, n30492,
         n30493, n30494, n30495, n30496, n30497, n30498, n30499, n30500,
         n30501, n30502, n30503, n30504, n30505, n30506, n30507, n30508,
         n30509, n30510, n30511, n30512, n30513, n30514, n30515, n30516,
         n30517, n30518, n30519, n30520, n30521, n30522, n30523, n30524,
         n30525, n30526, n30527, n30528, n30529, n30530, n30531, n30532,
         n30533, n30534, n30535, n30536, n30537, n30538, n30539, n30540,
         n30541, n30542, n30543, n30544, n30545, n30546, n30547, n30548,
         n30549, n30550, n30551, n30552, n30553, n30554, n30555, n30556,
         n30557, n30558, n30559, n30560, n30561, n30562, n30563, n30564,
         n30565, n30566, n30567, n30568, n30569, n30570, n30571, n30572,
         n30573, n30574, n30575, n30576, n30577, n30578, n30579, n30580,
         n30581, n30582, n30583, n30584, n30585, n30586, n30587, n30588,
         n30589, n30590, n30591, n30592, n30593, n30594, n30595, n30596,
         n30597, n30598, n30599, n30600, n30601, n30602, n30603, n30604,
         n30605, n30606, n30607, n30608, n30609, n30610, n30611, n30612,
         n30613, n30614, n30615, n30616, n30617, n30618, n30619, n30620,
         n30621, n30622, n30623, n30624, n30625, n30626, n30627, n30628,
         n30629, n30630, n30631, n30632, n30633, n30634, n30635, n30636,
         n30637, n30638, n30639, n30640, n30641, n30642, n30643, n30644,
         n30645, n30646, n30647, n30648, n30649, n30650, n30651, n30652,
         n30653, n30654, n30655, n30656, n30657, n30658, n30659, n30660,
         n30661, n30662, n30663, n30664, n30665, n30666, n30667, n30668,
         n30669, n30670, n30671, n30672, n30673, n30674, n30675, n30676,
         n30677, n30678, n30679, n30680, n30681, n30682, n30683, n30684,
         n30685, n30686, n30687, n30688, n30689, n30690, n30691, n30692,
         n30693, n30694, n30695, n30696, n30697, n30698, n30699, n30700,
         n30701, n30702, n30703, n30704, n30705, n30706, n30707, n30708,
         n30709, n30710, n30711, n30712, n30713, n30714, n30715, n30716,
         n30717, n30718, n30719, n30720, n30721, n30722, n30723, n30724,
         n30725, n30726, n30727, n30728, n30729, n30730, n30731, n30732,
         n30733, n30734, n30735, n30736, n30737, n30738, n30739, n30740,
         n30741, n30742, n30743, n30744, n30745, n30746, n30747, n30748,
         n30749, n30750, n30751, n30752, n30753, n30754, n30755, n30756,
         n30757, n30758, n30759, n30760, n30761, n30762, n30763, n30764,
         n30765, n30766, n30767, n30768, n30769, n30770, n30771, n30772,
         n30773, n30774, n30775, n30776, n30777, n30778, n30779, n30780,
         n30781, n30782, n30783, n30784, n30785, n30786, n30787, n30788,
         n30789, n30790, n30791, n30792, n30793, n30794, n30795, n30796,
         n30797, n30798, n30799, n30800, n30801, n30802, n30803, n30804,
         n30805, n30806, n30807, n30808, n30809, n30810, n30811, n30812,
         n30813, n30814, n30815, n30816, n30817, n30818, n30819, n30820,
         n30821, n30822, n30823, n30824, n30825, n30826, n30827, n30828,
         n30829, n30830, n30831, n30832, n30833, n30834, n30835, n30836,
         n30837, n30838, n30839, n30840, n30841, n30842, n30843, n30844,
         n30845, n30846, n30847, n30848, n30849, n30850, n30851, n30852,
         n30853, n30854, n30855, n30856, n30857, n30858, n30859, n30860,
         n30861, n30862, n30863, n30864, n30865, n30866, n30867, n30868,
         n30869, n30870, n30871, n30872, n30873, n30874, n30875, n30876,
         n30877, n30878, n30879, n30880, n30881, n30882, n30883, n30884,
         n30885, n30886, n30887, n30888, n30889, n30890, n30891, n30892,
         n30893, n30894, n30895, n30896, n30897, n30898, n30899, n30900,
         n30901, n30902, n30903, n30904, n30905, n30906, n30907, n30908,
         n30909, n30910, n30911, n30912, n30913, n30914, n30915, n30916,
         n30917, n30918, n30919, n30920, n30921, n30922, n30923, n30924,
         n30925, n30926, n30927, n30928, n30929, n30930, n30931, n30932,
         n30933, n30934, n30935, n30936, n30937, n30938, n30939, n30940,
         n30941, n30942, n30943, n30944, n30945, n30946, n30947, n30948,
         n30949, n30950, n30951, n30952, n30953, n30954, n30955, n30956,
         n30957, n30958, n30959, n30960, n30961, n30962, n30963, n30964,
         n30965, n30966, n30967, n30968, n30969, n30970, n30971, n30972,
         n30973, n30974, n30975, n30976, n30977, n30978, n30979, n30980,
         n30981, n30982, n30983, n30984, n30985, n30986, n30987, n30988,
         n30989, n30990, n30991, n30992, n30993, n30994, n30995, n30996,
         n30997, n30998, n30999, n31000, n31001, n31002, n31003, n31004,
         n31005, n31006, n31007, n31008, n31009, n31010, n31011, n31012,
         n31013, n31014, n31015, n31016, n31017, n31018, n31019, n31020,
         n31021, n31022, n31023, n31024, n31025, n31026, n31027, n31028,
         n31029, n31030, n31031, n31032, n31033, n31034, n31035, n31036,
         n31037, n31038, n31039, n31040, n31041, n31042, n31043, n31044,
         n31045, n31046, n31047, n31048, n31049, n31050, n31051, n31052,
         n31053, n31054, n31055, n31056, n31057, n31058, n31059, n31060,
         n31061, n31062, n31063, n31064, n31065, n31066, n31067, n31068,
         n31069, n31070, n31071, n31072, n31073, n31074, n31075, n31076,
         n31077, n31078, n31079, n31080, n31081, n31082, n31083, n31084,
         n31085, n31086, n31087, n31088, n31089, n31090, n31091, n31092,
         n31093, n31094, n31095, n31096, n31097, n31098, n31099, n31100,
         n31101, n31102, n31103, n31104, n31105, n31106, n31107, n31108,
         n31109, n31110, n31111, n31112, n31113, n31114, n31115, n31116,
         n31117, n31118, n31119, n31120, n31121, n31122, n31123, n31124,
         n31125, n31126, n31127, n31128, n31129, n31130, n31131, n31132,
         n31133, n31134, n31135, n31136, n31137, n31138, n31139, n31140,
         n31141, n31142, n31143, n31144, n31145, n31146, n31147, n31148,
         n31149, n31150, n31151, n31152, n31153, n31154, n31155, n31156,
         n31157, n31158, n31159, n31160, n31161, n31162, n31163, n31164,
         n31165, n31166, n31167, n31168, n31169, n31170, n31171, n31172,
         n31173, n31174, n31175, n31176, n31177, n31178, n31179, n31180,
         n31181, n31182, n31183, n31184, n31185, n31186, n31187, n31188,
         n31189, n31190, n31191, n31192, n31193, n31194, n31195, n31196,
         n31197, n31198, n31199, n31200, n31201, n31202, n31203, n31204,
         n31205, n31206, n31207, n31208, n31209, n31210, n31211, n31212,
         n31213, n31214, n31215, n31216, n31217, n31218, n31219, n31220,
         n31221, n31222, n31223, n31224, n31225, n31226, n31227, n31228,
         n31229, n31230, n31231, n31232, n31233, n31234, n31235, n31236,
         n31237, n31238, n31239, n31240, n31241, n31242, n31243, n31244,
         n31245, n31246, n31247, n31248, n31249, n31250, n31251, n31252,
         n31253, n31254, n31255, n31256, n31257, n31258, n31259, n31260,
         n31261, n31262, n31263, n31264, n31265, n31266, n31267, n31268,
         n31269, n31270, n31271, n31272, n31273, n31274, n31275, n31276,
         n31277, n31278, n31279, n31280, n31281, n31282, n31283, n31284,
         n31285, n31286, n31287, n31288, n31289, n31290, n31291, n31292,
         n31293, n31294, n31295, n31296, n31297, n31298, n31299, n31300,
         n31301, n31302, n31303, n31304, n31305, n31306, n31307, n31308,
         n31309, n31310, n31311, n31312, n31313, n31314, n31315, n31316,
         n31317, n31318, n31319, n31320, n31321, n31322, n31323, n31324,
         n31325, n31326, n31327, n31328, n31329, n31330, n31331, n31332,
         n31333, n31334, n31335, n31336, n31337, n31338, n31339, n31340,
         n31341, n31342, n31343, n31344, n31345, n31346, n31347, n31348,
         n31349, n31350, n31351, n31352, n31353, n31354, n31355, n31356,
         n31357, n31358, n31359, n31360, n31361, n31362, n31363, n31364,
         n31365, n31366, n31367, n31368, n31369, n31370, n31371, n31372,
         n31373, n31374, n31375, n31376, n31377, n31378, n31379, n31380,
         n31381, n31382, n31383, n31384, n31385, n31386, n31387, n31388,
         n31389, n31390, n31391, n31392, n31393, n31394, n31395, n31396,
         n31397, n31398, n31399, n31400, n31401, n31402, n31403, n31404,
         n31405, n31406, n31407, n31408, n31409, n31410, n31411, n31412,
         n31413, n31414, n31415, n31416, n31417, n31418, n31419, n31420,
         n31421, n31422, n31423, n31424, n31425, n31426, n31427, n31428,
         n31429, n31430, n31431, n31432, n31433, n31434, n31435, n31436,
         n31437, n31438, n31439, n31440, n31441, n31442, n31443, n31444,
         n31445, n31446, n31447, n31448, n31449, n31450, n31451, n31452,
         n31453, n31454, n31455, n31456, n31457, n31458, n31459, n31460,
         n31461, n31462, n31463, n31464, n31465, n31466, n31467, n31468,
         n31469, n31470, n31471, n31472, n31473, n31474, n31475, n31476,
         n31477, n31478, n31479, n31480, n31481, n31482, n31483, n31484,
         n31485, n31486, n31487, n31488, n31489, n31490, n31491, n31492,
         n31493, n31494, n31495, n31496, n31497, n31498, n31499, n31500,
         n31501, n31502, n31503, n31504, n31505, n31506, n31507, n31508,
         n31509, n31510, n31511, n31512, n31513, n31514, n31515, n31516,
         n31517, n31518, n31519, n31520, n31521, n31522, n31523, n31524,
         n31525, n31526, n31527, n31528, n31529, n31530, n31531, n31532,
         n31533, n31534, n31535, n31536, n31537, n31538, n31539, n31540,
         n31541, n31542, n31543, n31544, n31545, n31546, n31547, n31548,
         n31549, n31550, n31551, n31552, n31553, n31554, n31555, n31556,
         n31557, n31558, n31559, n31560, n31561, n31562, n31563, n31564,
         n31565, n31566, n31567, n31568, n31569, n31570, n31571, n31572,
         n31573, n31574, n31575, n31576, n31577, n31578, n31579, n31580,
         n31581, n31582, n31583, n31584, n31585, n31586, n31587, n31588,
         n31589, n31590, n31591, n31592, n31593, n31594, n31595, n31596,
         n31597, n31598, n31599, n31600, n31601, n31602, n31603, n31604,
         n31605, n31606, n31607, n31608, n31609, n31610, n31611, n31612,
         n31613, n31614, n31615, n31616, n31617, n31618, n31619, n31620,
         n31621, n31622, n31623, n31624, n31625, n31626, n31627, n31628,
         n31629, n31630, n31631, n31632, n31633, n31634, n31635, n31636,
         n31637, n31638, n31639, n31640, n31641, n31642, n31643, n31644,
         n31645, n31646, n31647, n31648, n31649, n31650, n31651, n31652,
         n31653, n31654, n31655, n31656, n31657, n31658, n31659, n31660,
         n31661, n31662, n31663, n31664, n31665, n31666, n31667, n31668,
         n31669, n31670, n31671, n31672, n31673, n31674, n31675, n31676,
         n31677, n31678, n31679, n31680, n31681, n31682, n31683, n31684,
         n31685, n31686, n31687, n31688, n31689, n31690, n31691, n31692,
         n31693, n31694, n31695, n31696, n31697, n31698, n31699, n31700,
         n31701, n31702, n31703, n31704, n31705, n31706, n31707, n31708,
         n31709, n31710, n31711, n31712, n31713, n31714, n31715, n31716,
         n31717, n31718, n31719, n31720, n31721, n31722, n31723, n31724,
         n31725, n31726, n31727, n31728, n31729, n31730, n31731, n31732,
         n31733, n31734, n31735, n31736, n31737, n31738, n31739, n31740,
         n31741, n31742, n31743, n31744, n31745, n31746, n31747, n31748,
         n31749, n31750, n31751, n31752, n31753, n31754, n31755, n31756,
         n31757, n31758, n31759, n31760, n31761, n31762, n31763, n31764,
         n31765, n31766, n31767, n31768, n31769, n31770, n31771, n31772,
         n31773, n31774, n31775, n31776, n31777, n31778, n31779, n31780,
         n31781, n31782, n31783, n31784, n31785, n31786, n31787, n31788,
         n31789, n31790, n31791, n31792, n31793, n31794, n31795, n31796,
         n31797, n31798, n31799, n31800, n31801, n31802, n31803, n31804,
         n31805, n31806, n31807, n31808, n31809, n31810, n31811, n31812,
         n31813, n31814, n31815, n31816, n31817, n31818, n31819, n31820,
         n31821, n31822, n31823, n31824, n31825, n31826, n31827, n31828,
         n31829, n31830, n31831, n31832, n31833, n31834, n31835, n31836,
         n31837, n31838, n31839, n31840, n31841, n31842, n31843, n31844,
         n31845, n31846, n31847, n31848, n31849, n31850, n31851, n31852,
         n31853, n31854, n31855, n31856, n31857, n31858, n31859, n31860,
         n31861, n31862, n31863, n31864, n31865, n31866, n31867, n31868,
         n31869, n31870, n31871, n31872, n31873, n31874, n31875, n31876,
         n31877, n31878, n31879, n31880, n31881, n31882, n31883, n31884,
         n31885, n31886, n31887, n31888, n31889, n31890, n31891, n31892,
         n31893, n31894, n31895, n31896, n31897, n31898, n31899, n31900,
         n31901, n31902, n31903, n31904, n31905, n31906, n31907, n31908,
         n31909, n31910, n31911, n31912, n31913, n31914, n31915, n31916,
         n31917, n31918, n31919, n31920, n31921, n31922, n31923, n31924,
         n31925, n31926, n31927, n31928, n31929, n31930, n31931, n31932,
         n31933, n31934, n31935, n31936, n31937, n31938, n31939, n31940,
         n31941, n31942, n31943, n31944, n31945, n31946, n31947, n31948,
         n31949, n31950, n31951, n31952, n31953, n31954, n31955, n31956,
         n31957, n31958, n31959, n31960, n31961, n31962, n31963, n31964,
         n31965, n31966, n31967, n31968, n31969, n31970, n31971, n31972,
         n31973, n31974, n31975, n31976, n31977, n31978, n31979, n31980,
         n31981, n31982, n31983, n31984, n31985, n31986, n31987, n31988,
         n31989, n31990, n31991, n31992, n31993, n31994, n31995, n31996,
         n31997, n31998, n31999, n32000, n32001, n32002, n32003, n32004,
         n32005, n32006, n32007, n32008, n32009, n32010, n32011, n32012,
         n32013, n32014, n32015, n32016, n32017, n32018, n32019, n32020,
         n32021, n32022, n32023, n32024, n32025, n32026, n32027, n32028,
         n32029, n32030, n32031, n32032, n32033, n32034, n32035, n32036,
         n32037, n32038, n32039, n32040, n32041, n32042, n32043, n32044,
         n32045, n32046, n32047, n32048, n32049, n32050, n32051, n32052,
         n32053, n32054, n32055, n32056, n32057, n32058, n32059, n32060,
         n32061, n32062, n32063, n32064, n32065, n32066, n32067, n32068,
         n32069, n32070, n32071, n32072, n32073, n32074, n32075, n32076,
         n32077, n32078, n32079, n32080, n32081, n32082, n32083, n32084,
         n32085, n32086, n32087, n32088, n32089, n32090, n32091, n32092,
         n32093, n32094, n32095, n32096, n32097, n32098, n32099, n32100,
         n32101, n32102, n32103, n32104, n32105, n32106, n32107, n32108,
         n32109, n32110, n32111, n32112, n32113, n32114, n32115, n32116,
         n32117, n32118, n32119, n32120, n32121, n32122, n32123, n32124,
         n32125, n32126, n32127, n32128, n32129, n32130, n32131, n32132,
         n32133, n32134, n32135, n32136, n32137, n32138, n32139, n32140,
         n32141, n32142, n32143, n32144, n32145, n32146, n32147, n32148,
         n32149, n32150, n32151, n32152, n32153, n32154, n32155, n32156,
         n32157, n32158, n32159, n32160, n32161, n32162, n32163, n32164,
         n32165, n32166, n32167, n32168, n32169, n32170, n32171, n32172,
         n32173, n32174, n32175, n32176, n32177, n32178, n32179, n32180,
         n32181, n32182, n32183, n32184, n32185, n32186, n32187, n32188,
         n32189, n32190, n32191, n32192, n32193, n32194, n32195, n32196,
         n32197, n32198, n32199, n32200, n32201, n32202, n32203, n32204,
         n32205, n32206, n32207, n32208, n32209, n32210, n32211, n32212,
         n32213, n32214, n32215, n32216, n32217, n32218, n32219, n32220,
         n32221, n32222, n32223, n32224, n32225, n32226, n32227, n32228,
         n32229, n32230, n32231, n32232, n32233, n32234, n32235, n32236,
         n32237, n32238, n32239, n32240, n32241, n32242, n32243, n32244,
         n32245, n32246, n32247, n32248, n32249, n32250, n32251, n32252,
         n32253, n32254, n32255, n32256, n32257, n32258, n32259, n32260,
         n32261, n32262, n32263, n32264, n32265, n32266, n32267, n32268,
         n32269, n32270, n32271, n32272, n32273, n32274, n32275, n32276,
         n32277, n32278, n32279, n32280, n32281, n32282, n32283, n32284,
         n32285, n32286, n32287, n32288, n32289, n32290, n32291, n32292,
         n32293, n32294, n32295, n32296, n32297, n32298, n32299, n32300,
         n32301, n32302, n32303, n32304, n32305, n32306, n32307, n32308,
         n32309, n32310, n32311, n32312, n32313, n32314, n32315, n32316,
         n32317, n32318, n32319, n32320, n32321, n32322, n32323, n32324,
         n32325, n32326, n32327, n32328, n32329, n32330, n32331, n32332,
         n32333, n32334, n32335, n32336, n32337, n32338, n32339, n32340,
         n32341, n32342, n32343, n32344, n32345, n32346, n32347, n32348,
         n32349, n32350, n32351, n32352, n32353, n32354, n32355, n32356,
         n32357, n32358, n32359, n32360, n32361, n32362, n32363, n32364,
         n32365, n32366, n32367, n32368, n32369, n32370, n32371, n32372,
         n32373, n32374, n32375, n32376, n32377, n32378, n32379, n32380,
         n32381, n32382, n32383, n32384, n32385, n32386, n32387, n32388,
         n32389, n32390, n32391, n32392, n32393, n32394, n32395, n32396,
         n32397, n32398, n32399, n32400, n32401, n32402, n32403, n32404,
         n32405, n32406, n32407, n32408, n32409, n32410, n32411, n32412,
         n32413, n32414, n32415, n32416, n32417, n32418, n32419, n32420,
         n32421, n32422, n32423, n32424, n32425, n32426, n32427, n32428,
         n32429, n32430, n32431, n32432, n32433, n32434, n32435, n32436,
         n32437, n32438, n32439, n32440, n32441, n32442, n32443, n32444,
         n32445, n32446, n32447, n32448, n32449, n32450, n32451, n32452,
         n32453, n32454, n32455, n32456, n32457, n32458, n32459, n32460,
         n32461, n32462, n32463, n32464, n32465, n32466, n32467, n32468,
         n32469, n32470, n32471, n32472, n32473, n32474, n32475, n32476,
         n32477, n32478, n32479, n32480, n32481, n32482, n32483, n32484,
         n32485, n32486, n32487, n32488, n32489, n32490, n32491, n32492,
         n32493, n32494, n32495, n32496, n32497, n32498, n32499, n32500,
         n32501, n32502, n32503, n32504, n32505, n32506, n32507, n32508,
         n32509, n32510, n32511, n32512, n32513, n32514, n32515, n32516,
         n32517, n32518, n32519, n32520, n32521, n32522, n32523, n32524,
         n32525, n32526, n32527, n32528, n32529, n32530, n32531, n32532,
         n32533, n32534, n32535, n32536, n32537, n32538, n32539, n32540,
         n32541, n32542, n32543, n32544, n32545, n32546, n32547, n32548,
         n32549, n32550, n32551, n32552, n32553, n32554, n32555, n32556,
         n32557, n32558, n32559, n32560, n32561, n32562, n32563, n32564,
         n32565, n32566, n32567, n32568, n32569, n32570, n32571, n32572,
         n32573, n32574, n32575, n32576, n32577, n32578, n32579, n32580,
         n32581, n32582, n32583, n32584, n32585, n32586, n32587, n32588,
         n32589, n32590, n32591, n32592, n32593, n32594, n32595, n32596,
         n32597, n32598, n32599, n32600, n32601, n32602, n32603, n32604,
         n32605, n32606, n32607, n32608, n32609, n32610, n32611, n32612,
         n32613, n32614, n32615, n32616, n32617, n32618, n32619, n32620,
         n32621, n32622, n32623, n32624, n32625, n32626, n32627, n32628,
         n32629, n32630, n32631, n32632, n32633, n32634, n32635, n32636,
         n32637, n32638, n32639, n32640, n32641, n32642, n32643, n32644,
         n32645, n32646, n32647, n32648, n32649, n32650, n32651, n32652,
         n32653, n32654, n32655, n32656, n32657, n32658, n32659, n32660,
         n32661, n32662, n32663, n32664, n32665, n32666, n32667, n32668,
         n32669, n32670, n32671, n32672, n32673, n32674, n32675, n32676,
         n32677, n32678, n32679, n32680, n32681, n32682, n32683, n32684,
         n32685, n32686, n32687, n32688, n32689, n32690, n32691, n32692,
         n32693, n32694, n32695, n32696, n32697, n32698, n32699, n32700,
         n32701, n32702, n32703, n32704, n32705, n32706, n32707, n32708,
         n32709, n32710, n32711, n32712, n32713, n32714, n32715, n32716,
         n32717, n32718, n32719, n32720, n32721, n32722, n32723, n32724,
         n32725, n32726, n32727, n32728, n32729, n32730, n32731, n32732,
         n32733, n32734, n32735, n32736, n32737, n32738, n32739, n32740,
         n32741, n32742, n32743, n32744, n32745, n32746, n32747, n32748,
         n32749, n32750, n32751, n32752, n32753, n32754, n32755, n32756,
         n32757, n32758, n32759, n32760, n32761, n32762, n32763, n32764,
         n32765, n32766, n32767, n32768, n32769, n32770, n32771, n32772,
         n32773, n32774, n32775, n32776, n32777, n32778, n32779, n32780,
         n32781, n32782, n32783, n32784, n32785, n32786, n32787, n32788,
         n32789, n32790, n32791, n32792, n32793, n32794, n32795, n32796,
         n32797, n32798, n32799, n32800, n32801, n32802, n32803, n32804,
         n32805, n32806, n32807, n32808, n32809, n32810, n32811, n32812,
         n32813, n32814, n32815, n32816, n32817, n32818, n32819, n32820,
         n32821, n32822, n32823, n32824, n32825, n32826, n32827, n32828,
         n32829, n32830, n32831, n32832, n32833, n32834, n32835, n32836,
         n32837, n32838, n32839, n32840, n32841, n32842, n32843, n32844,
         n32845, n32846, n32847, n32848, n32849, n32850, n32851, n32852,
         n32853, n32854, n32855, n32856, n32857, n32858, n32859, n32860,
         n32861, n32862, n32863, n32864, n32865, n32866, n32867, n32868,
         n32869, n32870, n32871, n32872, n32873, n32874, n32875, n32876,
         n32877, n32878, n32879, n32880, n32881, n32882, n32883, n32884,
         n32885, n32886, n32887, n32888, n32889, n32890, n32891, n32892,
         n32893, n32894, n32895, n32896, n32897, n32898, n32899, n32900,
         n32901, n32902, n32903, n32904, n32905, n32906, n32907, n32908,
         n32909, n32910, n32911, n32912, n32913, n32914, n32915, n32916,
         n32917, n32918, n32919, n32920, n32921, n32922, n32923, n32924,
         n32925, n32926, n32927, n32928, n32929, n32930, n32931, n32932,
         n32933, n32934, n32935, n32936, n32937, n32938, n32939, n32940,
         n32941, n32942, n32943, n32944, n32945, n32946, n32947, n32948,
         n32949, n32950, n32951, n32952, n32953, n32954, n32955, n32956,
         n32957, n32958, n32959, n32960, n32961, n32962, n32963, n32964,
         n32965, n32966, n32967, n32968, n32969, n32970, n32971, n32972,
         n32973, n32974, n32975, n32976, n32977, n32978, n32979, n32980,
         n32981, n32982, n32983, n32984, n32985, n32986, n32987, n32988,
         n32989, n32990, n32991, n32992, n32993, n32994, n32995, n32996,
         n32997, n32998, n32999, n33000, n33001, n33002, n33003, n33004,
         n33005, n33006, n33007, n33008, n33009, n33010, n33011, n33012,
         n33013, n33014, n33015, n33016, n33017, n33018, n33019, n33020,
         n33021, n33022, n33023, n33024, n33025, n33026, n33027, n33028,
         n33029, n33030, n33031, n33032, n33033, n33034, n33035, n33036,
         n33037, n33038, n33039, n33040, n33041, n33042, n33043, n33044,
         n33045, n33046, n33047, n33048, n33049, n33050, n33051, n33052,
         n33053, n33054, n33055, n33056, n33057, n33058, n33059, n33060,
         n33061, n33062, n33063, n33064, n33065, n33066, n33067, n33068,
         n33069, n33070, n33071, n33072, n33073, n33074, n33075, n33076,
         n33077, n33078, n33079, n33080, n33081, n33082, n33083, n33084,
         n33085, n33086, n33087, n33088, n33089, n33090, n33091, n33092,
         n33093, n33094, n33095, n33096, n33097, n33098, n33099, n33100,
         n33101, n33102, n33103, n33104, n33105, n33106, n33107, n33108,
         n33109, n33110, n33111, n33112, n33113, n33114, n33115, n33116,
         n33117, n33118, n33119, n33120, n33121, n33122, n33123, n33124,
         n33125, n33126, n33127, n33128, n33129, n33130, n33131, n33132,
         n33133, n33134, n33135, n33136, n33137, n33138, n33139, n33140,
         n33141, n33142, n33143, n33144, n33145, n33146, n33147, n33148,
         n33149, n33150, n33151, n33152, n33153, n33154, n33155, n33156,
         n33157, n33158, n33159, n33160, n33161, n33162, n33163, n33164,
         n33165, n33166, n33167, n33168, n33169, n33170, n33171, n33172,
         n33173, n33174, n33175, n33176, n33177, n33178, n33179, n33180,
         n33181, n33182, n33183, n33184, n33185, n33186, n33187, n33188,
         n33189, n33190, n33191, n33192, n33193, n33194, n33195, n33196,
         n33197, n33198, n33199, n33200, n33201, n33202, n33203, n33204,
         n33205, n33206, n33207, n33208, n33209, n33210, n33211, n33212,
         n33213, n33214, n33215, n33216, n33217, n33218, n33219, n33220,
         n33221, n33222, n33223, n33224, n33225, n33226, n33227, n33228,
         n33229, n33230, n33231, n33232, n33233, n33234, n33235, n33236,
         n33237, n33238, n33239, n33240, n33241, n33242, n33243, n33244,
         n33245, n33246, n33247, n33248, n33249, n33250, n33251, n33252,
         n33253, n33254, n33255, n33256, n33257, n33258, n33259, n33260,
         n33261, n33262, n33263, n33264, n33265, n33266, n33267, n33268,
         n33269, n33270, n33271, n33272, n33273, n33274, n33275, n33276,
         n33277, n33278, n33279, n33280, n33281, n33282, n33283, n33284,
         n33285, n33286, n33287, n33288, n33289, n33290, n33291, n33292,
         n33293, n33294, n33295, n33296, n33297, n33298, n33299, n33300,
         n33301, n33302, n33303, n33304, n33305, n33306, n33307, n33308,
         n33309, n33310, n33311, n33312, n33313, n33314, n33315, n33316,
         n33317, n33318, n33319, n33320, n33321, n33322, n33323, n33324,
         n33325, n33326, n33327, n33328, n33329, n33330, n33331, n33332,
         n33333, n33334, n33335, n33336, n33337, n33338, n33339, n33340,
         n33341, n33342, n33343, n33344, n33345, n33346, n33347, n33348,
         n33349, n33350, n33351, n33352, n33353, n33354, n33355, n33356,
         n33357, n33358, n33359, n33360, n33361, n33362, n33363, n33364,
         n33365, n33366, n33367, n33368, n33369, n33370, n33371, n33372,
         n33373, n33374, n33375, n33376, n33377, n33378, n33379, n33380,
         n33381, n33382, n33383, n33384, n33385, n33386, n33387, n33388,
         n33389, n33390, n33391, n33392, n33393, n33394, n33395, n33396,
         n33397, n33398, n33399, n33400, n33401, n33402, n33403, n33404,
         n33405, n33406, n33407, n33408, n33409, n33410, n33411, n33412,
         n33413, n33414, n33415, n33416, n33417, n33418, n33419, n33420,
         n33421, n33422, n33423, n33424, n33425, n33426, n33427, n33428,
         n33429, n33430, n33431, n33432, n33433, n33434, n33435, n33436,
         n33437, n33438, n33439, n33440, n33441, n33442, n33443, n33444,
         n33445, n33446, n33447, n33448, n33449, n33450, n33451, n33452,
         n33453, n33454, n33455, n33456, n33457, n33458, n33459, n33460,
         n33461, n33462, n33463, n33464, n33465, n33466, n33467, n33468,
         n33469, n33470, n33471, n33472, n33473, n33474, n33475, n33476,
         n33477, n33478, n33479, n33480, n33481, n33482, n33483, n33484,
         n33485, n33486, n33487, n33488, n33489, n33490, n33491, n33492,
         n33493, n33494, n33495, n33496, n33497, n33498, n33499, n33500,
         n33501, n33502, n33503, n33504, n33505, n33506, n33507, n33508,
         n33509, n33510, n33511, n33512, n33513, n33514, n33515, n33516,
         n33517, n33518, n33519, n33520, n33521, n33522, n33523, n33524,
         n33525, n33526, n33527, n33528, n33529, n33530, n33531, n33532,
         n33533, n33534, n33535, n33536, n33537, n33538, n33539, n33540,
         n33541, n33542, n33543, n33544, n33545, n33546, n33547, n33548,
         n33549, n33550, n33551, n33552, n33553, n33554, n33555, n33556,
         n33557, n33558, n33559, n33560, n33561, n33562, n33563, n33564,
         n33565, n33566, n33567, n33568, n33569, n33570, n33571, n33572,
         n33573, n33574, n33575, n33576, n33577, n33578, n33579, n33580,
         n33581, n33582, n33583, n33584, n33585, n33586, n33587, n33588,
         n33589, n33590, n33591, n33592, n33593, n33594, n33595, n33596,
         n33597, n33598, n33599, n33600, n33601, n33602, n33603, n33604,
         n33605, n33606, n33607, n33608, n33609, n33610, n33611, n33612,
         n33613, n33614, n33615, n33616, n33617, n33618, n33619, n33620,
         n33621, n33622, n33623, n33624, n33625, n33626, n33627, n33628,
         n33629, n33630, n33631, n33632, n33633, n33634, n33635, n33636,
         n33637, n33638, n33639, n33640, n33641, n33642, n33643, n33644,
         n33645, n33646, n33647, n33648, n33649, n33650, n33651, n33652,
         n33653, n33654, n33655, n33656, n33657, n33658, n33659, n33660,
         n33661, n33662, n33663, n33664, n33665, n33666, n33667, n33668,
         n33669, n33670, n33671, n33672, n33673, n33674, n33675, n33676,
         n33677, n33678, n33679, n33680, n33681, n33682, n33683, n33684,
         n33685, n33686, n33687, n33688, n33689, n33690, n33691, n33692,
         n33693, n33694, n33695, n33696, n33697, n33698, n33699, n33700,
         n33701, n33702, n33703, n33704, n33705, n33706, n33707, n33708,
         n33709, n33710, n33711, n33712, n33713, n33714, n33715, n33716,
         n33717, n33718, n33719, n33720, n33721, n33722, n33723, n33724,
         n33725, n33726, n33727, n33728, n33729, n33730, n33731, n33732,
         n33733, n33734, n33735, n33736, n33737, n33738, n33739, n33740,
         n33741, n33742, n33743, n33744, n33745, n33746, n33747, n33748,
         n33749, n33750, n33751, n33752, n33753, n33754, n33755, n33756,
         n33757, n33758, n33759, n33760, n33761, n33762, n33763, n33764,
         n33765, n33766, n33767, n33768, n33769, n33770, n33771, n33772,
         n33773, n33774, n33775, n33776, n33777, n33778, n33779, n33780,
         n33781, n33782, n33783, n33784, n33785, n33786, n33787, n33788,
         n33789, n33790, n33791, n33792, n33793, n33794, n33795, n33796,
         n33797, n33798, n33799, n33800, n33801, n33802, n33803, n33804,
         n33805, n33806, n33807, n33808, n33809, n33810, n33811, n33812,
         n33813, n33814, n33815, n33816, n33817, n33818, n33819, n33820,
         n33821, n33822, n33823, n33824, n33825, n33826, n33827, n33828,
         n33829, n33830, n33831, n33832, n33833, n33834, n33835, n33836,
         n33837, n33838, n33839, n33840, n33841, n33842, n33843, n33844,
         n33845, n33846, n33847, n33848, n33849, n33850, n33851, n33852,
         n33853, n33854, n33855, n33856, n33857, n33858, n33859, n33860,
         n33861, n33862, n33863, n33864, n33865, n33866, n33867, n33868,
         n33869, n33870, n33871, n33872, n33873, n33874, n33875, n33876,
         n33877, n33878, n33879, n33880, n33881, n33882, n33883, n33884,
         n33885, n33886, n33887, n33888, n33889, n33890, n33891, n33892,
         n33893, n33894, n33895, n33896, n33897, n33898, n33899, n33900,
         n33901, n33902, n33903, n33904, n33905, n33906, n33907, n33908,
         n33909, n33910, n33911, n33912, n33913, n33914, n33915, n33916,
         n33917, n33918, n33919, n33920, n33921, n33922, n33923, n33924,
         n33925, n33926, n33927, n33928, n33929, n33930, n33931, n33932,
         n33933, n33934, n33935, n33936, n33937, n33938, n33939, n33940,
         n33941, n33942, n33943, n33944, n33945, n33946, n33947, n33948,
         n33949, n33950, n33951, n33952, n33953, n33954, n33955, n33956,
         n33957, n33958, n33959, n33960, n33961, n33962, n33963, n33964,
         n33965, n33966, n33967, n33968, n33969, n33970, n33971, n33972,
         n33973, n33974, n33975, n33976, n33977, n33978, n33979, n33980,
         n33981, n33982, n33983, n33984, n33985, n33986, n33987, n33988,
         n33989, n33990, n33991, n33992, n33993, n33994, n33995, n33996,
         n33997, n33998, n33999, n34000, n34001, n34002, n34003, n34004,
         n34005, n34006, n34007, n34008, n34009, n34010, n34011, n34012,
         n34013, n34014, n34015, n34016, n34017, n34018, n34019, n34020,
         n34021, n34022, n34023, n34024, n34025, n34026, n34027, n34028,
         n34029, n34030, n34031, n34032, n34033, n34034, n34035, n34036,
         n34037, n34038, n34039, n34040, n34041, n34042, n34043, n34044,
         n34045, n34046, n34047, n34048, n34049, n34050, n34051, n34052,
         n34053, n34054, n34055, n34056, n34057, n34058, n34059, n34060,
         n34061, n34062, n34063, n34064, n34065, n34066, n34067, n34068,
         n34069, n34070, n34071, n34072, n34073, n34074, n34075, n34076,
         n34077, n34078, n34079, n34080, n34081, n34082, n34083, n34084,
         n34085, n34086, n34087, n34088, n34089, n34090, n34091, n34092,
         n34093, n34094, n34095, n34096, n34097, n34098, n34099, n34100,
         n34101, n34102, n34103, n34104, n34105, n34106, n34107, n34108,
         n34109, n34110, n34111, n34112, n34113, n34114, n34115, n34116,
         n34117, n34118, n34119, n34120, n34121, n34122, n34123, n34124,
         n34125, n34126, n34127, n34128, n34129, n34130, n34131, n34132,
         n34133, n34134, n34135, n34136, n34137, n34138, n34139, n34140,
         n34141, n34142, n34143, n34144, n34145, n34146, n34147, n34148,
         n34149, n34150, n34151, n34152, n34153, n34154, n34155, n34156,
         n34157, n34158, n34159, n34160, n34161, n34162, n34163, n34164,
         n34165, n34166, n34167, n34168, n34169, n34170, n34171, n34172,
         n34173, n34174, n34175, n34176, n34177, n34178, n34179, n34180,
         n34181, n34182, n34183, n34184, n34185, n34186, n34187, n34188,
         n34189, n34190, n34191, n34192, n34193, n34194, n34195, n34196,
         n34197, n34198, n34199, n34200, n34201, n34202, n34203, n34204,
         n34205, n34206, n34207, n34208, n34209, n34210, n34211, n34212,
         n34213, n34214, n34215, n34216, n34217, n34218, n34219, n34220,
         n34221, n34222, n34223, n34224, n34225, n34226, n34227, n34228,
         n34229, n34230, n34231, n34232, n34233, n34234, n34235, n34236,
         n34237, n34238, n34239, n34240, n34241, n34242, n34243, n34244,
         n34245, n34246, n34247, n34248, n34249, n34250, n34251, n34252,
         n34253, n34254, n34255, n34256, n34257, n34258, n34259, n34260,
         n34261, n34262, n34263, n34264, n34265, n34266, n34267, n34268,
         n34269, n34270, n34271, n34272, n34273, n34274, n34275, n34276,
         n34277, n34278, n34279, n34280, n34281, n34282, n34283, n34284,
         n34285, n34286, n34287, n34288, n34289, n34290, n34291, n34292,
         n34293, n34294, n34295, n34296, n34297, n34298, n34299, n34300,
         n34301, n34302, n34303, n34304, n34305, n34306, n34307, n34308,
         n34309, n34310, n34311, n34312, n34313, n34314, n34315, n34316,
         n34317, n34318, n34319, n34320, n34321, n34322, n34323, n34324,
         n34325, n34326, n34327, n34328, n34329, n34330, n34331, n34332,
         n34333, n34334, n34335, n34336, n34337, n34338, n34339, n34340,
         n34341, n34342, n34343, n34344, n34345, n34346, n34347, n34348,
         n34349, n34350, n34351, n34352, n34353, n34354, n34355, n34356,
         n34357, n34358, n34359, n34360, n34361, n34362, n34363, n34364,
         n34365, n34366, n34367, n34368, n34369, n34370, n34371, n34372,
         n34373, n34374, n34375, n34376, n34377, n34378, n34379, n34380,
         n34381, n34382, n34383, n34384, n34385, n34386, n34387, n34388,
         n34389, n34390, n34391, n34392, n34393, n34394, n34395, n34396,
         n34397, n34398, n34399, n34400, n34401, n34402, n34403, n34404,
         n34405, n34406, n34407, n34408, n34409, n34410, n34411, n34412,
         n34413, n34414, n34415, n34416, n34417, n34418, n34419, n34420,
         n34421, n34422, n34423, n34424, n34425, n34426, n34427, n34428,
         n34429, n34430, n34431, n34432, n34433, n34434, n34435, n34436,
         n34437, n34438, n34439, n34440, n34441, n34442, n34443, n34444,
         n34445, n34446, n34447, n34448, n34449, n34450, n34451, n34452,
         n34453, n34454, n34455, n34456, n34457, n34458, n34459, n34460,
         n34461, n34462, n34463, n34464, n34465, n34466, n34467, n34468,
         n34469, n34470, n34471, n34472, n34473, n34474, n34475, n34476,
         n34477, n34478, n34479, n34480, n34481, n34482, n34483, n34484,
         n34485, n34486, n34487, n34488, n34489, n34490, n34491, n34492,
         n34493, n34494, n34495, n34496, n34497, n34498, n34499, n34500,
         n34501, n34502, n34503, n34504, n34505, n34506, n34507, n34508,
         n34509, n34510, n34511, n34512, n34513, n34514, n34515, n34516,
         n34517, n34518, n34519, n34520, n34521, n34522, n34523, n34524,
         n34525, n34526, n34527, n34528, n34529, n34530, n34531, n34532,
         n34533, n34534, n34535, n34536, n34537, n34538, n34539, n34540,
         n34541, n34542, n34543, n34544, n34545, n34546, n34547, n34548,
         n34549, n34550, n34551, n34552, n34553, n34554, n34555, n34556,
         n34557, n34558, n34559, n34560, n34561, n34562, n34563, n34564,
         n34565, n34566, n34567, n34568, n34569, n34570, n34571, n34572,
         n34573, n34574, n34575, n34576, n34577, n34578, n34579, n34580,
         n34581, n34582, n34583, n34584, n34585, n34586, n34587, n34588,
         n34589, n34590, n34591, n34592, n34593, n34594, n34595, n34596,
         n34597, n34598, n34599, n34600, n34601, n34602, n34603, n34604,
         n34605, n34606, n34607, n34608, n34609, n34610, n34611, n34612,
         n34613, n34614, n34615, n34616, n34617, n34618, n34619, n34620,
         n34621, n34622, n34623, n34624, n34625, n34626, n34627, n34628,
         n34629, n34630, n34631, n34632, n34633, n34634, n34635, n34636,
         n34637, n34638, n34639, n34640, n34641, n34642, n34643, n34644,
         n34645, n34646, n34647, n34648, n34649, n34650, n34651, n34652,
         n34653, n34654, n34655, n34656, n34657, n34658, n34659, n34660,
         n34661, n34662, n34663, n34664, n34665, n34666, n34667, n34668,
         n34669, n34670, n34671, n34672, n34673, n34674, n34675, n34676,
         n34677, n34678, n34679, n34680, n34681, n34682, n34683, n34684,
         n34685, n34686, n34687, n34688, n34689, n34690, n34691, n34692,
         n34693, n34694, n34695, n34696, n34697;
  wire   [31:0] m0s0_data_i;
  wire   [31:0] m0s0_data_o;
  wire   [31:0] m0s0_addr;
  wire   [3:0] m0s0_sel;
  wire   [31:0] m0s1_data_i;
  wire   [31:0] m0s2_data_i;
  wire   [31:0] m0s3_data_i;
  wire   [31:0] m0s4_data_i;
  wire   [31:0] m0s5_data_i;
  wire   [31:0] m0s6_data_i;
  wire   [31:0] m0s7_data_i;
  wire   [31:0] m0s8_data_i;
  wire   [31:0] m0s9_data_i;
  wire   [31:0] m0s10_data_i;
  wire   [31:0] m0s11_data_i;
  wire   [31:0] m0s12_data_i;
  wire   [31:0] m0s13_data_i;
  wire   [31:0] m0s14_data_i;
  wire   [31:0] m1s0_data_o;
  wire   [31:0] m1s0_addr;
  wire   [3:0] m1s0_sel;
  wire   [31:0] m2s0_data_o;
  wire   [31:0] m2s0_addr;
  wire   [3:0] m2s0_sel;
  wire   [31:0] m3s0_data_o;
  wire   [31:0] m3s0_addr;
  wire   [3:0] m3s0_sel;
  wire   [31:0] m4s0_data_o;
  wire   [31:0] m4s0_addr;
  wire   [3:0] m4s0_sel;
  wire   [31:0] m5s0_data_o;
  wire   [31:0] m5s0_addr;
  wire   [3:0] m5s0_sel;
  wire   [31:0] m6s0_data_o;
  wire   [31:0] m6s0_addr;
  wire   [3:0] m6s0_sel;
  wire   [31:0] m7s0_data_o;
  wire   [31:0] m7s0_addr;
  wire   [3:0] m7s0_sel;
  wire   [2:0] \s0/msel/gnt_p3 ;
  wire   [2:0] \s0/msel/gnt_p2 ;
  wire   [2:0] \s0/msel/gnt_p1 ;
  wire   [2:0] \s0/msel/gnt_p0 ;
  wire   [1:0] \s0/msel/pri_out ;
  wire   [2:0] \s1/msel/gnt_p3 ;
  wire   [2:0] \s1/msel/gnt_p2 ;
  wire   [2:0] \s1/msel/gnt_p1 ;
  wire   [2:0] \s1/msel/gnt_p0 ;
  wire   [1:0] \s1/msel/pri_out ;
  wire   [2:0] \s2/msel/gnt_p3 ;
  wire   [2:0] \s2/msel/gnt_p2 ;
  wire   [2:0] \s2/msel/gnt_p1 ;
  wire   [2:0] \s2/msel/gnt_p0 ;
  wire   [1:0] \s2/msel/pri_out ;
  wire   [2:0] \s3/msel/gnt_p3 ;
  wire   [2:0] \s3/msel/gnt_p2 ;
  wire   [2:0] \s3/msel/gnt_p1 ;
  wire   [2:0] \s3/msel/gnt_p0 ;
  wire   [1:0] \s3/msel/pri_out ;
  wire   [2:0] \s4/msel/gnt_p3 ;
  wire   [2:0] \s4/msel/gnt_p2 ;
  wire   [2:0] \s4/msel/gnt_p1 ;
  wire   [2:0] \s4/msel/gnt_p0 ;
  wire   [1:0] \s4/msel/pri_out ;
  wire   [2:0] \s5/msel/gnt_p3 ;
  wire   [2:0] \s5/msel/gnt_p2 ;
  wire   [2:0] \s5/msel/gnt_p1 ;
  wire   [2:0] \s5/msel/gnt_p0 ;
  wire   [1:0] \s5/msel/pri_out ;
  wire   [2:0] \s6/msel/gnt_p3 ;
  wire   [2:0] \s6/msel/gnt_p2 ;
  wire   [2:0] \s6/msel/gnt_p1 ;
  wire   [2:0] \s6/msel/gnt_p0 ;
  wire   [1:0] \s6/msel/pri_out ;
  wire   [2:0] \s7/msel/gnt_p3 ;
  wire   [2:0] \s7/msel/gnt_p2 ;
  wire   [2:0] \s7/msel/gnt_p1 ;
  wire   [2:0] \s7/msel/gnt_p0 ;
  wire   [1:0] \s7/msel/pri_out ;
  wire   [2:0] \s8/msel/gnt_p3 ;
  wire   [2:0] \s8/msel/gnt_p2 ;
  wire   [2:0] \s8/msel/gnt_p1 ;
  wire   [2:0] \s8/msel/gnt_p0 ;
  wire   [1:0] \s8/msel/pri_out ;
  wire   [2:0] \s9/msel/gnt_p3 ;
  wire   [2:0] \s9/msel/gnt_p2 ;
  wire   [2:0] \s9/msel/gnt_p1 ;
  wire   [2:0] \s9/msel/gnt_p0 ;
  wire   [1:0] \s9/msel/pri_out ;
  wire   [2:0] \s10/msel/gnt_p3 ;
  wire   [2:0] \s10/msel/gnt_p2 ;
  wire   [2:0] \s10/msel/gnt_p1 ;
  wire   [2:0] \s10/msel/gnt_p0 ;
  wire   [1:0] \s10/msel/pri_out ;
  wire   [2:0] \s11/msel/gnt_p3 ;
  wire   [2:0] \s11/msel/gnt_p2 ;
  wire   [2:0] \s11/msel/gnt_p1 ;
  wire   [2:0] \s11/msel/gnt_p0 ;
  wire   [1:0] \s11/msel/pri_out ;
  wire   [2:0] \s12/msel/gnt_p3 ;
  wire   [2:0] \s12/msel/gnt_p2 ;
  wire   [2:0] \s12/msel/gnt_p1 ;
  wire   [2:0] \s12/msel/gnt_p0 ;
  wire   [1:0] \s12/msel/pri_out ;
  wire   [2:0] \s13/msel/gnt_p3 ;
  wire   [2:0] \s13/msel/gnt_p2 ;
  wire   [2:0] \s13/msel/gnt_p1 ;
  wire   [2:0] \s13/msel/gnt_p0 ;
  wire   [1:0] \s13/msel/pri_out ;
  wire   [2:0] \s14/msel/gnt_p3 ;
  wire   [2:0] \s14/msel/gnt_p2 ;
  wire   [2:0] \s14/msel/gnt_p1 ;
  wire   [2:0] \s14/msel/gnt_p0 ;
  wire   [1:0] \s14/msel/pri_out ;
  wire   [2:0] \s15/msel/gnt_p3 ;
  wire   [2:0] \s15/msel/gnt_p2 ;
  wire   [2:0] \s15/msel/gnt_p1 ;
  wire   [2:0] \s15/msel/gnt_p0 ;
  wire   [1:0] \s15/msel/pri_out ;
  wire   [15:0] \rf/rf_dout ;
  assign m0s0_data_i[31] = s0_data_i[31];
  assign m0s0_data_i[30] = s0_data_i[30];
  assign m0s0_data_i[29] = s0_data_i[29];
  assign m0s0_data_i[28] = s0_data_i[28];
  assign m0s0_data_i[27] = s0_data_i[27];
  assign m0s0_data_i[26] = s0_data_i[26];
  assign m0s0_data_i[25] = s0_data_i[25];
  assign m0s0_data_i[24] = s0_data_i[24];
  assign m0s0_data_i[23] = s0_data_i[23];
  assign m0s0_data_i[22] = s0_data_i[22];
  assign m0s0_data_i[21] = s0_data_i[21];
  assign m0s0_data_i[20] = s0_data_i[20];
  assign m0s0_data_i[19] = s0_data_i[19];
  assign m0s0_data_i[18] = s0_data_i[18];
  assign m0s0_data_i[17] = s0_data_i[17];
  assign m0s0_data_i[16] = s0_data_i[16];
  assign m0s0_data_i[15] = s0_data_i[15];
  assign m0s0_data_i[14] = s0_data_i[14];
  assign m0s0_data_i[13] = s0_data_i[13];
  assign m0s0_data_i[12] = s0_data_i[12];
  assign m0s0_data_i[11] = s0_data_i[11];
  assign m0s0_data_i[10] = s0_data_i[10];
  assign m0s0_data_i[9] = s0_data_i[9];
  assign m0s0_data_i[8] = s0_data_i[8];
  assign m0s0_data_i[7] = s0_data_i[7];
  assign m0s0_data_i[6] = s0_data_i[6];
  assign m0s0_data_i[5] = s0_data_i[5];
  assign m0s0_data_i[4] = s0_data_i[4];
  assign m0s0_data_i[3] = s0_data_i[3];
  assign m0s0_data_i[2] = s0_data_i[2];
  assign m0s0_data_i[1] = s0_data_i[1];
  assign m0s0_data_i[0] = s0_data_i[0];
  assign m0s0_data_o[31] = m0_data_i[31];
  assign m0s0_data_o[30] = m0_data_i[30];
  assign m0s0_data_o[29] = m0_data_i[29];
  assign m0s0_data_o[28] = m0_data_i[28];
  assign m0s0_data_o[27] = m0_data_i[27];
  assign m0s0_data_o[26] = m0_data_i[26];
  assign m0s0_data_o[25] = m0_data_i[25];
  assign m0s0_data_o[24] = m0_data_i[24];
  assign m0s0_data_o[23] = m0_data_i[23];
  assign m0s0_data_o[22] = m0_data_i[22];
  assign m0s0_data_o[21] = m0_data_i[21];
  assign m0s0_data_o[20] = m0_data_i[20];
  assign m0s0_data_o[19] = m0_data_i[19];
  assign m0s0_data_o[18] = m0_data_i[18];
  assign m0s0_data_o[17] = m0_data_i[17];
  assign m0s0_data_o[16] = m0_data_i[16];
  assign m0s0_data_o[15] = m0_data_i[15];
  assign m0s0_data_o[14] = m0_data_i[14];
  assign m0s0_data_o[13] = m0_data_i[13];
  assign m0s0_data_o[12] = m0_data_i[12];
  assign m0s0_data_o[11] = m0_data_i[11];
  assign m0s0_data_o[10] = m0_data_i[10];
  assign m0s0_data_o[9] = m0_data_i[9];
  assign m0s0_data_o[8] = m0_data_i[8];
  assign m0s0_data_o[7] = m0_data_i[7];
  assign m0s0_data_o[6] = m0_data_i[6];
  assign m0s0_data_o[5] = m0_data_i[5];
  assign m0s0_data_o[4] = m0_data_i[4];
  assign m0s0_data_o[3] = m0_data_i[3];
  assign m0s0_data_o[2] = m0_data_i[2];
  assign m0s0_data_o[1] = m0_data_i[1];
  assign m0s0_data_o[0] = m0_data_i[0];
  assign m0s0_addr[31] = m0_addr_i[31];
  assign m0s0_addr[30] = m0_addr_i[30];
  assign m0s0_addr[29] = m0_addr_i[29];
  assign m0s0_addr[28] = m0_addr_i[28];
  assign m0s0_addr[27] = m0_addr_i[27];
  assign m0s0_addr[26] = m0_addr_i[26];
  assign m0s0_addr[25] = m0_addr_i[25];
  assign m0s0_addr[24] = m0_addr_i[24];
  assign m0s0_addr[23] = m0_addr_i[23];
  assign m0s0_addr[22] = m0_addr_i[22];
  assign m0s0_addr[21] = m0_addr_i[21];
  assign m0s0_addr[20] = m0_addr_i[20];
  assign m0s0_addr[19] = m0_addr_i[19];
  assign m0s0_addr[18] = m0_addr_i[18];
  assign m0s0_addr[17] = m0_addr_i[17];
  assign m0s0_addr[16] = m0_addr_i[16];
  assign m0s0_addr[15] = m0_addr_i[15];
  assign m0s0_addr[14] = m0_addr_i[14];
  assign m0s0_addr[13] = m0_addr_i[13];
  assign m0s0_addr[12] = m0_addr_i[12];
  assign m0s0_addr[11] = m0_addr_i[11];
  assign m0s0_addr[10] = m0_addr_i[10];
  assign m0s0_addr[9] = m0_addr_i[9];
  assign m0s0_addr[8] = m0_addr_i[8];
  assign m0s0_addr[7] = m0_addr_i[7];
  assign m0s0_addr[6] = m0_addr_i[6];
  assign m0s0_addr[5] = m0_addr_i[5];
  assign m0s0_addr[4] = m0_addr_i[4];
  assign m0s0_addr[3] = m0_addr_i[3];
  assign m0s0_addr[2] = m0_addr_i[2];
  assign m0s0_addr[1] = m0_addr_i[1];
  assign m0s0_addr[0] = m0_addr_i[0];
  assign m0s0_sel[3] = m0_sel_i[3];
  assign m0s0_sel[2] = m0_sel_i[2];
  assign m0s0_sel[1] = m0_sel_i[1];
  assign m0s0_sel[0] = m0_sel_i[0];
  assign m0s0_we = m0_we_i;
  assign m0s1_data_i[31] = s1_data_i[31];
  assign m0s1_data_i[30] = s1_data_i[30];
  assign m0s1_data_i[29] = s1_data_i[29];
  assign m0s1_data_i[28] = s1_data_i[28];
  assign m0s1_data_i[27] = s1_data_i[27];
  assign m0s1_data_i[26] = s1_data_i[26];
  assign m0s1_data_i[25] = s1_data_i[25];
  assign m0s1_data_i[24] = s1_data_i[24];
  assign m0s1_data_i[23] = s1_data_i[23];
  assign m0s1_data_i[22] = s1_data_i[22];
  assign m0s1_data_i[21] = s1_data_i[21];
  assign m0s1_data_i[20] = s1_data_i[20];
  assign m0s1_data_i[19] = s1_data_i[19];
  assign m0s1_data_i[18] = s1_data_i[18];
  assign m0s1_data_i[17] = s1_data_i[17];
  assign m0s1_data_i[16] = s1_data_i[16];
  assign m0s1_data_i[15] = s1_data_i[15];
  assign m0s1_data_i[14] = s1_data_i[14];
  assign m0s1_data_i[13] = s1_data_i[13];
  assign m0s1_data_i[12] = s1_data_i[12];
  assign m0s1_data_i[11] = s1_data_i[11];
  assign m0s1_data_i[10] = s1_data_i[10];
  assign m0s1_data_i[9] = s1_data_i[9];
  assign m0s1_data_i[8] = s1_data_i[8];
  assign m0s1_data_i[7] = s1_data_i[7];
  assign m0s1_data_i[6] = s1_data_i[6];
  assign m0s1_data_i[5] = s1_data_i[5];
  assign m0s1_data_i[4] = s1_data_i[4];
  assign m0s1_data_i[3] = s1_data_i[3];
  assign m0s1_data_i[2] = s1_data_i[2];
  assign m0s1_data_i[1] = s1_data_i[1];
  assign m0s1_data_i[0] = s1_data_i[0];
  assign m0s2_data_i[31] = s2_data_i[31];
  assign m0s2_data_i[30] = s2_data_i[30];
  assign m0s2_data_i[29] = s2_data_i[29];
  assign m0s2_data_i[28] = s2_data_i[28];
  assign m0s2_data_i[27] = s2_data_i[27];
  assign m0s2_data_i[26] = s2_data_i[26];
  assign m0s2_data_i[25] = s2_data_i[25];
  assign m0s2_data_i[24] = s2_data_i[24];
  assign m0s2_data_i[23] = s2_data_i[23];
  assign m0s2_data_i[22] = s2_data_i[22];
  assign m0s2_data_i[21] = s2_data_i[21];
  assign m0s2_data_i[20] = s2_data_i[20];
  assign m0s2_data_i[19] = s2_data_i[19];
  assign m0s2_data_i[18] = s2_data_i[18];
  assign m0s2_data_i[17] = s2_data_i[17];
  assign m0s2_data_i[16] = s2_data_i[16];
  assign m0s2_data_i[15] = s2_data_i[15];
  assign m0s2_data_i[14] = s2_data_i[14];
  assign m0s2_data_i[13] = s2_data_i[13];
  assign m0s2_data_i[12] = s2_data_i[12];
  assign m0s2_data_i[11] = s2_data_i[11];
  assign m0s2_data_i[10] = s2_data_i[10];
  assign m0s2_data_i[9] = s2_data_i[9];
  assign m0s2_data_i[8] = s2_data_i[8];
  assign m0s2_data_i[7] = s2_data_i[7];
  assign m0s2_data_i[6] = s2_data_i[6];
  assign m0s2_data_i[5] = s2_data_i[5];
  assign m0s2_data_i[4] = s2_data_i[4];
  assign m0s2_data_i[3] = s2_data_i[3];
  assign m0s2_data_i[2] = s2_data_i[2];
  assign m0s2_data_i[1] = s2_data_i[1];
  assign m0s2_data_i[0] = s2_data_i[0];
  assign m0s3_data_i[31] = s3_data_i[31];
  assign m0s3_data_i[30] = s3_data_i[30];
  assign m0s3_data_i[29] = s3_data_i[29];
  assign m0s3_data_i[28] = s3_data_i[28];
  assign m0s3_data_i[27] = s3_data_i[27];
  assign m0s3_data_i[26] = s3_data_i[26];
  assign m0s3_data_i[25] = s3_data_i[25];
  assign m0s3_data_i[24] = s3_data_i[24];
  assign m0s3_data_i[23] = s3_data_i[23];
  assign m0s3_data_i[22] = s3_data_i[22];
  assign m0s3_data_i[21] = s3_data_i[21];
  assign m0s3_data_i[20] = s3_data_i[20];
  assign m0s3_data_i[19] = s3_data_i[19];
  assign m0s3_data_i[18] = s3_data_i[18];
  assign m0s3_data_i[17] = s3_data_i[17];
  assign m0s3_data_i[16] = s3_data_i[16];
  assign m0s3_data_i[15] = s3_data_i[15];
  assign m0s3_data_i[14] = s3_data_i[14];
  assign m0s3_data_i[13] = s3_data_i[13];
  assign m0s3_data_i[12] = s3_data_i[12];
  assign m0s3_data_i[11] = s3_data_i[11];
  assign m0s3_data_i[10] = s3_data_i[10];
  assign m0s3_data_i[9] = s3_data_i[9];
  assign m0s3_data_i[8] = s3_data_i[8];
  assign m0s3_data_i[7] = s3_data_i[7];
  assign m0s3_data_i[6] = s3_data_i[6];
  assign m0s3_data_i[5] = s3_data_i[5];
  assign m0s3_data_i[4] = s3_data_i[4];
  assign m0s3_data_i[3] = s3_data_i[3];
  assign m0s3_data_i[2] = s3_data_i[2];
  assign m0s3_data_i[1] = s3_data_i[1];
  assign m0s3_data_i[0] = s3_data_i[0];
  assign m0s4_data_i[31] = s4_data_i[31];
  assign m0s4_data_i[30] = s4_data_i[30];
  assign m0s4_data_i[29] = s4_data_i[29];
  assign m0s4_data_i[28] = s4_data_i[28];
  assign m0s4_data_i[27] = s4_data_i[27];
  assign m0s4_data_i[26] = s4_data_i[26];
  assign m0s4_data_i[25] = s4_data_i[25];
  assign m0s4_data_i[24] = s4_data_i[24];
  assign m0s4_data_i[23] = s4_data_i[23];
  assign m0s4_data_i[22] = s4_data_i[22];
  assign m0s4_data_i[21] = s4_data_i[21];
  assign m0s4_data_i[20] = s4_data_i[20];
  assign m0s4_data_i[19] = s4_data_i[19];
  assign m0s4_data_i[18] = s4_data_i[18];
  assign m0s4_data_i[17] = s4_data_i[17];
  assign m0s4_data_i[16] = s4_data_i[16];
  assign m0s4_data_i[15] = s4_data_i[15];
  assign m0s4_data_i[14] = s4_data_i[14];
  assign m0s4_data_i[13] = s4_data_i[13];
  assign m0s4_data_i[12] = s4_data_i[12];
  assign m0s4_data_i[11] = s4_data_i[11];
  assign m0s4_data_i[10] = s4_data_i[10];
  assign m0s4_data_i[9] = s4_data_i[9];
  assign m0s4_data_i[8] = s4_data_i[8];
  assign m0s4_data_i[7] = s4_data_i[7];
  assign m0s4_data_i[6] = s4_data_i[6];
  assign m0s4_data_i[5] = s4_data_i[5];
  assign m0s4_data_i[4] = s4_data_i[4];
  assign m0s4_data_i[3] = s4_data_i[3];
  assign m0s4_data_i[2] = s4_data_i[2];
  assign m0s4_data_i[1] = s4_data_i[1];
  assign m0s4_data_i[0] = s4_data_i[0];
  assign m0s5_data_i[31] = s5_data_i[31];
  assign m0s5_data_i[30] = s5_data_i[30];
  assign m0s5_data_i[29] = s5_data_i[29];
  assign m0s5_data_i[28] = s5_data_i[28];
  assign m0s5_data_i[27] = s5_data_i[27];
  assign m0s5_data_i[26] = s5_data_i[26];
  assign m0s5_data_i[25] = s5_data_i[25];
  assign m0s5_data_i[24] = s5_data_i[24];
  assign m0s5_data_i[23] = s5_data_i[23];
  assign m0s5_data_i[22] = s5_data_i[22];
  assign m0s5_data_i[21] = s5_data_i[21];
  assign m0s5_data_i[20] = s5_data_i[20];
  assign m0s5_data_i[19] = s5_data_i[19];
  assign m0s5_data_i[18] = s5_data_i[18];
  assign m0s5_data_i[17] = s5_data_i[17];
  assign m0s5_data_i[16] = s5_data_i[16];
  assign m0s5_data_i[15] = s5_data_i[15];
  assign m0s5_data_i[14] = s5_data_i[14];
  assign m0s5_data_i[13] = s5_data_i[13];
  assign m0s5_data_i[12] = s5_data_i[12];
  assign m0s5_data_i[11] = s5_data_i[11];
  assign m0s5_data_i[10] = s5_data_i[10];
  assign m0s5_data_i[9] = s5_data_i[9];
  assign m0s5_data_i[8] = s5_data_i[8];
  assign m0s5_data_i[7] = s5_data_i[7];
  assign m0s5_data_i[6] = s5_data_i[6];
  assign m0s5_data_i[5] = s5_data_i[5];
  assign m0s5_data_i[4] = s5_data_i[4];
  assign m0s5_data_i[3] = s5_data_i[3];
  assign m0s5_data_i[2] = s5_data_i[2];
  assign m0s5_data_i[1] = s5_data_i[1];
  assign m0s5_data_i[0] = s5_data_i[0];
  assign m0s6_data_i[31] = s6_data_i[31];
  assign m0s6_data_i[30] = s6_data_i[30];
  assign m0s6_data_i[29] = s6_data_i[29];
  assign m0s6_data_i[28] = s6_data_i[28];
  assign m0s6_data_i[27] = s6_data_i[27];
  assign m0s6_data_i[26] = s6_data_i[26];
  assign m0s6_data_i[25] = s6_data_i[25];
  assign m0s6_data_i[24] = s6_data_i[24];
  assign m0s6_data_i[23] = s6_data_i[23];
  assign m0s6_data_i[22] = s6_data_i[22];
  assign m0s6_data_i[21] = s6_data_i[21];
  assign m0s6_data_i[20] = s6_data_i[20];
  assign m0s6_data_i[19] = s6_data_i[19];
  assign m0s6_data_i[18] = s6_data_i[18];
  assign m0s6_data_i[17] = s6_data_i[17];
  assign m0s6_data_i[16] = s6_data_i[16];
  assign m0s6_data_i[15] = s6_data_i[15];
  assign m0s6_data_i[14] = s6_data_i[14];
  assign m0s6_data_i[13] = s6_data_i[13];
  assign m0s6_data_i[12] = s6_data_i[12];
  assign m0s6_data_i[11] = s6_data_i[11];
  assign m0s6_data_i[10] = s6_data_i[10];
  assign m0s6_data_i[9] = s6_data_i[9];
  assign m0s6_data_i[8] = s6_data_i[8];
  assign m0s6_data_i[7] = s6_data_i[7];
  assign m0s6_data_i[6] = s6_data_i[6];
  assign m0s6_data_i[5] = s6_data_i[5];
  assign m0s6_data_i[4] = s6_data_i[4];
  assign m0s6_data_i[3] = s6_data_i[3];
  assign m0s6_data_i[2] = s6_data_i[2];
  assign m0s6_data_i[1] = s6_data_i[1];
  assign m0s6_data_i[0] = s6_data_i[0];
  assign m0s7_data_i[31] = s7_data_i[31];
  assign m0s7_data_i[30] = s7_data_i[30];
  assign m0s7_data_i[29] = s7_data_i[29];
  assign m0s7_data_i[28] = s7_data_i[28];
  assign m0s7_data_i[27] = s7_data_i[27];
  assign m0s7_data_i[26] = s7_data_i[26];
  assign m0s7_data_i[25] = s7_data_i[25];
  assign m0s7_data_i[24] = s7_data_i[24];
  assign m0s7_data_i[23] = s7_data_i[23];
  assign m0s7_data_i[22] = s7_data_i[22];
  assign m0s7_data_i[21] = s7_data_i[21];
  assign m0s7_data_i[20] = s7_data_i[20];
  assign m0s7_data_i[19] = s7_data_i[19];
  assign m0s7_data_i[18] = s7_data_i[18];
  assign m0s7_data_i[17] = s7_data_i[17];
  assign m0s7_data_i[16] = s7_data_i[16];
  assign m0s7_data_i[15] = s7_data_i[15];
  assign m0s7_data_i[14] = s7_data_i[14];
  assign m0s7_data_i[13] = s7_data_i[13];
  assign m0s7_data_i[12] = s7_data_i[12];
  assign m0s7_data_i[11] = s7_data_i[11];
  assign m0s7_data_i[10] = s7_data_i[10];
  assign m0s7_data_i[9] = s7_data_i[9];
  assign m0s7_data_i[8] = s7_data_i[8];
  assign m0s7_data_i[7] = s7_data_i[7];
  assign m0s7_data_i[6] = s7_data_i[6];
  assign m0s7_data_i[5] = s7_data_i[5];
  assign m0s7_data_i[4] = s7_data_i[4];
  assign m0s7_data_i[3] = s7_data_i[3];
  assign m0s7_data_i[2] = s7_data_i[2];
  assign m0s7_data_i[1] = s7_data_i[1];
  assign m0s7_data_i[0] = s7_data_i[0];
  assign m0s8_data_i[31] = s8_data_i[31];
  assign m0s8_data_i[30] = s8_data_i[30];
  assign m0s8_data_i[29] = s8_data_i[29];
  assign m0s8_data_i[28] = s8_data_i[28];
  assign m0s8_data_i[27] = s8_data_i[27];
  assign m0s8_data_i[26] = s8_data_i[26];
  assign m0s8_data_i[25] = s8_data_i[25];
  assign m0s8_data_i[24] = s8_data_i[24];
  assign m0s8_data_i[23] = s8_data_i[23];
  assign m0s8_data_i[22] = s8_data_i[22];
  assign m0s8_data_i[21] = s8_data_i[21];
  assign m0s8_data_i[20] = s8_data_i[20];
  assign m0s8_data_i[19] = s8_data_i[19];
  assign m0s8_data_i[18] = s8_data_i[18];
  assign m0s8_data_i[17] = s8_data_i[17];
  assign m0s8_data_i[16] = s8_data_i[16];
  assign m0s8_data_i[15] = s8_data_i[15];
  assign m0s8_data_i[14] = s8_data_i[14];
  assign m0s8_data_i[13] = s8_data_i[13];
  assign m0s8_data_i[12] = s8_data_i[12];
  assign m0s8_data_i[11] = s8_data_i[11];
  assign m0s8_data_i[10] = s8_data_i[10];
  assign m0s8_data_i[9] = s8_data_i[9];
  assign m0s8_data_i[8] = s8_data_i[8];
  assign m0s8_data_i[7] = s8_data_i[7];
  assign m0s8_data_i[6] = s8_data_i[6];
  assign m0s8_data_i[5] = s8_data_i[5];
  assign m0s8_data_i[4] = s8_data_i[4];
  assign m0s8_data_i[3] = s8_data_i[3];
  assign m0s8_data_i[2] = s8_data_i[2];
  assign m0s8_data_i[1] = s8_data_i[1];
  assign m0s8_data_i[0] = s8_data_i[0];
  assign m0s9_data_i[31] = s9_data_i[31];
  assign m0s9_data_i[30] = s9_data_i[30];
  assign m0s9_data_i[29] = s9_data_i[29];
  assign m0s9_data_i[28] = s9_data_i[28];
  assign m0s9_data_i[27] = s9_data_i[27];
  assign m0s9_data_i[26] = s9_data_i[26];
  assign m0s9_data_i[25] = s9_data_i[25];
  assign m0s9_data_i[24] = s9_data_i[24];
  assign m0s9_data_i[23] = s9_data_i[23];
  assign m0s9_data_i[22] = s9_data_i[22];
  assign m0s9_data_i[21] = s9_data_i[21];
  assign m0s9_data_i[20] = s9_data_i[20];
  assign m0s9_data_i[19] = s9_data_i[19];
  assign m0s9_data_i[18] = s9_data_i[18];
  assign m0s9_data_i[17] = s9_data_i[17];
  assign m0s9_data_i[16] = s9_data_i[16];
  assign m0s9_data_i[15] = s9_data_i[15];
  assign m0s9_data_i[14] = s9_data_i[14];
  assign m0s9_data_i[13] = s9_data_i[13];
  assign m0s9_data_i[12] = s9_data_i[12];
  assign m0s9_data_i[11] = s9_data_i[11];
  assign m0s9_data_i[10] = s9_data_i[10];
  assign m0s9_data_i[9] = s9_data_i[9];
  assign m0s9_data_i[8] = s9_data_i[8];
  assign m0s9_data_i[7] = s9_data_i[7];
  assign m0s9_data_i[6] = s9_data_i[6];
  assign m0s9_data_i[5] = s9_data_i[5];
  assign m0s9_data_i[4] = s9_data_i[4];
  assign m0s9_data_i[3] = s9_data_i[3];
  assign m0s9_data_i[2] = s9_data_i[2];
  assign m0s9_data_i[1] = s9_data_i[1];
  assign m0s9_data_i[0] = s9_data_i[0];
  assign m0s10_data_i[31] = s10_data_i[31];
  assign m0s10_data_i[30] = s10_data_i[30];
  assign m0s10_data_i[29] = s10_data_i[29];
  assign m0s10_data_i[28] = s10_data_i[28];
  assign m0s10_data_i[27] = s10_data_i[27];
  assign m0s10_data_i[26] = s10_data_i[26];
  assign m0s10_data_i[25] = s10_data_i[25];
  assign m0s10_data_i[24] = s10_data_i[24];
  assign m0s10_data_i[23] = s10_data_i[23];
  assign m0s10_data_i[22] = s10_data_i[22];
  assign m0s10_data_i[21] = s10_data_i[21];
  assign m0s10_data_i[20] = s10_data_i[20];
  assign m0s10_data_i[19] = s10_data_i[19];
  assign m0s10_data_i[18] = s10_data_i[18];
  assign m0s10_data_i[17] = s10_data_i[17];
  assign m0s10_data_i[16] = s10_data_i[16];
  assign m0s10_data_i[15] = s10_data_i[15];
  assign m0s10_data_i[14] = s10_data_i[14];
  assign m0s10_data_i[13] = s10_data_i[13];
  assign m0s10_data_i[12] = s10_data_i[12];
  assign m0s10_data_i[11] = s10_data_i[11];
  assign m0s10_data_i[10] = s10_data_i[10];
  assign m0s10_data_i[9] = s10_data_i[9];
  assign m0s10_data_i[8] = s10_data_i[8];
  assign m0s10_data_i[7] = s10_data_i[7];
  assign m0s10_data_i[6] = s10_data_i[6];
  assign m0s10_data_i[5] = s10_data_i[5];
  assign m0s10_data_i[4] = s10_data_i[4];
  assign m0s10_data_i[3] = s10_data_i[3];
  assign m0s10_data_i[2] = s10_data_i[2];
  assign m0s10_data_i[1] = s10_data_i[1];
  assign m0s10_data_i[0] = s10_data_i[0];
  assign m0s11_data_i[31] = s11_data_i[31];
  assign m0s11_data_i[30] = s11_data_i[30];
  assign m0s11_data_i[29] = s11_data_i[29];
  assign m0s11_data_i[28] = s11_data_i[28];
  assign m0s11_data_i[27] = s11_data_i[27];
  assign m0s11_data_i[26] = s11_data_i[26];
  assign m0s11_data_i[25] = s11_data_i[25];
  assign m0s11_data_i[24] = s11_data_i[24];
  assign m0s11_data_i[23] = s11_data_i[23];
  assign m0s11_data_i[22] = s11_data_i[22];
  assign m0s11_data_i[21] = s11_data_i[21];
  assign m0s11_data_i[20] = s11_data_i[20];
  assign m0s11_data_i[19] = s11_data_i[19];
  assign m0s11_data_i[18] = s11_data_i[18];
  assign m0s11_data_i[17] = s11_data_i[17];
  assign m0s11_data_i[16] = s11_data_i[16];
  assign m0s11_data_i[15] = s11_data_i[15];
  assign m0s11_data_i[14] = s11_data_i[14];
  assign m0s11_data_i[13] = s11_data_i[13];
  assign m0s11_data_i[12] = s11_data_i[12];
  assign m0s11_data_i[11] = s11_data_i[11];
  assign m0s11_data_i[10] = s11_data_i[10];
  assign m0s11_data_i[9] = s11_data_i[9];
  assign m0s11_data_i[8] = s11_data_i[8];
  assign m0s11_data_i[7] = s11_data_i[7];
  assign m0s11_data_i[6] = s11_data_i[6];
  assign m0s11_data_i[5] = s11_data_i[5];
  assign m0s11_data_i[4] = s11_data_i[4];
  assign m0s11_data_i[3] = s11_data_i[3];
  assign m0s11_data_i[2] = s11_data_i[2];
  assign m0s11_data_i[1] = s11_data_i[1];
  assign m0s11_data_i[0] = s11_data_i[0];
  assign m0s12_data_i[31] = s12_data_i[31];
  assign m0s12_data_i[30] = s12_data_i[30];
  assign m0s12_data_i[29] = s12_data_i[29];
  assign m0s12_data_i[28] = s12_data_i[28];
  assign m0s12_data_i[27] = s12_data_i[27];
  assign m0s12_data_i[26] = s12_data_i[26];
  assign m0s12_data_i[25] = s12_data_i[25];
  assign m0s12_data_i[24] = s12_data_i[24];
  assign m0s12_data_i[23] = s12_data_i[23];
  assign m0s12_data_i[22] = s12_data_i[22];
  assign m0s12_data_i[21] = s12_data_i[21];
  assign m0s12_data_i[20] = s12_data_i[20];
  assign m0s12_data_i[19] = s12_data_i[19];
  assign m0s12_data_i[18] = s12_data_i[18];
  assign m0s12_data_i[17] = s12_data_i[17];
  assign m0s12_data_i[16] = s12_data_i[16];
  assign m0s12_data_i[15] = s12_data_i[15];
  assign m0s12_data_i[14] = s12_data_i[14];
  assign m0s12_data_i[13] = s12_data_i[13];
  assign m0s12_data_i[12] = s12_data_i[12];
  assign m0s12_data_i[11] = s12_data_i[11];
  assign m0s12_data_i[10] = s12_data_i[10];
  assign m0s12_data_i[9] = s12_data_i[9];
  assign m0s12_data_i[8] = s12_data_i[8];
  assign m0s12_data_i[7] = s12_data_i[7];
  assign m0s12_data_i[6] = s12_data_i[6];
  assign m0s12_data_i[5] = s12_data_i[5];
  assign m0s12_data_i[4] = s12_data_i[4];
  assign m0s12_data_i[3] = s12_data_i[3];
  assign m0s12_data_i[2] = s12_data_i[2];
  assign m0s12_data_i[1] = s12_data_i[1];
  assign m0s12_data_i[0] = s12_data_i[0];
  assign m0s13_data_i[31] = s13_data_i[31];
  assign m0s13_data_i[30] = s13_data_i[30];
  assign m0s13_data_i[29] = s13_data_i[29];
  assign m0s13_data_i[28] = s13_data_i[28];
  assign m0s13_data_i[27] = s13_data_i[27];
  assign m0s13_data_i[26] = s13_data_i[26];
  assign m0s13_data_i[25] = s13_data_i[25];
  assign m0s13_data_i[24] = s13_data_i[24];
  assign m0s13_data_i[23] = s13_data_i[23];
  assign m0s13_data_i[22] = s13_data_i[22];
  assign m0s13_data_i[21] = s13_data_i[21];
  assign m0s13_data_i[20] = s13_data_i[20];
  assign m0s13_data_i[19] = s13_data_i[19];
  assign m0s13_data_i[18] = s13_data_i[18];
  assign m0s13_data_i[17] = s13_data_i[17];
  assign m0s13_data_i[16] = s13_data_i[16];
  assign m0s13_data_i[15] = s13_data_i[15];
  assign m0s13_data_i[14] = s13_data_i[14];
  assign m0s13_data_i[13] = s13_data_i[13];
  assign m0s13_data_i[12] = s13_data_i[12];
  assign m0s13_data_i[11] = s13_data_i[11];
  assign m0s13_data_i[10] = s13_data_i[10];
  assign m0s13_data_i[9] = s13_data_i[9];
  assign m0s13_data_i[8] = s13_data_i[8];
  assign m0s13_data_i[7] = s13_data_i[7];
  assign m0s13_data_i[6] = s13_data_i[6];
  assign m0s13_data_i[5] = s13_data_i[5];
  assign m0s13_data_i[4] = s13_data_i[4];
  assign m0s13_data_i[3] = s13_data_i[3];
  assign m0s13_data_i[2] = s13_data_i[2];
  assign m0s13_data_i[1] = s13_data_i[1];
  assign m0s13_data_i[0] = s13_data_i[0];
  assign m0s14_data_i[31] = s14_data_i[31];
  assign m0s14_data_i[30] = s14_data_i[30];
  assign m0s14_data_i[29] = s14_data_i[29];
  assign m0s14_data_i[28] = s14_data_i[28];
  assign m0s14_data_i[27] = s14_data_i[27];
  assign m0s14_data_i[26] = s14_data_i[26];
  assign m0s14_data_i[25] = s14_data_i[25];
  assign m0s14_data_i[24] = s14_data_i[24];
  assign m0s14_data_i[23] = s14_data_i[23];
  assign m0s14_data_i[22] = s14_data_i[22];
  assign m0s14_data_i[21] = s14_data_i[21];
  assign m0s14_data_i[20] = s14_data_i[20];
  assign m0s14_data_i[19] = s14_data_i[19];
  assign m0s14_data_i[18] = s14_data_i[18];
  assign m0s14_data_i[17] = s14_data_i[17];
  assign m0s14_data_i[16] = s14_data_i[16];
  assign m0s14_data_i[15] = s14_data_i[15];
  assign m0s14_data_i[14] = s14_data_i[14];
  assign m0s14_data_i[13] = s14_data_i[13];
  assign m0s14_data_i[12] = s14_data_i[12];
  assign m0s14_data_i[11] = s14_data_i[11];
  assign m0s14_data_i[10] = s14_data_i[10];
  assign m0s14_data_i[9] = s14_data_i[9];
  assign m0s14_data_i[8] = s14_data_i[8];
  assign m0s14_data_i[7] = s14_data_i[7];
  assign m0s14_data_i[6] = s14_data_i[6];
  assign m0s14_data_i[5] = s14_data_i[5];
  assign m0s14_data_i[4] = s14_data_i[4];
  assign m0s14_data_i[3] = s14_data_i[3];
  assign m0s14_data_i[2] = s14_data_i[2];
  assign m0s14_data_i[1] = s14_data_i[1];
  assign m0s14_data_i[0] = s14_data_i[0];
  assign m1s0_data_o[31] = m1_data_i[31];
  assign m1s0_data_o[30] = m1_data_i[30];
  assign m1s0_data_o[29] = m1_data_i[29];
  assign m1s0_data_o[28] = m1_data_i[28];
  assign m1s0_data_o[27] = m1_data_i[27];
  assign m1s0_data_o[26] = m1_data_i[26];
  assign m1s0_data_o[25] = m1_data_i[25];
  assign m1s0_data_o[24] = m1_data_i[24];
  assign m1s0_data_o[23] = m1_data_i[23];
  assign m1s0_data_o[22] = m1_data_i[22];
  assign m1s0_data_o[21] = m1_data_i[21];
  assign m1s0_data_o[20] = m1_data_i[20];
  assign m1s0_data_o[19] = m1_data_i[19];
  assign m1s0_data_o[18] = m1_data_i[18];
  assign m1s0_data_o[17] = m1_data_i[17];
  assign m1s0_data_o[16] = m1_data_i[16];
  assign m1s0_data_o[15] = m1_data_i[15];
  assign m1s0_data_o[14] = m1_data_i[14];
  assign m1s0_data_o[13] = m1_data_i[13];
  assign m1s0_data_o[12] = m1_data_i[12];
  assign m1s0_data_o[11] = m1_data_i[11];
  assign m1s0_data_o[10] = m1_data_i[10];
  assign m1s0_data_o[9] = m1_data_i[9];
  assign m1s0_data_o[8] = m1_data_i[8];
  assign m1s0_data_o[7] = m1_data_i[7];
  assign m1s0_data_o[6] = m1_data_i[6];
  assign m1s0_data_o[5] = m1_data_i[5];
  assign m1s0_data_o[4] = m1_data_i[4];
  assign m1s0_data_o[3] = m1_data_i[3];
  assign m1s0_data_o[2] = m1_data_i[2];
  assign m1s0_data_o[1] = m1_data_i[1];
  assign m1s0_data_o[0] = m1_data_i[0];
  assign m1s0_addr[31] = m1_addr_i[31];
  assign m1s0_addr[30] = m1_addr_i[30];
  assign m1s0_addr[29] = m1_addr_i[29];
  assign m1s0_addr[28] = m1_addr_i[28];
  assign m1s0_addr[27] = m1_addr_i[27];
  assign m1s0_addr[26] = m1_addr_i[26];
  assign m1s0_addr[25] = m1_addr_i[25];
  assign m1s0_addr[24] = m1_addr_i[24];
  assign m1s0_addr[23] = m1_addr_i[23];
  assign m1s0_addr[22] = m1_addr_i[22];
  assign m1s0_addr[21] = m1_addr_i[21];
  assign m1s0_addr[20] = m1_addr_i[20];
  assign m1s0_addr[19] = m1_addr_i[19];
  assign m1s0_addr[18] = m1_addr_i[18];
  assign m1s0_addr[17] = m1_addr_i[17];
  assign m1s0_addr[16] = m1_addr_i[16];
  assign m1s0_addr[15] = m1_addr_i[15];
  assign m1s0_addr[14] = m1_addr_i[14];
  assign m1s0_addr[13] = m1_addr_i[13];
  assign m1s0_addr[12] = m1_addr_i[12];
  assign m1s0_addr[11] = m1_addr_i[11];
  assign m1s0_addr[10] = m1_addr_i[10];
  assign m1s0_addr[9] = m1_addr_i[9];
  assign m1s0_addr[8] = m1_addr_i[8];
  assign m1s0_addr[7] = m1_addr_i[7];
  assign m1s0_addr[6] = m1_addr_i[6];
  assign m1s0_addr[5] = m1_addr_i[5];
  assign m1s0_addr[4] = m1_addr_i[4];
  assign m1s0_addr[3] = m1_addr_i[3];
  assign m1s0_addr[2] = m1_addr_i[2];
  assign m1s0_addr[1] = m1_addr_i[1];
  assign m1s0_addr[0] = m1_addr_i[0];
  assign m1s0_sel[3] = m1_sel_i[3];
  assign m1s0_sel[2] = m1_sel_i[2];
  assign m1s0_sel[1] = m1_sel_i[1];
  assign m1s0_sel[0] = m1_sel_i[0];
  assign m1s0_we = m1_we_i;
  assign m2s0_data_o[31] = m2_data_i[31];
  assign m2s0_data_o[30] = m2_data_i[30];
  assign m2s0_data_o[29] = m2_data_i[29];
  assign m2s0_data_o[28] = m2_data_i[28];
  assign m2s0_data_o[27] = m2_data_i[27];
  assign m2s0_data_o[26] = m2_data_i[26];
  assign m2s0_data_o[25] = m2_data_i[25];
  assign m2s0_data_o[24] = m2_data_i[24];
  assign m2s0_data_o[23] = m2_data_i[23];
  assign m2s0_data_o[22] = m2_data_i[22];
  assign m2s0_data_o[21] = m2_data_i[21];
  assign m2s0_data_o[20] = m2_data_i[20];
  assign m2s0_data_o[19] = m2_data_i[19];
  assign m2s0_data_o[18] = m2_data_i[18];
  assign m2s0_data_o[17] = m2_data_i[17];
  assign m2s0_data_o[16] = m2_data_i[16];
  assign m2s0_data_o[15] = m2_data_i[15];
  assign m2s0_data_o[14] = m2_data_i[14];
  assign m2s0_data_o[13] = m2_data_i[13];
  assign m2s0_data_o[12] = m2_data_i[12];
  assign m2s0_data_o[11] = m2_data_i[11];
  assign m2s0_data_o[10] = m2_data_i[10];
  assign m2s0_data_o[9] = m2_data_i[9];
  assign m2s0_data_o[8] = m2_data_i[8];
  assign m2s0_data_o[7] = m2_data_i[7];
  assign m2s0_data_o[6] = m2_data_i[6];
  assign m2s0_data_o[5] = m2_data_i[5];
  assign m2s0_data_o[4] = m2_data_i[4];
  assign m2s0_data_o[3] = m2_data_i[3];
  assign m2s0_data_o[2] = m2_data_i[2];
  assign m2s0_data_o[1] = m2_data_i[1];
  assign m2s0_data_o[0] = m2_data_i[0];
  assign m2s0_addr[31] = m2_addr_i[31];
  assign m2s0_addr[30] = m2_addr_i[30];
  assign m2s0_addr[29] = m2_addr_i[29];
  assign m2s0_addr[28] = m2_addr_i[28];
  assign m2s0_addr[27] = m2_addr_i[27];
  assign m2s0_addr[26] = m2_addr_i[26];
  assign m2s0_addr[25] = m2_addr_i[25];
  assign m2s0_addr[24] = m2_addr_i[24];
  assign m2s0_addr[23] = m2_addr_i[23];
  assign m2s0_addr[22] = m2_addr_i[22];
  assign m2s0_addr[21] = m2_addr_i[21];
  assign m2s0_addr[20] = m2_addr_i[20];
  assign m2s0_addr[19] = m2_addr_i[19];
  assign m2s0_addr[18] = m2_addr_i[18];
  assign m2s0_addr[17] = m2_addr_i[17];
  assign m2s0_addr[16] = m2_addr_i[16];
  assign m2s0_addr[15] = m2_addr_i[15];
  assign m2s0_addr[14] = m2_addr_i[14];
  assign m2s0_addr[13] = m2_addr_i[13];
  assign m2s0_addr[12] = m2_addr_i[12];
  assign m2s0_addr[11] = m2_addr_i[11];
  assign m2s0_addr[10] = m2_addr_i[10];
  assign m2s0_addr[9] = m2_addr_i[9];
  assign m2s0_addr[8] = m2_addr_i[8];
  assign m2s0_addr[7] = m2_addr_i[7];
  assign m2s0_addr[6] = m2_addr_i[6];
  assign m2s0_addr[5] = m2_addr_i[5];
  assign m2s0_addr[4] = m2_addr_i[4];
  assign m2s0_addr[3] = m2_addr_i[3];
  assign m2s0_addr[2] = m2_addr_i[2];
  assign m2s0_addr[1] = m2_addr_i[1];
  assign m2s0_addr[0] = m2_addr_i[0];
  assign m2s0_sel[3] = m2_sel_i[3];
  assign m2s0_sel[2] = m2_sel_i[2];
  assign m2s0_sel[1] = m2_sel_i[1];
  assign m2s0_sel[0] = m2_sel_i[0];
  assign m2s0_we = m2_we_i;
  assign m3s0_data_o[31] = m3_data_i[31];
  assign m3s0_data_o[30] = m3_data_i[30];
  assign m3s0_data_o[29] = m3_data_i[29];
  assign m3s0_data_o[28] = m3_data_i[28];
  assign m3s0_data_o[27] = m3_data_i[27];
  assign m3s0_data_o[26] = m3_data_i[26];
  assign m3s0_data_o[25] = m3_data_i[25];
  assign m3s0_data_o[24] = m3_data_i[24];
  assign m3s0_data_o[23] = m3_data_i[23];
  assign m3s0_data_o[22] = m3_data_i[22];
  assign m3s0_data_o[21] = m3_data_i[21];
  assign m3s0_data_o[20] = m3_data_i[20];
  assign m3s0_data_o[19] = m3_data_i[19];
  assign m3s0_data_o[18] = m3_data_i[18];
  assign m3s0_data_o[17] = m3_data_i[17];
  assign m3s0_data_o[16] = m3_data_i[16];
  assign m3s0_data_o[15] = m3_data_i[15];
  assign m3s0_data_o[14] = m3_data_i[14];
  assign m3s0_data_o[13] = m3_data_i[13];
  assign m3s0_data_o[12] = m3_data_i[12];
  assign m3s0_data_o[11] = m3_data_i[11];
  assign m3s0_data_o[10] = m3_data_i[10];
  assign m3s0_data_o[9] = m3_data_i[9];
  assign m3s0_data_o[8] = m3_data_i[8];
  assign m3s0_data_o[7] = m3_data_i[7];
  assign m3s0_data_o[6] = m3_data_i[6];
  assign m3s0_data_o[5] = m3_data_i[5];
  assign m3s0_data_o[4] = m3_data_i[4];
  assign m3s0_data_o[3] = m3_data_i[3];
  assign m3s0_data_o[2] = m3_data_i[2];
  assign m3s0_data_o[1] = m3_data_i[1];
  assign m3s0_data_o[0] = m3_data_i[0];
  assign m3s0_addr[31] = m3_addr_i[31];
  assign m3s0_addr[30] = m3_addr_i[30];
  assign m3s0_addr[29] = m3_addr_i[29];
  assign m3s0_addr[28] = m3_addr_i[28];
  assign m3s0_addr[27] = m3_addr_i[27];
  assign m3s0_addr[26] = m3_addr_i[26];
  assign m3s0_addr[25] = m3_addr_i[25];
  assign m3s0_addr[24] = m3_addr_i[24];
  assign m3s0_addr[23] = m3_addr_i[23];
  assign m3s0_addr[22] = m3_addr_i[22];
  assign m3s0_addr[21] = m3_addr_i[21];
  assign m3s0_addr[20] = m3_addr_i[20];
  assign m3s0_addr[19] = m3_addr_i[19];
  assign m3s0_addr[18] = m3_addr_i[18];
  assign m3s0_addr[17] = m3_addr_i[17];
  assign m3s0_addr[16] = m3_addr_i[16];
  assign m3s0_addr[15] = m3_addr_i[15];
  assign m3s0_addr[14] = m3_addr_i[14];
  assign m3s0_addr[13] = m3_addr_i[13];
  assign m3s0_addr[12] = m3_addr_i[12];
  assign m3s0_addr[11] = m3_addr_i[11];
  assign m3s0_addr[10] = m3_addr_i[10];
  assign m3s0_addr[9] = m3_addr_i[9];
  assign m3s0_addr[8] = m3_addr_i[8];
  assign m3s0_addr[7] = m3_addr_i[7];
  assign m3s0_addr[6] = m3_addr_i[6];
  assign m3s0_addr[5] = m3_addr_i[5];
  assign m3s0_addr[4] = m3_addr_i[4];
  assign m3s0_addr[3] = m3_addr_i[3];
  assign m3s0_addr[2] = m3_addr_i[2];
  assign m3s0_addr[1] = m3_addr_i[1];
  assign m3s0_addr[0] = m3_addr_i[0];
  assign m3s0_sel[3] = m3_sel_i[3];
  assign m3s0_sel[2] = m3_sel_i[2];
  assign m3s0_sel[1] = m3_sel_i[1];
  assign m3s0_sel[0] = m3_sel_i[0];
  assign m3s0_we = m3_we_i;
  assign m4s0_data_o[31] = m4_data_i[31];
  assign m4s0_data_o[30] = m4_data_i[30];
  assign m4s0_data_o[29] = m4_data_i[29];
  assign m4s0_data_o[28] = m4_data_i[28];
  assign m4s0_data_o[27] = m4_data_i[27];
  assign m4s0_data_o[26] = m4_data_i[26];
  assign m4s0_data_o[25] = m4_data_i[25];
  assign m4s0_data_o[24] = m4_data_i[24];
  assign m4s0_data_o[23] = m4_data_i[23];
  assign m4s0_data_o[22] = m4_data_i[22];
  assign m4s0_data_o[21] = m4_data_i[21];
  assign m4s0_data_o[20] = m4_data_i[20];
  assign m4s0_data_o[19] = m4_data_i[19];
  assign m4s0_data_o[18] = m4_data_i[18];
  assign m4s0_data_o[17] = m4_data_i[17];
  assign m4s0_data_o[16] = m4_data_i[16];
  assign m4s0_data_o[15] = m4_data_i[15];
  assign m4s0_data_o[14] = m4_data_i[14];
  assign m4s0_data_o[13] = m4_data_i[13];
  assign m4s0_data_o[12] = m4_data_i[12];
  assign m4s0_data_o[11] = m4_data_i[11];
  assign m4s0_data_o[10] = m4_data_i[10];
  assign m4s0_data_o[9] = m4_data_i[9];
  assign m4s0_data_o[8] = m4_data_i[8];
  assign m4s0_data_o[7] = m4_data_i[7];
  assign m4s0_data_o[6] = m4_data_i[6];
  assign m4s0_data_o[5] = m4_data_i[5];
  assign m4s0_data_o[4] = m4_data_i[4];
  assign m4s0_data_o[3] = m4_data_i[3];
  assign m4s0_data_o[2] = m4_data_i[2];
  assign m4s0_data_o[1] = m4_data_i[1];
  assign m4s0_data_o[0] = m4_data_i[0];
  assign m4s0_addr[31] = m4_addr_i[31];
  assign m4s0_addr[30] = m4_addr_i[30];
  assign m4s0_addr[29] = m4_addr_i[29];
  assign m4s0_addr[28] = m4_addr_i[28];
  assign m4s0_addr[27] = m4_addr_i[27];
  assign m4s0_addr[26] = m4_addr_i[26];
  assign m4s0_addr[25] = m4_addr_i[25];
  assign m4s0_addr[24] = m4_addr_i[24];
  assign m4s0_addr[23] = m4_addr_i[23];
  assign m4s0_addr[22] = m4_addr_i[22];
  assign m4s0_addr[21] = m4_addr_i[21];
  assign m4s0_addr[20] = m4_addr_i[20];
  assign m4s0_addr[19] = m4_addr_i[19];
  assign m4s0_addr[18] = m4_addr_i[18];
  assign m4s0_addr[17] = m4_addr_i[17];
  assign m4s0_addr[16] = m4_addr_i[16];
  assign m4s0_addr[15] = m4_addr_i[15];
  assign m4s0_addr[14] = m4_addr_i[14];
  assign m4s0_addr[13] = m4_addr_i[13];
  assign m4s0_addr[12] = m4_addr_i[12];
  assign m4s0_addr[11] = m4_addr_i[11];
  assign m4s0_addr[10] = m4_addr_i[10];
  assign m4s0_addr[9] = m4_addr_i[9];
  assign m4s0_addr[8] = m4_addr_i[8];
  assign m4s0_addr[7] = m4_addr_i[7];
  assign m4s0_addr[6] = m4_addr_i[6];
  assign m4s0_addr[5] = m4_addr_i[5];
  assign m4s0_addr[4] = m4_addr_i[4];
  assign m4s0_addr[3] = m4_addr_i[3];
  assign m4s0_addr[2] = m4_addr_i[2];
  assign m4s0_addr[1] = m4_addr_i[1];
  assign m4s0_addr[0] = m4_addr_i[0];
  assign m4s0_sel[3] = m4_sel_i[3];
  assign m4s0_sel[2] = m4_sel_i[2];
  assign m4s0_sel[1] = m4_sel_i[1];
  assign m4s0_sel[0] = m4_sel_i[0];
  assign m4s0_we = m4_we_i;
  assign m5s0_data_o[31] = m5_data_i[31];
  assign m5s0_data_o[30] = m5_data_i[30];
  assign m5s0_data_o[29] = m5_data_i[29];
  assign m5s0_data_o[28] = m5_data_i[28];
  assign m5s0_data_o[27] = m5_data_i[27];
  assign m5s0_data_o[26] = m5_data_i[26];
  assign m5s0_data_o[25] = m5_data_i[25];
  assign m5s0_data_o[24] = m5_data_i[24];
  assign m5s0_data_o[23] = m5_data_i[23];
  assign m5s0_data_o[22] = m5_data_i[22];
  assign m5s0_data_o[21] = m5_data_i[21];
  assign m5s0_data_o[20] = m5_data_i[20];
  assign m5s0_data_o[19] = m5_data_i[19];
  assign m5s0_data_o[18] = m5_data_i[18];
  assign m5s0_data_o[17] = m5_data_i[17];
  assign m5s0_data_o[16] = m5_data_i[16];
  assign m5s0_data_o[15] = m5_data_i[15];
  assign m5s0_data_o[14] = m5_data_i[14];
  assign m5s0_data_o[13] = m5_data_i[13];
  assign m5s0_data_o[12] = m5_data_i[12];
  assign m5s0_data_o[11] = m5_data_i[11];
  assign m5s0_data_o[10] = m5_data_i[10];
  assign m5s0_data_o[9] = m5_data_i[9];
  assign m5s0_data_o[8] = m5_data_i[8];
  assign m5s0_data_o[7] = m5_data_i[7];
  assign m5s0_data_o[6] = m5_data_i[6];
  assign m5s0_data_o[5] = m5_data_i[5];
  assign m5s0_data_o[4] = m5_data_i[4];
  assign m5s0_data_o[3] = m5_data_i[3];
  assign m5s0_data_o[2] = m5_data_i[2];
  assign m5s0_data_o[1] = m5_data_i[1];
  assign m5s0_data_o[0] = m5_data_i[0];
  assign m5s0_addr[31] = m5_addr_i[31];
  assign m5s0_addr[30] = m5_addr_i[30];
  assign m5s0_addr[29] = m5_addr_i[29];
  assign m5s0_addr[28] = m5_addr_i[28];
  assign m5s0_addr[27] = m5_addr_i[27];
  assign m5s0_addr[26] = m5_addr_i[26];
  assign m5s0_addr[25] = m5_addr_i[25];
  assign m5s0_addr[24] = m5_addr_i[24];
  assign m5s0_addr[23] = m5_addr_i[23];
  assign m5s0_addr[22] = m5_addr_i[22];
  assign m5s0_addr[21] = m5_addr_i[21];
  assign m5s0_addr[20] = m5_addr_i[20];
  assign m5s0_addr[19] = m5_addr_i[19];
  assign m5s0_addr[18] = m5_addr_i[18];
  assign m5s0_addr[17] = m5_addr_i[17];
  assign m5s0_addr[16] = m5_addr_i[16];
  assign m5s0_addr[15] = m5_addr_i[15];
  assign m5s0_addr[14] = m5_addr_i[14];
  assign m5s0_addr[13] = m5_addr_i[13];
  assign m5s0_addr[12] = m5_addr_i[12];
  assign m5s0_addr[11] = m5_addr_i[11];
  assign m5s0_addr[10] = m5_addr_i[10];
  assign m5s0_addr[9] = m5_addr_i[9];
  assign m5s0_addr[8] = m5_addr_i[8];
  assign m5s0_addr[7] = m5_addr_i[7];
  assign m5s0_addr[6] = m5_addr_i[6];
  assign m5s0_addr[5] = m5_addr_i[5];
  assign m5s0_addr[4] = m5_addr_i[4];
  assign m5s0_addr[3] = m5_addr_i[3];
  assign m5s0_addr[2] = m5_addr_i[2];
  assign m5s0_addr[1] = m5_addr_i[1];
  assign m5s0_addr[0] = m5_addr_i[0];
  assign m5s0_sel[3] = m5_sel_i[3];
  assign m5s0_sel[2] = m5_sel_i[2];
  assign m5s0_sel[1] = m5_sel_i[1];
  assign m5s0_sel[0] = m5_sel_i[0];
  assign m5s0_we = m5_we_i;
  assign m6s0_data_o[31] = m6_data_i[31];
  assign m6s0_data_o[30] = m6_data_i[30];
  assign m6s0_data_o[29] = m6_data_i[29];
  assign m6s0_data_o[28] = m6_data_i[28];
  assign m6s0_data_o[27] = m6_data_i[27];
  assign m6s0_data_o[26] = m6_data_i[26];
  assign m6s0_data_o[25] = m6_data_i[25];
  assign m6s0_data_o[24] = m6_data_i[24];
  assign m6s0_data_o[23] = m6_data_i[23];
  assign m6s0_data_o[22] = m6_data_i[22];
  assign m6s0_data_o[21] = m6_data_i[21];
  assign m6s0_data_o[20] = m6_data_i[20];
  assign m6s0_data_o[19] = m6_data_i[19];
  assign m6s0_data_o[18] = m6_data_i[18];
  assign m6s0_data_o[17] = m6_data_i[17];
  assign m6s0_data_o[16] = m6_data_i[16];
  assign m6s0_data_o[15] = m6_data_i[15];
  assign m6s0_data_o[14] = m6_data_i[14];
  assign m6s0_data_o[13] = m6_data_i[13];
  assign m6s0_data_o[12] = m6_data_i[12];
  assign m6s0_data_o[11] = m6_data_i[11];
  assign m6s0_data_o[10] = m6_data_i[10];
  assign m6s0_data_o[9] = m6_data_i[9];
  assign m6s0_data_o[8] = m6_data_i[8];
  assign m6s0_data_o[7] = m6_data_i[7];
  assign m6s0_data_o[6] = m6_data_i[6];
  assign m6s0_data_o[5] = m6_data_i[5];
  assign m6s0_data_o[4] = m6_data_i[4];
  assign m6s0_data_o[3] = m6_data_i[3];
  assign m6s0_data_o[2] = m6_data_i[2];
  assign m6s0_data_o[1] = m6_data_i[1];
  assign m6s0_data_o[0] = m6_data_i[0];
  assign m6s0_addr[31] = m6_addr_i[31];
  assign m6s0_addr[30] = m6_addr_i[30];
  assign m6s0_addr[29] = m6_addr_i[29];
  assign m6s0_addr[28] = m6_addr_i[28];
  assign m6s0_addr[27] = m6_addr_i[27];
  assign m6s0_addr[26] = m6_addr_i[26];
  assign m6s0_addr[25] = m6_addr_i[25];
  assign m6s0_addr[24] = m6_addr_i[24];
  assign m6s0_addr[23] = m6_addr_i[23];
  assign m6s0_addr[22] = m6_addr_i[22];
  assign m6s0_addr[21] = m6_addr_i[21];
  assign m6s0_addr[20] = m6_addr_i[20];
  assign m6s0_addr[19] = m6_addr_i[19];
  assign m6s0_addr[18] = m6_addr_i[18];
  assign m6s0_addr[17] = m6_addr_i[17];
  assign m6s0_addr[16] = m6_addr_i[16];
  assign m6s0_addr[15] = m6_addr_i[15];
  assign m6s0_addr[14] = m6_addr_i[14];
  assign m6s0_addr[13] = m6_addr_i[13];
  assign m6s0_addr[12] = m6_addr_i[12];
  assign m6s0_addr[11] = m6_addr_i[11];
  assign m6s0_addr[10] = m6_addr_i[10];
  assign m6s0_addr[9] = m6_addr_i[9];
  assign m6s0_addr[8] = m6_addr_i[8];
  assign m6s0_addr[7] = m6_addr_i[7];
  assign m6s0_addr[6] = m6_addr_i[6];
  assign m6s0_addr[5] = m6_addr_i[5];
  assign m6s0_addr[4] = m6_addr_i[4];
  assign m6s0_addr[3] = m6_addr_i[3];
  assign m6s0_addr[2] = m6_addr_i[2];
  assign m6s0_addr[1] = m6_addr_i[1];
  assign m6s0_addr[0] = m6_addr_i[0];
  assign m6s0_sel[3] = m6_sel_i[3];
  assign m6s0_sel[2] = m6_sel_i[2];
  assign m6s0_sel[1] = m6_sel_i[1];
  assign m6s0_sel[0] = m6_sel_i[0];
  assign m6s0_we = m6_we_i;
  assign m7s0_data_o[31] = m7_data_i[31];
  assign m7s0_data_o[30] = m7_data_i[30];
  assign m7s0_data_o[29] = m7_data_i[29];
  assign m7s0_data_o[28] = m7_data_i[28];
  assign m7s0_data_o[27] = m7_data_i[27];
  assign m7s0_data_o[26] = m7_data_i[26];
  assign m7s0_data_o[25] = m7_data_i[25];
  assign m7s0_data_o[24] = m7_data_i[24];
  assign m7s0_data_o[23] = m7_data_i[23];
  assign m7s0_data_o[22] = m7_data_i[22];
  assign m7s0_data_o[21] = m7_data_i[21];
  assign m7s0_data_o[20] = m7_data_i[20];
  assign m7s0_data_o[19] = m7_data_i[19];
  assign m7s0_data_o[18] = m7_data_i[18];
  assign m7s0_data_o[17] = m7_data_i[17];
  assign m7s0_data_o[16] = m7_data_i[16];
  assign m7s0_data_o[15] = m7_data_i[15];
  assign m7s0_data_o[14] = m7_data_i[14];
  assign m7s0_data_o[13] = m7_data_i[13];
  assign m7s0_data_o[12] = m7_data_i[12];
  assign m7s0_data_o[11] = m7_data_i[11];
  assign m7s0_data_o[10] = m7_data_i[10];
  assign m7s0_data_o[9] = m7_data_i[9];
  assign m7s0_data_o[8] = m7_data_i[8];
  assign m7s0_data_o[7] = m7_data_i[7];
  assign m7s0_data_o[6] = m7_data_i[6];
  assign m7s0_data_o[5] = m7_data_i[5];
  assign m7s0_data_o[4] = m7_data_i[4];
  assign m7s0_data_o[3] = m7_data_i[3];
  assign m7s0_data_o[2] = m7_data_i[2];
  assign m7s0_data_o[1] = m7_data_i[1];
  assign m7s0_data_o[0] = m7_data_i[0];
  assign m7s0_addr[31] = m7_addr_i[31];
  assign m7s0_addr[30] = m7_addr_i[30];
  assign m7s0_addr[29] = m7_addr_i[29];
  assign m7s0_addr[28] = m7_addr_i[28];
  assign m7s0_addr[27] = m7_addr_i[27];
  assign m7s0_addr[26] = m7_addr_i[26];
  assign m7s0_addr[25] = m7_addr_i[25];
  assign m7s0_addr[24] = m7_addr_i[24];
  assign m7s0_addr[23] = m7_addr_i[23];
  assign m7s0_addr[22] = m7_addr_i[22];
  assign m7s0_addr[21] = m7_addr_i[21];
  assign m7s0_addr[20] = m7_addr_i[20];
  assign m7s0_addr[19] = m7_addr_i[19];
  assign m7s0_addr[18] = m7_addr_i[18];
  assign m7s0_addr[17] = m7_addr_i[17];
  assign m7s0_addr[16] = m7_addr_i[16];
  assign m7s0_addr[15] = m7_addr_i[15];
  assign m7s0_addr[14] = m7_addr_i[14];
  assign m7s0_addr[13] = m7_addr_i[13];
  assign m7s0_addr[12] = m7_addr_i[12];
  assign m7s0_addr[11] = m7_addr_i[11];
  assign m7s0_addr[10] = m7_addr_i[10];
  assign m7s0_addr[9] = m7_addr_i[9];
  assign m7s0_addr[8] = m7_addr_i[8];
  assign m7s0_addr[7] = m7_addr_i[7];
  assign m7s0_addr[6] = m7_addr_i[6];
  assign m7s0_addr[5] = m7_addr_i[5];
  assign m7s0_addr[4] = m7_addr_i[4];
  assign m7s0_addr[3] = m7_addr_i[3];
  assign m7s0_addr[2] = m7_addr_i[2];
  assign m7s0_addr[1] = m7_addr_i[1];
  assign m7s0_addr[0] = m7_addr_i[0];
  assign m7s0_sel[3] = m7_sel_i[3];
  assign m7s0_sel[2] = m7_sel_i[2];
  assign m7s0_sel[1] = m7_sel_i[1];
  assign m7s0_sel[0] = m7_sel_i[0];
  assign m7s0_we = m7_we_i;

  DFFARX1 \m0/s15_cyc_o_reg  ( .D(n18177), .CLK(clock), .RSTB(n34690), .Q(
        m0s15_cyc) );
  DFFARX1 \m0/s14_cyc_o_reg  ( .D(n18176), .CLK(clock), .RSTB(n34690), .Q(
        m0s14_cyc) );
  DFFARX1 \m0/s13_cyc_o_reg  ( .D(n18175), .CLK(clock), .RSTB(n34678), .Q(
        m0s13_cyc) );
  DFFARX1 \m0/s12_cyc_o_reg  ( .D(n18174), .CLK(clock), .RSTB(n34691), .Q(
        m0s12_cyc) );
  DFFARX1 \m0/s11_cyc_o_reg  ( .D(n18173), .CLK(clock), .RSTB(n34687), .Q(
        m0s11_cyc) );
  DFFARX1 \m0/s10_cyc_o_reg  ( .D(n18172), .CLK(clock), .RSTB(n34686), .Q(
        m0s10_cyc) );
  DFFARX1 \m0/s9_cyc_o_reg  ( .D(n18171), .CLK(clock), .RSTB(n34680), .Q(
        m0s9_cyc) );
  DFFARX1 \m0/s8_cyc_o_reg  ( .D(n18170), .CLK(clock), .RSTB(n34682), .Q(
        m0s8_cyc) );
  DFFARX1 \m0/s7_cyc_o_reg  ( .D(n18169), .CLK(clock), .RSTB(n34694), .Q(
        m0s7_cyc) );
  DFFARX1 \m0/s6_cyc_o_reg  ( .D(n18168), .CLK(clock), .RSTB(n34683), .Q(
        m0s6_cyc) );
  DFFARX1 \m0/s5_cyc_o_reg  ( .D(n18167), .CLK(clock), .RSTB(n34697), .Q(
        m0s5_cyc) );
  DFFARX1 \m0/s4_cyc_o_reg  ( .D(n18166), .CLK(clock), .RSTB(n34684), .Q(
        m0s4_cyc) );
  DFFARX1 \m0/s3_cyc_o_reg  ( .D(n18165), .CLK(clock), .RSTB(n34683), .Q(
        m0s3_cyc) );
  DFFARX1 \m0/s2_cyc_o_reg  ( .D(n18164), .CLK(clock), .RSTB(n34695), .Q(
        m0s2_cyc) );
  DFFARX1 \m0/s1_cyc_o_reg  ( .D(n18163), .CLK(clock), .RSTB(n34690), .Q(
        m0s1_cyc) );
  DFFARX1 \m0/s0_cyc_o_reg  ( .D(n18162), .CLK(clock), .RSTB(n34685), .Q(
        m0s0_cyc) );
  DFFARX1 \m1/s15_cyc_o_reg  ( .D(n18161), .CLK(clock), .RSTB(n34687), .Q(
        m1s15_cyc) );
  DFFARX1 \m1/s14_cyc_o_reg  ( .D(n18160), .CLK(clock), .RSTB(n34696), .Q(
        m1s14_cyc) );
  DFFARX1 \m1/s13_cyc_o_reg  ( .D(n18159), .CLK(clock), .RSTB(n34678), .Q(
        m1s13_cyc) );
  DFFARX1 \m1/s12_cyc_o_reg  ( .D(n18158), .CLK(clock), .RSTB(n34678), .Q(
        m1s12_cyc) );
  DFFARX1 \m1/s11_cyc_o_reg  ( .D(n18157), .CLK(clock), .RSTB(n34677), .Q(
        m1s11_cyc) );
  DFFARX1 \m1/s10_cyc_o_reg  ( .D(n18156), .CLK(clock), .RSTB(n34687), .Q(
        m1s10_cyc) );
  DFFARX1 \m1/s9_cyc_o_reg  ( .D(n18155), .CLK(clock), .RSTB(n34691), .Q(
        m1s9_cyc) );
  DFFARX1 \m1/s8_cyc_o_reg  ( .D(n18154), .CLK(clock), .RSTB(n34688), .Q(
        m1s8_cyc) );
  DFFARX1 \m1/s7_cyc_o_reg  ( .D(n18153), .CLK(clock), .RSTB(n34680), .Q(
        m1s7_cyc) );
  DFFARX1 \m1/s6_cyc_o_reg  ( .D(n18152), .CLK(clock), .RSTB(n34682), .Q(
        m1s6_cyc) );
  DFFARX1 \m1/s5_cyc_o_reg  ( .D(n18151), .CLK(clock), .RSTB(n34686), .Q(
        m1s5_cyc) );
  DFFARX1 \m1/s4_cyc_o_reg  ( .D(n18150), .CLK(clock), .RSTB(n34691), .Q(
        m1s4_cyc) );
  DFFARX1 \m1/s3_cyc_o_reg  ( .D(n18149), .CLK(clock), .RSTB(n34684), .Q(
        m1s3_cyc) );
  DFFARX1 \m1/s2_cyc_o_reg  ( .D(n18148), .CLK(clock), .RSTB(n34679), .Q(
        m1s2_cyc) );
  DFFARX1 \m1/s1_cyc_o_reg  ( .D(n18147), .CLK(clock), .RSTB(n34686), .Q(
        m1s1_cyc) );
  DFFARX1 \m1/s0_cyc_o_reg  ( .D(n18146), .CLK(clock), .RSTB(n34692), .Q(
        m1s0_cyc) );
  DFFARX1 \m2/s15_cyc_o_reg  ( .D(n18145), .CLK(clock), .RSTB(n34689), .Q(
        m2s15_cyc) );
  DFFARX1 \m2/s14_cyc_o_reg  ( .D(n18144), .CLK(clock), .RSTB(n34685), .Q(
        m2s14_cyc) );
  DFFARX1 \m2/s13_cyc_o_reg  ( .D(n18143), .CLK(clock), .RSTB(n34695), .Q(
        m2s13_cyc) );
  DFFARX1 \m2/s12_cyc_o_reg  ( .D(n18142), .CLK(clock), .RSTB(n34678), .Q(
        m2s12_cyc) );
  DFFARX1 \m2/s11_cyc_o_reg  ( .D(n18141), .CLK(clock), .RSTB(n34688), .Q(
        m2s11_cyc) );
  DFFARX1 \m2/s10_cyc_o_reg  ( .D(n18140), .CLK(clock), .RSTB(n34677), .Q(
        m2s10_cyc) );
  DFFARX1 \m2/s9_cyc_o_reg  ( .D(n18139), .CLK(clock), .RSTB(n34681), .Q(
        m2s9_cyc) );
  DFFARX1 \m2/s8_cyc_o_reg  ( .D(n18138), .CLK(clock), .RSTB(n34686), .Q(
        m2s8_cyc) );
  DFFARX1 \m2/s7_cyc_o_reg  ( .D(n18137), .CLK(clock), .RSTB(n34692), .Q(
        m2s7_cyc) );
  DFFARX1 \m2/s6_cyc_o_reg  ( .D(n18136), .CLK(clock), .RSTB(n34694), .Q(
        m2s6_cyc) );
  DFFARX1 \m2/s5_cyc_o_reg  ( .D(n18135), .CLK(clock), .RSTB(n34679), .Q(
        m2s5_cyc) );
  DFFARX1 \m2/s4_cyc_o_reg  ( .D(n18134), .CLK(clock), .RSTB(n34695), .Q(
        m2s4_cyc) );
  DFFARX1 \m2/s3_cyc_o_reg  ( .D(n18133), .CLK(clock), .RSTB(n34696), .Q(
        m2s3_cyc) );
  DFFARX1 \m2/s2_cyc_o_reg  ( .D(n18132), .CLK(clock), .RSTB(n34678), .Q(
        m2s2_cyc) );
  DFFARX1 \m2/s1_cyc_o_reg  ( .D(n18131), .CLK(clock), .RSTB(n34697), .Q(
        m2s1_cyc) );
  DFFARX1 \m2/s0_cyc_o_reg  ( .D(n18130), .CLK(clock), .RSTB(n34677), .Q(
        m2s0_cyc) );
  DFFARX1 \m3/s15_cyc_o_reg  ( .D(n18129), .CLK(clock), .RSTB(n34681), .Q(
        m3s15_cyc) );
  DFFARX1 \m3/s14_cyc_o_reg  ( .D(n18128), .CLK(clock), .RSTB(n34696), .Q(
        m3s14_cyc) );
  DFFARX1 \m3/s13_cyc_o_reg  ( .D(n18127), .CLK(clock), .RSTB(n34678), .Q(
        m3s13_cyc) );
  DFFARX1 \m3/s12_cyc_o_reg  ( .D(n18126), .CLK(clock), .RSTB(n34688), .Q(
        m3s12_cyc) );
  DFFARX1 \m3/s11_cyc_o_reg  ( .D(n18125), .CLK(clock), .RSTB(n34694), .Q(
        m3s11_cyc) );
  DFFARX1 \m3/s10_cyc_o_reg  ( .D(n18124), .CLK(clock), .RSTB(n34689), .Q(
        m3s10_cyc) );
  DFFARX1 \m3/s9_cyc_o_reg  ( .D(n18123), .CLK(clock), .RSTB(n34690), .Q(
        m3s9_cyc) );
  DFFARX1 \m3/s8_cyc_o_reg  ( .D(n18122), .CLK(clock), .RSTB(n34684), .Q(
        m3s8_cyc) );
  DFFARX1 \m3/s7_cyc_o_reg  ( .D(n18121), .CLK(clock), .RSTB(n34678), .Q(
        m3s7_cyc) );
  DFFARX1 \m3/s6_cyc_o_reg  ( .D(n18120), .CLK(clock), .RSTB(n34691), .Q(
        m3s6_cyc) );
  DFFARX1 \m3/s5_cyc_o_reg  ( .D(n18119), .CLK(clock), .RSTB(n34690), .Q(
        m3s5_cyc) );
  DFFARX1 \m3/s4_cyc_o_reg  ( .D(n18118), .CLK(clock), .RSTB(n34680), .Q(
        m3s4_cyc) );
  DFFARX1 \m3/s3_cyc_o_reg  ( .D(n18117), .CLK(clock), .RSTB(n34682), .Q(
        m3s3_cyc) );
  DFFARX1 \m3/s2_cyc_o_reg  ( .D(n18116), .CLK(clock), .RSTB(n34691), .Q(
        m3s2_cyc) );
  DFFARX1 \m3/s1_cyc_o_reg  ( .D(n18115), .CLK(clock), .RSTB(n34683), .Q(
        m3s1_cyc) );
  DFFARX1 \m3/s0_cyc_o_reg  ( .D(n18114), .CLK(clock), .RSTB(n34686), .Q(
        m3s0_cyc) );
  DFFARX1 \m4/s15_cyc_o_reg  ( .D(n18113), .CLK(clock), .RSTB(n34687), .Q(
        m4s15_cyc) );
  DFFARX1 \m4/s14_cyc_o_reg  ( .D(n18112), .CLK(clock), .RSTB(n34688), .Q(
        m4s14_cyc) );
  DFFARX1 \m4/s13_cyc_o_reg  ( .D(n18111), .CLK(clock), .RSTB(n34685), .Q(
        m4s13_cyc) );
  DFFARX1 \m4/s12_cyc_o_reg  ( .D(n18110), .CLK(clock), .RSTB(n34679), .Q(
        m4s12_cyc) );
  DFFARX1 \m4/s11_cyc_o_reg  ( .D(n18109), .CLK(clock), .RSTB(n34678), .Q(
        m4s11_cyc) );
  DFFARX1 \m4/s10_cyc_o_reg  ( .D(n18108), .CLK(clock), .RSTB(n34685), .Q(
        m4s10_cyc) );
  DFFARX1 \m4/s9_cyc_o_reg  ( .D(n18107), .CLK(clock), .RSTB(n34677), .Q(
        m4s9_cyc) );
  DFFARX1 \m4/s8_cyc_o_reg  ( .D(n18106), .CLK(clock), .RSTB(n34678), .Q(
        m4s8_cyc) );
  DFFARX1 \m4/s7_cyc_o_reg  ( .D(n18105), .CLK(clock), .RSTB(n34683), .Q(
        m4s7_cyc) );
  DFFARX1 \m4/s6_cyc_o_reg  ( .D(n18104), .CLK(clock), .RSTB(n34690), .Q(
        m4s6_cyc) );
  DFFARX1 \m4/s5_cyc_o_reg  ( .D(n18103), .CLK(clock), .RSTB(n34692), .Q(
        m4s5_cyc) );
  DFFARX1 \m4/s4_cyc_o_reg  ( .D(n18102), .CLK(clock), .RSTB(n34696), .Q(
        m4s4_cyc) );
  DFFARX1 \m4/s3_cyc_o_reg  ( .D(n18101), .CLK(clock), .RSTB(n34678), .Q(
        m4s3_cyc) );
  DFFARX1 \m4/s2_cyc_o_reg  ( .D(n18100), .CLK(clock), .RSTB(n34697), .Q(
        m4s2_cyc) );
  DFFARX1 \m4/s1_cyc_o_reg  ( .D(n18099), .CLK(clock), .RSTB(n34678), .Q(
        m4s1_cyc) );
  DFFARX1 \m4/s0_cyc_o_reg  ( .D(n18098), .CLK(clock), .RSTB(n34681), .Q(
        m4s0_cyc) );
  DFFARX1 \m5/s15_cyc_o_reg  ( .D(n18097), .CLK(clock), .RSTB(n34693), .Q(
        m5s15_cyc) );
  DFFARX1 \m5/s14_cyc_o_reg  ( .D(n18096), .CLK(clock), .RSTB(n34685), .Q(
        m5s14_cyc) );
  DFFARX1 \m5/s13_cyc_o_reg  ( .D(n18095), .CLK(clock), .RSTB(n34687), .Q(
        m5s13_cyc) );
  DFFARX1 \m5/s12_cyc_o_reg  ( .D(n18094), .CLK(clock), .RSTB(n34680), .Q(
        m5s12_cyc) );
  DFFARX1 \m5/s11_cyc_o_reg  ( .D(n18093), .CLK(clock), .RSTB(n34688), .Q(
        m5s11_cyc) );
  DFFARX1 \m5/s10_cyc_o_reg  ( .D(n18092), .CLK(clock), .RSTB(n34686), .Q(
        m5s10_cyc) );
  DFFARX1 \m5/s9_cyc_o_reg  ( .D(n18091), .CLK(clock), .RSTB(n34689), .Q(
        m5s9_cyc) );
  DFFARX1 \m5/s8_cyc_o_reg  ( .D(n18090), .CLK(clock), .RSTB(n34691), .Q(
        m5s8_cyc) );
  DFFARX1 \m5/s7_cyc_o_reg  ( .D(n18089), .CLK(clock), .RSTB(n34680), .Q(
        m5s7_cyc) );
  DFFARX1 \m5/s6_cyc_o_reg  ( .D(n18088), .CLK(clock), .RSTB(n34682), .Q(
        m5s6_cyc) );
  DFFARX1 \m5/s5_cyc_o_reg  ( .D(n18087), .CLK(clock), .RSTB(n34692), .Q(
        m5s5_cyc) );
  DFFARX1 \m5/s4_cyc_o_reg  ( .D(n18086), .CLK(clock), .RSTB(n34683), .Q(
        m5s4_cyc) );
  DFFARX1 \m5/s3_cyc_o_reg  ( .D(n18085), .CLK(clock), .RSTB(n34695), .Q(
        m5s3_cyc) );
  DFFARX1 \m5/s2_cyc_o_reg  ( .D(n18084), .CLK(clock), .RSTB(n34684), .Q(
        m5s2_cyc) );
  DFFARX1 \m5/s1_cyc_o_reg  ( .D(n18083), .CLK(clock), .RSTB(n34686), .Q(
        m5s1_cyc) );
  DFFARX1 \m5/s0_cyc_o_reg  ( .D(n18082), .CLK(clock), .RSTB(n34681), .Q(
        m5s0_cyc) );
  DFFARX1 \m6/s15_cyc_o_reg  ( .D(n18081), .CLK(clock), .RSTB(n34685), .Q(
        m6s15_cyc) );
  DFFARX1 \m6/s14_cyc_o_reg  ( .D(n18080), .CLK(clock), .RSTB(n34694), .Q(
        m6s14_cyc) );
  DFFARX1 \m6/s13_cyc_o_reg  ( .D(n18079), .CLK(clock), .RSTB(n34687), .Q(
        m6s13_cyc) );
  DFFARX1 \m6/s12_cyc_o_reg  ( .D(n18078), .CLK(clock), .RSTB(n34692), .Q(
        m6s12_cyc) );
  DFFARX1 \m6/s11_cyc_o_reg  ( .D(n18077), .CLK(clock), .RSTB(n34692), .Q(
        m6s11_cyc) );
  DFFARX1 \m6/s10_cyc_o_reg  ( .D(n18076), .CLK(clock), .RSTB(n34694), .Q(
        m6s10_cyc) );
  DFFARX1 \m6/s9_cyc_o_reg  ( .D(n18075), .CLK(clock), .RSTB(n34679), .Q(
        m6s9_cyc) );
  DFFARX1 \m6/s8_cyc_o_reg  ( .D(n18074), .CLK(clock), .RSTB(n34695), .Q(
        m6s8_cyc) );
  DFFARX1 \m6/s7_cyc_o_reg  ( .D(n18073), .CLK(clock), .RSTB(n34696), .Q(
        m6s7_cyc) );
  DFFARX1 \m6/s6_cyc_o_reg  ( .D(n18072), .CLK(clock), .RSTB(n34685), .Q(
        m6s6_cyc) );
  DFFARX1 \m6/s5_cyc_o_reg  ( .D(n18071), .CLK(clock), .RSTB(n34697), .Q(
        m6s5_cyc) );
  DFFARX1 \m6/s4_cyc_o_reg  ( .D(n18070), .CLK(clock), .RSTB(n34677), .Q(
        m6s4_cyc) );
  DFFARX1 \m6/s3_cyc_o_reg  ( .D(n18069), .CLK(clock), .RSTB(n34681), .Q(
        m6s3_cyc) );
  DFFARX1 \m6/s2_cyc_o_reg  ( .D(n18068), .CLK(clock), .RSTB(n34693), .Q(
        m6s2_cyc) );
  DFFARX1 \m6/s1_cyc_o_reg  ( .D(n18067), .CLK(clock), .RSTB(n34689), .Q(
        m6s1_cyc) );
  DFFARX1 \m6/s0_cyc_o_reg  ( .D(n18066), .CLK(clock), .RSTB(n34690), .Q(
        m6s0_cyc) );
  DFFARX1 \m7/s15_cyc_o_reg  ( .D(n18065), .CLK(clock), .RSTB(n34682), .Q(
        m7s15_cyc) );
  DFFARX1 \m7/s14_cyc_o_reg  ( .D(n18064), .CLK(clock), .RSTB(n34685), .Q(
        m7s14_cyc) );
  DFFARX1 \m7/s13_cyc_o_reg  ( .D(n18063), .CLK(clock), .RSTB(n34691), .Q(
        m7s13_cyc) );
  DFFARX1 \m7/s12_cyc_o_reg  ( .D(n18062), .CLK(clock), .RSTB(n34680), .Q(
        m7s12_cyc) );
  DFFARX1 \m7/s11_cyc_o_reg  ( .D(n18061), .CLK(clock), .RSTB(n34682), .Q(
        m7s11_cyc) );
  DFFARX1 \m7/s10_cyc_o_reg  ( .D(n18060), .CLK(clock), .RSTB(n34683), .Q(
        m7s10_cyc) );
  DFFARX1 \m7/s9_cyc_o_reg  ( .D(n18059), .CLK(clock), .RSTB(n34683), .Q(
        m7s9_cyc) );
  DFFARX1 \m7/s8_cyc_o_reg  ( .D(n18058), .CLK(clock), .RSTB(n34679), .Q(
        m7s8_cyc) );
  DFFARX1 \m7/s7_cyc_o_reg  ( .D(n18057), .CLK(clock), .RSTB(n34684), .Q(
        m7s7_cyc) );
  DFFARX1 \m7/s6_cyc_o_reg  ( .D(n18056), .CLK(clock), .RSTB(n34686), .Q(
        m7s6_cyc) );
  DFFARX1 \m7/s5_cyc_o_reg  ( .D(n18055), .CLK(clock), .RSTB(n34677), .Q(
        m7s5_cyc) );
  DFFARX1 \m7/s4_cyc_o_reg  ( .D(n18054), .CLK(clock), .RSTB(n34677), .Q(
        m7s4_cyc) );
  DFFARX1 \m7/s3_cyc_o_reg  ( .D(n18053), .CLK(clock), .RSTB(n34692), .Q(
        m7s3_cyc) );
  DFFARX1 \m7/s2_cyc_o_reg  ( .D(n18052), .CLK(clock), .RSTB(n34685), .Q(
        m7s2_cyc) );
  DFFARX1 \m7/s1_cyc_o_reg  ( .D(n18051), .CLK(clock), .RSTB(n34693), .Q(
        m7s1_cyc) );
  DFFARX1 \m7/s0_cyc_o_reg  ( .D(n18050), .CLK(clock), .RSTB(n34688), .Q(
        m7s0_cyc) );
  DFFARX1 \s0/msel/arb1/state_reg[0]  ( .D(n18028), .CLK(clock), .RSTB(n34694), 
        .Q(\s0/msel/gnt_p1 [0]), .QN(n34250) );
  DFFARX1 \s0/msel/arb1/state_reg[1]  ( .D(n18029), .CLK(clock), .RSTB(n34679), 
        .Q(\s0/msel/gnt_p1 [1]), .QN(n34669) );
  DFFARX1 \s0/msel/arb1/state_reg[2]  ( .D(n18030), .CLK(clock), .RSTB(n34695), 
        .Q(\s0/msel/gnt_p1 [2]), .QN(n34432) );
  DFFARX1 \s0/msel/arb0/state_reg[0]  ( .D(n18025), .CLK(clock), .RSTB(n34696), 
        .Q(\s0/msel/gnt_p0 [0]), .QN(n34240) );
  DFFARX1 \s0/msel/arb0/state_reg[1]  ( .D(n18026), .CLK(clock), .RSTB(n34684), 
        .Q(\s0/msel/gnt_p0 [1]), .QN(n34453) );
  DFFARX1 \s0/msel/arb0/state_reg[2]  ( .D(n18027), .CLK(clock), .RSTB(n34697), 
        .Q(\s0/msel/gnt_p0 [2]), .QN(n34440) );
  DFFARX1 \s0/msel/arb3/state_reg[0]  ( .D(n18031), .CLK(clock), .RSTB(n34685), 
        .Q(\s0/msel/gnt_p3 [0]), .QN(n34259) );
  DFFARX1 \s0/msel/arb3/state_reg[1]  ( .D(n18032), .CLK(clock), .RSTB(n34677), 
        .Q(\s0/msel/gnt_p3 [1]), .QN(n34423) );
  DFFARX1 \s0/msel/arb3/state_reg[2]  ( .D(n18033), .CLK(clock), .RSTB(n34677), 
        .Q(\s0/msel/gnt_p3 [2]), .QN(n34549) );
  DFFARX1 \s0/msel/arb2/state_reg[0]  ( .D(n18022), .CLK(clock), .RSTB(n34677), 
        .Q(\s0/msel/gnt_p2 [0]), .QN(n34290) );
  DFFARX1 \s0/msel/arb2/state_reg[1]  ( .D(n18023), .CLK(clock), .RSTB(n34677), 
        .Q(\s0/msel/gnt_p2 [1]), .QN(n34286) );
  DFFARX1 \s0/msel/arb2/state_reg[2]  ( .D(n18024), .CLK(clock), .RSTB(n34677), 
        .Q(\s0/msel/gnt_p2 [2]), .QN(n34473) );
  DFFARX1 \s2/msel/arb1/state_reg[0]  ( .D(n17972), .CLK(clock), .RSTB(n34677), 
        .Q(\s2/msel/gnt_p1 [0]), .QN(n34241) );
  DFFARX1 \s2/msel/arb1/state_reg[1]  ( .D(n17973), .CLK(clock), .RSTB(n34677), 
        .Q(\s2/msel/gnt_p1 [1]), .QN(n34383) );
  DFFARX1 \s2/msel/arb1/state_reg[2]  ( .D(n17974), .CLK(clock), .RSTB(n34677), 
        .Q(\s2/msel/gnt_p1 [2]), .QN(n34438) );
  DFFARX1 \s2/msel/arb0/state_reg[0]  ( .D(n17969), .CLK(clock), .RSTB(n34677), 
        .Q(\s2/msel/gnt_p0 [0]), .QN(n34554) );
  DFFARX1 \s2/msel/arb0/state_reg[1]  ( .D(n17970), .CLK(clock), .RSTB(n34677), 
        .Q(\s2/msel/gnt_p0 [1]), .QN(n34670) );
  DFFARX1 \s2/msel/arb0/state_reg[2]  ( .D(n17971), .CLK(clock), .RSTB(n34677), 
        .Q(\s2/msel/gnt_p0 [2]), .QN(n34291) );
  DFFARX1 \s2/msel/arb3/state_reg[0]  ( .D(n17975), .CLK(clock), .RSTB(n34677), 
        .Q(\s2/msel/gnt_p3 [0]), .QN(n34277) );
  DFFARX1 \s2/msel/arb3/state_reg[1]  ( .D(n17976), .CLK(clock), .RSTB(n34692), 
        .Q(\s2/msel/gnt_p3 [1]), .QN(n34395) );
  DFFARX1 \s2/msel/arb3/state_reg[2]  ( .D(n17977), .CLK(clock), .RSTB(n34689), 
        .Q(\s2/msel/gnt_p3 [2]), .QN(n34548) );
  DFFARX1 \s2/msel/arb2/state_reg[0]  ( .D(n17966), .CLK(clock), .RSTB(n34690), 
        .Q(\s2/msel/gnt_p2 [0]), .QN(n34609) );
  DFFARX1 \s2/msel/arb2/state_reg[1]  ( .D(n17967), .CLK(clock), .RSTB(n34687), 
        .Q(\s2/msel/gnt_p2 [1]), .QN(n34268) );
  DFFARX1 \s2/msel/arb2/state_reg[2]  ( .D(n17968), .CLK(clock), .RSTB(n34693), 
        .Q(\s2/msel/gnt_p2 [2]), .QN(n34391) );
  DFFARX1 \s1/msel/arb1/state_reg[0]  ( .D(n18000), .CLK(clock), .RSTB(n34691), 
        .Q(\s1/msel/gnt_p1 [0]), .QN(n34673) );
  DFFARX1 \s1/msel/arb1/state_reg[1]  ( .D(n18001), .CLK(clock), .RSTB(n34680), 
        .Q(\s1/msel/gnt_p1 [1]), .QN(n34392) );
  DFFARX1 \s1/msel/arb1/state_reg[2]  ( .D(n18002), .CLK(clock), .RSTB(n34682), 
        .Q(\s1/msel/gnt_p1 [2]), .QN(n34446) );
  DFFARX1 \s1/msel/arb0/state_reg[0]  ( .D(n17997), .CLK(clock), .RSTB(n34677), 
        .Q(\s1/msel/gnt_p0 [0]), .QN(n34233) );
  DFFARX1 \s1/msel/arb0/state_reg[1]  ( .D(n17998), .CLK(clock), .RSTB(n34683), 
        .Q(\s1/msel/gnt_p0 [1]), .QN(n34285) );
  DFFARX1 \s1/msel/arb0/state_reg[2]  ( .D(n17999), .CLK(clock), .RSTB(n34694), 
        .Q(\s1/msel/gnt_p0 [2]), .QN(n34454) );
  DFFARX1 \s1/msel/arb3/state_reg[0]  ( .D(n18003), .CLK(clock), .RSTB(n34684), 
        .Q(\s1/msel/gnt_p3 [0]), .QN(n34280) );
  DFFARX1 \s1/msel/arb3/state_reg[1]  ( .D(n18004), .CLK(clock), .RSTB(n34692), 
        .Q(\s1/msel/gnt_p3 [1]), .QN(n34427) );
  DFFARX1 \s1/msel/arb3/state_reg[2]  ( .D(n18005), .CLK(clock), .RSTB(n34684), 
        .Q(\s1/msel/gnt_p3 [2]), .QN(n34428) );
  DFFARX1 \s1/msel/arb2/state_reg[0]  ( .D(n17994), .CLK(clock), .RSTB(n34686), 
        .Q(\s1/msel/gnt_p2 [0]), .QN(n34385) );
  DFFARX1 \s1/msel/arb2/state_reg[1]  ( .D(n17995), .CLK(clock), .RSTB(n34694), 
        .Q(\s1/msel/gnt_p2 [1]), .QN(n34445) );
  DFFARX1 \s1/msel/arb2/state_reg[2]  ( .D(n17996), .CLK(clock), .RSTB(n34679), 
        .Q(\s1/msel/gnt_p2 [2]), .QN(n34437) );
  DFFARX1 \s3/msel/arb1/state_reg[0]  ( .D(n17944), .CLK(clock), .RSTB(n34695), 
        .Q(\s3/msel/gnt_p1 [0]), .QN(n34658) );
  DFFARX1 \s3/msel/arb1/state_reg[1]  ( .D(n17945), .CLK(clock), .RSTB(n34696), 
        .Q(\s3/msel/gnt_p1 [1]), .QN(n34388) );
  DFFARX1 \s3/msel/arb1/state_reg[2]  ( .D(n17946), .CLK(clock), .RSTB(n34683), 
        .Q(\s3/msel/gnt_p1 [2]), .QN(n34418) );
  DFFARX1 \s3/msel/arb0/state_reg[0]  ( .D(n17941), .CLK(clock), .RSTB(n34697), 
        .Q(\s3/msel/gnt_p0 [0]), .QN(n34393) );
  DFFARX1 \s3/msel/arb0/state_reg[1]  ( .D(n17942), .CLK(clock), .RSTB(n34684), 
        .Q(\s3/msel/gnt_p0 [1]), .QN(n34263) );
  DFFARX1 \s3/msel/arb0/state_reg[2]  ( .D(n17943), .CLK(clock), .RSTB(n34693), 
        .Q(\s3/msel/gnt_p0 [2]), .QN(n34413) );
  DFFARX1 \s3/msel/arb3/state_reg[0]  ( .D(n17947), .CLK(clock), .RSTB(n34687), 
        .Q(\s3/msel/gnt_p3 [0]), .QN(n34665) );
  DFFARX1 \s3/msel/arb3/state_reg[1]  ( .D(n17948), .CLK(clock), .RSTB(n34680), 
        .Q(\s3/msel/gnt_p3 [1]), .QN(n34404) );
  DFFARX1 \s3/msel/arb3/state_reg[2]  ( .D(n17949), .CLK(clock), .RSTB(n34680), 
        .Q(\s3/msel/gnt_p3 [2]), .QN(n34458) );
  DFFARX1 \s3/msel/arb2/state_reg[0]  ( .D(n17938), .CLK(clock), .RSTB(n34680), 
        .Q(\s3/msel/gnt_p2 [0]), .QN(n34416) );
  DFFARX1 \s3/msel/arb2/state_reg[1]  ( .D(n17939), .CLK(clock), .RSTB(n34680), 
        .Q(\s3/msel/gnt_p2 [1]), .QN(n34287) );
  DFFARX1 \s3/msel/arb2/state_reg[2]  ( .D(n17940), .CLK(clock), .RSTB(n34680), 
        .Q(\s3/msel/gnt_p2 [2]), .QN(n34650) );
  DFFARX1 \s4/msel/arb1/state_reg[0]  ( .D(n17916), .CLK(clock), .RSTB(n34680), 
        .Q(\s4/msel/gnt_p1 [0]), .QN(n34246) );
  DFFARX1 \s4/msel/arb1/state_reg[1]  ( .D(n17917), .CLK(clock), .RSTB(n34680), 
        .Q(\s4/msel/gnt_p1 [1]), .QN(n34389) );
  DFFARX1 \s4/msel/arb1/state_reg[2]  ( .D(n17918), .CLK(clock), .RSTB(n34680), 
        .Q(\s4/msel/gnt_p1 [2]), .QN(n34459) );
  DFFARX1 \s4/msel/arb0/state_reg[0]  ( .D(n17913), .CLK(clock), .RSTB(n34691), 
        .Q(\s4/msel/gnt_p0 [0]), .QN(n34378) );
  DFFARX1 \s4/msel/arb0/state_reg[1]  ( .D(n17914), .CLK(clock), .RSTB(n34680), 
        .Q(\s4/msel/gnt_p0 [1]), .QN(n34232) );
  DFFARX1 \s4/msel/arb0/state_reg[2]  ( .D(n17915), .CLK(clock), .RSTB(n34682), 
        .Q(\s4/msel/gnt_p0 [2]), .QN(n34457) );
  DFFARX1 \s4/msel/arb3/state_reg[0]  ( .D(n17919), .CLK(clock), .RSTB(n34678), 
        .Q(\s4/msel/gnt_p3 [0]), .QN(n34455) );
  DFFARX1 \s4/msel/arb3/state_reg[1]  ( .D(n17920), .CLK(clock), .RSTB(n34683), 
        .Q(\s4/msel/gnt_p3 [1]), .QN(n34656) );
  DFFARX1 \s4/msel/arb3/state_reg[2]  ( .D(n17921), .CLK(clock), .RSTB(n34686), 
        .Q(\s4/msel/gnt_p3 [2]), .QN(n34465) );
  DFFARX1 \s4/msel/arb2/state_reg[0]  ( .D(n17910), .CLK(clock), .RSTB(n34684), 
        .Q(\s4/msel/gnt_p2 [0]), .QN(n34408) );
  DFFARX1 \s4/msel/arb2/state_reg[1]  ( .D(n17911), .CLK(clock), .RSTB(n34682), 
        .Q(\s4/msel/gnt_p2 [1]), .QN(n34279) );
  DFFARX1 \s4/msel/arb2/state_reg[2]  ( .D(n17912), .CLK(clock), .RSTB(n34685), 
        .Q(\s4/msel/gnt_p2 [2]), .QN(n34607) );
  DFFARX1 \s6/msel/arb1/state_reg[0]  ( .D(n17860), .CLK(clock), .RSTB(n34686), 
        .Q(\s6/msel/gnt_p1 [0]), .QN(n34243) );
  DFFARX1 \s6/msel/arb1/state_reg[1]  ( .D(n17861), .CLK(clock), .RSTB(n34678), 
        .Q(\s6/msel/gnt_p1 [1]), .QN(n34666) );
  DFFARX1 \s6/msel/arb1/state_reg[2]  ( .D(n17862), .CLK(clock), .RSTB(n34677), 
        .Q(\s6/msel/gnt_p1 [2]), .QN(n34597) );
  DFFARX1 \s6/msel/arb0/state_reg[0]  ( .D(n17857), .CLK(clock), .RSTB(n34696), 
        .Q(\s6/msel/gnt_p0 [0]), .QN(n34671) );
  DFFARX1 \s6/msel/arb0/state_reg[1]  ( .D(n17858), .CLK(clock), .RSTB(n34682), 
        .Q(\s6/msel/gnt_p0 [1]), .QN(n34675) );
  DFFARX1 \s6/msel/arb0/state_reg[2]  ( .D(n17859), .CLK(clock), .RSTB(n34697), 
        .Q(\s6/msel/gnt_p0 [2]), .QN(n34402) );
  DFFARX1 \s6/msel/arb3/state_reg[0]  ( .D(n17863), .CLK(clock), .RSTB(n34683), 
        .Q(\s6/msel/gnt_p3 [0]), .QN(n34449) );
  DFFARX1 \s6/msel/arb3/state_reg[1]  ( .D(n17864), .CLK(clock), .RSTB(n34693), 
        .Q(\s6/msel/gnt_p3 [1]), .QN(n34270) );
  DFFARX1 \s6/msel/arb3/state_reg[2]  ( .D(n17865), .CLK(clock), .RSTB(n34681), 
        .Q(\s6/msel/gnt_p3 [2]), .QN(n34640) );
  DFFARX1 \s6/msel/arb2/state_reg[0]  ( .D(n17854), .CLK(clock), .RSTB(n34687), 
        .Q(\s6/msel/gnt_p2 [0]), .QN(n34224) );
  DFFARX1 \s6/msel/arb2/state_reg[1]  ( .D(n17855), .CLK(clock), .RSTB(n34680), 
        .Q(\s6/msel/gnt_p2 [1]), .QN(n34254) );
  DFFARX1 \s6/msel/arb2/state_reg[2]  ( .D(n17856), .CLK(clock), .RSTB(n34688), 
        .Q(\s6/msel/gnt_p2 [2]), .QN(n34461) );
  DFFARX1 \s5/msel/arb1/state_reg[0]  ( .D(n17888), .CLK(clock), .RSTB(n34689), 
        .Q(\s5/msel/gnt_p1 [0]), .QN(n34657) );
  DFFARX1 \s5/msel/arb1/state_reg[1]  ( .D(n17889), .CLK(clock), .RSTB(n34690), 
        .Q(\s5/msel/gnt_p1 [1]), .QN(n34252) );
  DFFARX1 \s5/msel/arb1/state_reg[2]  ( .D(n17890), .CLK(clock), .RSTB(n34691), 
        .Q(\s5/msel/gnt_p1 [2]), .QN(n34371) );
  DFFARX1 \s5/msel/arb0/state_reg[0]  ( .D(n17885), .CLK(clock), .RSTB(n34683), 
        .Q(\s5/msel/gnt_p0 [0]), .QN(n34398) );
  DFFARX1 \s5/msel/arb0/state_reg[1]  ( .D(n17886), .CLK(clock), .RSTB(n34678), 
        .Q(\s5/msel/gnt_p0 [1]), .QN(n34415) );
  DFFARX1 \s5/msel/arb0/state_reg[2]  ( .D(n17887), .CLK(clock), .RSTB(n34677), 
        .Q(\s5/msel/gnt_p0 [2]), .QN(n34258) );
  DFFARX1 \s5/msel/arb3/state_reg[0]  ( .D(n17891), .CLK(clock), .RSTB(n34685), 
        .Q(\s5/msel/gnt_p3 [0]), .QN(n34409) );
  DFFARX1 \s5/msel/arb3/state_reg[1]  ( .D(n17892), .CLK(clock), .RSTB(n34692), 
        .Q(\s5/msel/gnt_p3 [1]), .QN(n34227) );
  DFFARX1 \s5/msel/arb3/state_reg[2]  ( .D(n17893), .CLK(clock), .RSTB(n34682), 
        .Q(\s5/msel/gnt_p3 [2]), .QN(n34275) );
  DFFARX1 \s5/msel/arb2/state_reg[0]  ( .D(n17882), .CLK(clock), .RSTB(n34686), 
        .Q(\s5/msel/gnt_p2 [0]), .QN(n34256) );
  DFFARX1 \s5/msel/arb2/state_reg[1]  ( .D(n17883), .CLK(clock), .RSTB(n34694), 
        .Q(\s5/msel/gnt_p2 [1]), .QN(n34396) );
  DFFARX1 \s5/msel/arb2/state_reg[2]  ( .D(n17884), .CLK(clock), .RSTB(n34679), 
        .Q(\s5/msel/gnt_p2 [2]), .QN(n34426) );
  DFFARX1 \s7/msel/arb1/state_reg[0]  ( .D(n17832), .CLK(clock), .RSTB(n34695), 
        .Q(\s7/msel/gnt_p1 [0]), .QN(n34245) );
  DFFARX1 \s7/msel/arb1/state_reg[1]  ( .D(n17833), .CLK(clock), .RSTB(n34696), 
        .Q(\s7/msel/gnt_p1 [1]), .QN(n34439) );
  DFFARX1 \s7/msel/arb1/state_reg[2]  ( .D(n17834), .CLK(clock), .RSTB(n34680), 
        .Q(\s7/msel/gnt_p1 [2]), .QN(n34424) );
  DFFARX1 \s7/msel/arb0/state_reg[0]  ( .D(n17829), .CLK(clock), .RSTB(n34691), 
        .Q(\s7/msel/gnt_p0 [0]), .QN(n34289) );
  DFFARX1 \s7/msel/arb0/state_reg[1]  ( .D(n17830), .CLK(clock), .RSTB(n34680), 
        .Q(\s7/msel/gnt_p0 [1]), .QN(n34414) );
  DFFARX1 \s7/msel/arb0/state_reg[2]  ( .D(n17831), .CLK(clock), .RSTB(n34682), 
        .Q(\s7/msel/gnt_p0 [2]), .QN(n34550) );
  DFFARX1 \s7/msel/arb3/state_reg[0]  ( .D(n17835), .CLK(clock), .RSTB(n34685), 
        .Q(\s7/msel/gnt_p3 [0]), .QN(n34410) );
  DFFARX1 \s7/msel/arb3/state_reg[1]  ( .D(n17836), .CLK(clock), .RSTB(n34683), 
        .Q(\s7/msel/gnt_p3 [1]), .QN(n34262) );
  DFFARX1 \s7/msel/arb3/state_reg[2]  ( .D(n17837), .CLK(clock), .RSTB(n34692), 
        .Q(\s7/msel/gnt_p3 [2]), .QN(n34380) );
  DFFARX1 \s7/msel/arb2/state_reg[0]  ( .D(n17826), .CLK(clock), .RSTB(n34684), 
        .Q(\s7/msel/gnt_p2 [0]), .QN(n34429) );
  DFFARX1 \s7/msel/arb2/state_reg[1]  ( .D(n17827), .CLK(clock), .RSTB(n34685), 
        .Q(\s7/msel/gnt_p2 [1]), .QN(n34274) );
  DFFARX1 \s7/msel/arb2/state_reg[2]  ( .D(n17828), .CLK(clock), .RSTB(n34690), 
        .Q(\s7/msel/gnt_p2 [2]), .QN(n34435) );
  DFFARX1 \s8/msel/arb1/state_reg[0]  ( .D(n17804), .CLK(clock), .RSTB(n34678), 
        .Q(\s8/msel/gnt_p1 [0]), .QN(n34229) );
  DFFARX1 \s8/msel/arb1/state_reg[1]  ( .D(n17805), .CLK(clock), .RSTB(n34677), 
        .Q(\s8/msel/gnt_p1 [1]), .QN(n34276) );
  DFFARX1 \s8/msel/arb1/state_reg[2]  ( .D(n17806), .CLK(clock), .RSTB(n34684), 
        .Q(\s8/msel/gnt_p1 [2]), .QN(n34420) );
  DFFARX1 \s8/msel/arb0/state_reg[0]  ( .D(n17801), .CLK(clock), .RSTB(n34680), 
        .Q(\s8/msel/gnt_p0 [0]) );
  DFFARX1 \s8/msel/arb0/state_reg[1]  ( .D(n17802), .CLK(clock), .RSTB(n34693), 
        .Q(\s8/msel/gnt_p0 [1]), .QN(n34654) );
  DFFARX1 \s8/msel/arb0/state_reg[2]  ( .D(n17803), .CLK(clock), .RSTB(n34681), 
        .Q(\s8/msel/gnt_p0 [2]), .QN(n34403) );
  DFFARX1 \s8/msel/arb3/state_reg[0]  ( .D(n17807), .CLK(clock), .RSTB(n34687), 
        .Q(\s8/msel/gnt_p3 [0]), .QN(n34228) );
  DFFARX1 \s8/msel/arb3/state_reg[1]  ( .D(n17808), .CLK(clock), .RSTB(n34688), 
        .Q(\s8/msel/gnt_p3 [1]), .QN(n34223) );
  DFFARX1 \s8/msel/arb3/state_reg[2]  ( .D(n17809), .CLK(clock), .RSTB(n34689), 
        .Q(\s8/msel/gnt_p3 [2]), .QN(n34456) );
  DFFARX1 \s8/msel/arb2/state_reg[0]  ( .D(n17798), .CLK(clock), .RSTB(n34690), 
        .Q(\s8/msel/gnt_p2 [0]), .QN(n34467) );
  DFFARX1 \s8/msel/arb2/state_reg[1]  ( .D(n17799), .CLK(clock), .RSTB(n34691), 
        .Q(\s8/msel/gnt_p2 [1]), .QN(n34273) );
  DFFARX1 \s8/msel/arb2/state_reg[2]  ( .D(n17800), .CLK(clock), .RSTB(n34680), 
        .Q(\s8/msel/gnt_p2 [2]), .QN(n34430) );
  DFFARX1 \s10/msel/arb1/state_reg[0]  ( .D(n17748), .CLK(clock), .RSTB(n34682), .Q(\s10/msel/gnt_p1 [0]), .QN(n34434) );
  DFFARX1 \s10/msel/arb1/state_reg[1]  ( .D(n17749), .CLK(clock), .RSTB(n34684), .Q(\s10/msel/gnt_p1 [1]), .QN(n34253) );
  DFFARX1 \s10/msel/arb1/state_reg[2]  ( .D(n17750), .CLK(clock), .RSTB(n34683), .Q(\s10/msel/gnt_p1 [2]), .QN(n34610) );
  DFFARX1 \s10/msel/arb0/state_reg[0]  ( .D(n17745), .CLK(clock), .RSTB(n34679), .Q(\s10/msel/gnt_p0 [0]), .QN(n34417) );
  DFFARX1 \s10/msel/arb0/state_reg[1]  ( .D(n17746), .CLK(clock), .RSTB(n34695), .Q(\s10/msel/gnt_p0 [1]), .QN(n34257) );
  DFFARX1 \s10/msel/arb0/state_reg[2]  ( .D(n17747), .CLK(clock), .RSTB(n34696), .Q(\s10/msel/gnt_p0 [2]), .QN(n34451) );
  DFFARX1 \s10/msel/arb3/state_reg[0]  ( .D(n17751), .CLK(clock), .RSTB(n34690), .Q(\s10/msel/gnt_p3 [0]), .QN(n34464) );
  DFFARX1 \s10/msel/arb3/state_reg[1]  ( .D(n17752), .CLK(clock), .RSTB(n34697), .Q(\s10/msel/gnt_p3 [1]), .QN(n34251) );
  DFFARX1 \s10/msel/arb3/state_reg[2]  ( .D(n17753), .CLK(clock), .RSTB(n34693), .Q(\s10/msel/gnt_p3 [2]), .QN(n34472) );
  DFFARX1 \s10/msel/arb2/state_reg[0]  ( .D(n17742), .CLK(clock), .RSTB(n34681), .Q(\s10/msel/gnt_p2 [0]), .QN(n34463) );
  DFFARX1 \s10/msel/arb2/state_reg[1]  ( .D(n17743), .CLK(clock), .RSTB(n34687), .Q(\s10/msel/gnt_p2 [1]), .QN(n34255) );
  DFFARX1 \s10/msel/arb2/state_reg[2]  ( .D(n17744), .CLK(clock), .RSTB(n34688), .Q(\s10/msel/gnt_p2 [2]), .QN(n34405) );
  DFFARX1 \s9/msel/arb1/state_reg[0]  ( .D(n17776), .CLK(clock), .RSTB(n34689), 
        .Q(\s9/msel/gnt_p1 [0]), .QN(n34260) );
  DFFARX1 \s9/msel/arb1/state_reg[1]  ( .D(n17777), .CLK(clock), .RSTB(n34690), 
        .Q(\s9/msel/gnt_p1 [1]), .QN(n34400) );
  DFFARX1 \s9/msel/arb1/state_reg[2]  ( .D(n17778), .CLK(clock), .RSTB(n34692), 
        .Q(\s9/msel/gnt_p1 [2]), .QN(n34442) );
  DFFARX1 \s9/msel/arb0/state_reg[0]  ( .D(n17773), .CLK(clock), .RSTB(n34690), 
        .Q(\s9/msel/gnt_p0 [0]), .QN(n34436) );
  DFFARX1 \s9/msel/arb0/state_reg[1]  ( .D(n17774), .CLK(clock), .RSTB(n34686), 
        .Q(\s9/msel/gnt_p0 [1]), .QN(n34266) );
  DFFARX1 \s9/msel/arb0/state_reg[2]  ( .D(n17775), .CLK(clock), .RSTB(n34694), 
        .Q(\s9/msel/gnt_p0 [2]), .QN(n34284) );
  DFFARX1 \s9/msel/arb3/state_reg[0]  ( .D(n17779), .CLK(clock), .RSTB(n34679), 
        .Q(\s9/msel/gnt_p3 [0]), .QN(n34282) );
  DFFARX1 \s9/msel/arb3/state_reg[1]  ( .D(n17780), .CLK(clock), .RSTB(n34695), 
        .Q(\s9/msel/gnt_p3 [1]), .QN(n34225) );
  DFFARX1 \s9/msel/arb3/state_reg[2]  ( .D(n17781), .CLK(clock), .RSTB(n34696), 
        .Q(\s9/msel/gnt_p3 [2]), .QN(n34560) );
  DFFARX1 \s9/msel/arb2/state_reg[0]  ( .D(n17770), .CLK(clock), .RSTB(n34689), 
        .Q(\s9/msel/gnt_p2 [0]), .QN(n34462) );
  DFFARX1 \s9/msel/arb2/state_reg[1]  ( .D(n17771), .CLK(clock), .RSTB(n34697), 
        .Q(\s9/msel/gnt_p2 [1]), .QN(n34466) );
  DFFARX1 \s9/msel/arb2/state_reg[2]  ( .D(n17772), .CLK(clock), .RSTB(n34693), 
        .Q(\s9/msel/gnt_p2 [2]), .QN(n34469) );
  DFFARX1 \s13/msel/arb1/state_reg[0]  ( .D(n17664), .CLK(clock), .RSTB(n34681), .Q(\s13/msel/gnt_p1 [0]), .QN(n34248) );
  DFFARX1 \s13/msel/arb1/state_reg[1]  ( .D(n17665), .CLK(clock), .RSTB(n34687), .Q(\s13/msel/gnt_p1 [1]), .QN(n34411) );
  DFFARX1 \s13/msel/arb1/state_reg[2]  ( .D(n17666), .CLK(clock), .RSTB(n34680), .Q(\s13/msel/gnt_p1 [2]), .QN(n34471) );
  DFFARX1 \s13/msel/arb0/state_reg[0]  ( .D(n17661), .CLK(clock), .RSTB(n34692), .Q(\s13/msel/gnt_p0 [0]), .QN(n34653) );
  DFFARX1 \s13/msel/arb0/state_reg[1]  ( .D(n17662), .CLK(clock), .RSTB(n34689), .Q(\s13/msel/gnt_p0 [1]), .QN(n34264) );
  DFFARX1 \s13/msel/arb0/state_reg[2]  ( .D(n17663), .CLK(clock), .RSTB(n34686), .Q(\s13/msel/gnt_p0 [2]), .QN(n34292) );
  DFFARX1 \s13/msel/arb3/state_reg[0]  ( .D(n17667), .CLK(clock), .RSTB(n34688), .Q(\s13/msel/gnt_p3 [0]), .QN(n34267) );
  DFFARX1 \s13/msel/arb3/state_reg[1]  ( .D(n17668), .CLK(clock), .RSTB(n34694), .Q(\s13/msel/gnt_p3 [1]), .QN(n34384) );
  DFFARX1 \s13/msel/arb3/state_reg[2]  ( .D(n17669), .CLK(clock), .RSTB(n34679), .Q(\s13/msel/gnt_p3 [2]), .QN(n34431) );
  DFFARX1 \s13/msel/arb2/state_reg[0]  ( .D(n17658), .CLK(clock), .RSTB(n34695), .Q(\s13/msel/gnt_p2 [0]), .QN(n34288) );
  DFFARX1 \s13/msel/arb2/state_reg[1]  ( .D(n17659), .CLK(clock), .RSTB(n34696), .Q(\s13/msel/gnt_p2 [1]), .QN(n34234) );
  DFFARX1 \s13/msel/arb2/state_reg[2]  ( .D(n17660), .CLK(clock), .RSTB(n34697), .Q(\s13/msel/gnt_p2 [2]), .QN(n34608) );
  DFFARX1 \s12/msel/arb1/state_reg[0]  ( .D(n17692), .CLK(clock), .RSTB(n34693), .Q(\s12/msel/gnt_p1 [0]), .QN(n34664) );
  DFFARX1 \s12/msel/arb1/state_reg[1]  ( .D(n17693), .CLK(clock), .RSTB(n34681), .Q(\s12/msel/gnt_p1 [1]), .QN(n34545) );
  DFFARX1 \s12/msel/arb1/state_reg[2]  ( .D(n17694), .CLK(clock), .RSTB(n34679), .Q(\s12/msel/gnt_p1 [2]), .QN(n34397) );
  DFFARX1 \s12/msel/arb0/state_reg[0]  ( .D(n17689), .CLK(clock), .RSTB(n34679), .Q(\s12/msel/gnt_p0 [0]), .QN(n34443) );
  DFFARX1 \s12/msel/arb0/state_reg[1]  ( .D(n17690), .CLK(clock), .RSTB(n34679), .Q(\s12/msel/gnt_p0 [1]), .QN(n34278) );
  DFFARX1 \s12/msel/arb0/state_reg[2]  ( .D(n17691), .CLK(clock), .RSTB(n34679), .Q(\s12/msel/gnt_p0 [2]), .QN(n34382) );
  DFFARX1 \s12/msel/arb3/state_reg[0]  ( .D(n17695), .CLK(clock), .RSTB(n34679), .Q(\s12/msel/gnt_p3 [0]), .QN(n34269) );
  DFFARX1 \s12/msel/arb3/state_reg[1]  ( .D(n17696), .CLK(clock), .RSTB(n34679), .Q(\s12/msel/gnt_p3 [1]), .QN(n34230) );
  DFFARX1 \s12/msel/arb3/state_reg[2]  ( .D(n17697), .CLK(clock), .RSTB(n34679), .Q(\s12/msel/gnt_p3 [2]), .QN(n34450) );
  DFFARX1 \s12/msel/arb2/state_reg[0]  ( .D(n17686), .CLK(clock), .RSTB(n34679), .Q(\s12/msel/gnt_p2 [0]), .QN(n34244) );
  DFFARX1 \s12/msel/arb2/state_reg[1]  ( .D(n17687), .CLK(clock), .RSTB(n34679), .Q(\s12/msel/gnt_p2 [1]), .QN(n34422) );
  DFFARX1 \s12/msel/arb2/state_reg[2]  ( .D(n17688), .CLK(clock), .RSTB(n34679), .Q(\s12/msel/gnt_p2 [2]), .QN(n34553) );
  DFFARX1 \s14/msel/arb1/state_reg[0]  ( .D(n17636), .CLK(clock), .RSTB(n34679), .Q(\s14/msel/gnt_p1 [0]), .QN(n34394) );
  DFFARX1 \s14/msel/arb1/state_reg[1]  ( .D(n17637), .CLK(clock), .RSTB(n34679), .Q(\s14/msel/gnt_p1 [1]), .QN(n34242) );
  DFFARX1 \s14/msel/arb1/state_reg[2]  ( .D(n17638), .CLK(clock), .RSTB(n34692), .Q(\s14/msel/gnt_p1 [2]), .QN(n34386) );
  DFFARX1 \s14/msel/arb0/state_reg[0]  ( .D(n17633), .CLK(clock), .RSTB(n34686), .Q(\s14/msel/gnt_p0 [0]), .QN(n34639) );
  DFFARX1 \s14/msel/arb0/state_reg[1]  ( .D(n17634), .CLK(clock), .RSTB(n34687), .Q(\s14/msel/gnt_p0 [1]), .QN(n34247) );
  DFFARX1 \s14/msel/arb0/state_reg[2]  ( .D(n17635), .CLK(clock), .RSTB(n34688), .Q(\s14/msel/gnt_p0 [2]), .QN(n34387) );
  DFFARX1 \s14/msel/arb3/state_reg[0]  ( .D(n17639), .CLK(clock), .RSTB(n34694), .Q(\s14/msel/gnt_p3 [0]), .QN(n34468) );
  DFFARX1 \s14/msel/arb3/state_reg[1]  ( .D(n17640), .CLK(clock), .RSTB(n34679), .Q(\s14/msel/gnt_p3 [1]), .QN(n34447) );
  DFFARX1 \s14/msel/arb3/state_reg[2]  ( .D(n17641), .CLK(clock), .RSTB(n34695), .Q(\s14/msel/gnt_p3 [2]), .QN(n34281) );
  DFFARX1 \s14/msel/arb2/state_reg[0]  ( .D(n17630), .CLK(clock), .RSTB(n34696), .Q(\s14/msel/gnt_p2 [0]), .QN(n34271) );
  DFFARX1 \s14/msel/arb2/state_reg[1]  ( .D(n17631), .CLK(clock), .RSTB(n34697), .Q(\s14/msel/gnt_p2 [1]), .QN(n34381) );
  DFFARX1 \s14/msel/arb2/state_reg[2]  ( .D(n17632), .CLK(clock), .RSTB(n34693), .Q(\s14/msel/gnt_p2 [2]), .QN(n34460) );
  DFFARX1 \s11/msel/arb1/state_reg[0]  ( .D(n17720), .CLK(clock), .RSTB(n34681), .Q(\s11/msel/gnt_p1 [0]), .QN(n34655) );
  DFFARX1 \s11/msel/arb1/state_reg[1]  ( .D(n17721), .CLK(clock), .RSTB(n34689), .Q(\s11/msel/gnt_p1 [1]), .QN(n34390) );
  DFFARX1 \s11/msel/arb1/state_reg[2]  ( .D(n17722), .CLK(clock), .RSTB(n34678), .Q(\s11/msel/gnt_p1 [2]), .QN(n34425) );
  DFFARX1 \s11/msel/arb0/state_reg[0]  ( .D(n17717), .CLK(clock), .RSTB(n34678), .Q(\s11/msel/gnt_p0 [0]), .QN(n34249) );
  DFFARX1 \s11/msel/arb0/state_reg[1]  ( .D(n17718), .CLK(clock), .RSTB(n34678), .Q(\s11/msel/gnt_p0 [1]), .QN(n34668) );
  DFFARX1 \s11/msel/arb0/state_reg[2]  ( .D(n17719), .CLK(clock), .RSTB(n34678), .Q(\s11/msel/gnt_p0 [2]), .QN(n34452) );
  DFFARX1 \s11/msel/arb3/state_reg[0]  ( .D(n17723), .CLK(clock), .RSTB(n34678), .Q(\s11/msel/gnt_p3 [0]), .QN(n34399) );
  DFFARX1 \s11/msel/arb3/state_reg[1]  ( .D(n17724), .CLK(clock), .RSTB(n34678), .Q(\s11/msel/gnt_p3 [1]), .QN(n34419) );
  DFFARX1 \s11/msel/arb3/state_reg[2]  ( .D(n17725), .CLK(clock), .RSTB(n34678), .Q(\s11/msel/gnt_p3 [2]), .QN(n34444) );
  DFFARX1 \s11/msel/arb2/state_reg[0]  ( .D(n17714), .CLK(clock), .RSTB(n34678), .Q(\s11/msel/gnt_p2 [0]), .QN(n34470) );
  DFFARX1 \s11/msel/arb2/state_reg[1]  ( .D(n17715), .CLK(clock), .RSTB(n34678), .Q(\s11/msel/gnt_p2 [1]), .QN(n34407) );
  DFFARX1 \s11/msel/arb2/state_reg[2]  ( .D(n17716), .CLK(clock), .RSTB(n34678), .Q(\s11/msel/gnt_p2 [2]), .QN(n34401) );
  DFFARX1 \s15/msel/arb1/state_reg[0]  ( .D(n17608), .CLK(clock), .RSTB(n34678), .Q(\s15/msel/gnt_p1 [0]), .QN(n34272) );
  DFFARX1 \s15/msel/arb1/state_reg[1]  ( .D(n17609), .CLK(clock), .RSTB(n34678), .Q(\s15/msel/gnt_p1 [1]), .QN(n34412) );
  DFFARX1 \s15/msel/arb1/state_reg[2]  ( .D(n17610), .CLK(clock), .RSTB(n34697), .Q(\s15/msel/gnt_p1 [2]), .QN(n34448) );
  DFFARX1 \s15/msel/arb0/state_reg[0]  ( .D(n17605), .CLK(clock), .RSTB(n34688), .Q(\s15/msel/gnt_p0 [0]), .QN(n34261) );
  DFFARX1 \s15/msel/arb0/state_reg[1]  ( .D(n17606), .CLK(clock), .RSTB(n34679), .Q(\s15/msel/gnt_p0 [1]), .QN(n34226) );
  DFFARX1 \s15/msel/arb0/state_reg[2]  ( .D(n17607), .CLK(clock), .RSTB(n34689), .Q(\s15/msel/gnt_p0 [2]), .QN(n34441) );
  DFFARX1 \s15/msel/arb3/state_reg[0]  ( .D(n17611), .CLK(clock), .RSTB(n34690), .Q(\s15/msel/gnt_p3 [0]), .QN(n34283) );
  DFFARX1 \s15/msel/arb3/state_reg[1]  ( .D(n17612), .CLK(clock), .RSTB(n34689), .Q(\s15/msel/gnt_p3 [1]), .QN(n34421) );
  DFFARX1 \s15/msel/arb3/state_reg[2]  ( .D(n17613), .CLK(clock), .RSTB(n34677), .Q(\s15/msel/gnt_p3 [2]), .QN(n34433) );
  DFFARX1 \s15/msel/arb2/state_reg[0]  ( .D(n17601), .CLK(clock), .RSTB(n34691), .Q(\s15/msel/gnt_p2 [0]), .QN(n34231) );
  DFFARX1 \s15/msel/arb2/state_reg[1]  ( .D(n17603), .CLK(clock), .RSTB(n34681), .Q(\s15/msel/gnt_p2 [1]), .QN(n34265) );
  DFFARX1 \s15/msel/arb2/state_reg[2]  ( .D(n17604), .CLK(clock), .RSTB(n34680), .Q(\s15/msel/gnt_p2 [2]), .QN(n34406) );
  DFFX1 \s0/m7_cyc_r_reg  ( .D(m7s0_cyc), .CLK(clock), .Q(\s0/m7_cyc_r ) );
  DFFX1 \s0/m6_cyc_r_reg  ( .D(m6s0_cyc), .CLK(clock), .Q(\s0/m6_cyc_r ) );
  DFFX1 \s0/m5_cyc_r_reg  ( .D(m5s0_cyc), .CLK(clock), .Q(\s0/m5_cyc_r ) );
  DFFX1 \s0/m4_cyc_r_reg  ( .D(m4s0_cyc), .CLK(clock), .Q(\s0/m4_cyc_r ) );
  DFFX1 \s0/m3_cyc_r_reg  ( .D(m3s0_cyc), .CLK(clock), .Q(\s0/m3_cyc_r ) );
  DFFX1 \s0/m2_cyc_r_reg  ( .D(m2s0_cyc), .CLK(clock), .Q(\s0/m2_cyc_r ) );
  DFFX1 \s0/m1_cyc_r_reg  ( .D(m1s0_cyc), .CLK(clock), .Q(\s0/m1_cyc_r ) );
  DFFX1 \s0/m0_cyc_r_reg  ( .D(m0s0_cyc), .CLK(clock), .Q(\s0/m0_cyc_r ) );
  DFFX1 \s0/next_reg  ( .D(n18193), .CLK(clock), .Q(\s0/next ) );
  DFFX1 \s1/m7_cyc_r_reg  ( .D(m7s1_cyc), .CLK(clock), .Q(\s1/m7_cyc_r ) );
  DFFX1 \s1/m6_cyc_r_reg  ( .D(m6s1_cyc), .CLK(clock), .Q(\s1/m6_cyc_r ) );
  DFFX1 \s1/m5_cyc_r_reg  ( .D(m5s1_cyc), .CLK(clock), .Q(\s1/m5_cyc_r ) );
  DFFX1 \s1/m4_cyc_r_reg  ( .D(m4s1_cyc), .CLK(clock), .Q(\s1/m4_cyc_r ) );
  DFFX1 \s1/m3_cyc_r_reg  ( .D(m3s1_cyc), .CLK(clock), .Q(\s1/m3_cyc_r ) );
  DFFX1 \s1/m2_cyc_r_reg  ( .D(m2s1_cyc), .CLK(clock), .Q(\s1/m2_cyc_r ) );
  DFFX1 \s1/m1_cyc_r_reg  ( .D(m1s1_cyc), .CLK(clock), .Q(\s1/m1_cyc_r ) );
  DFFX1 \s1/m0_cyc_r_reg  ( .D(m0s1_cyc), .CLK(clock), .Q(\s1/m0_cyc_r ) );
  DFFX1 \s1/next_reg  ( .D(n18192), .CLK(clock), .Q(\s1/next ) );
  DFFX1 \s2/m7_cyc_r_reg  ( .D(m7s2_cyc), .CLK(clock), .Q(\s2/m7_cyc_r ) );
  DFFX1 \s2/m6_cyc_r_reg  ( .D(m6s2_cyc), .CLK(clock), .Q(\s2/m6_cyc_r ) );
  DFFX1 \s2/m5_cyc_r_reg  ( .D(m5s2_cyc), .CLK(clock), .Q(\s2/m5_cyc_r ) );
  DFFX1 \s2/m4_cyc_r_reg  ( .D(m4s2_cyc), .CLK(clock), .Q(\s2/m4_cyc_r ) );
  DFFX1 \s2/m3_cyc_r_reg  ( .D(m3s2_cyc), .CLK(clock), .Q(\s2/m3_cyc_r ) );
  DFFX1 \s2/m2_cyc_r_reg  ( .D(m2s2_cyc), .CLK(clock), .Q(\s2/m2_cyc_r ) );
  DFFX1 \s2/m1_cyc_r_reg  ( .D(m1s2_cyc), .CLK(clock), .Q(\s2/m1_cyc_r ) );
  DFFX1 \s2/m0_cyc_r_reg  ( .D(m0s2_cyc), .CLK(clock), .Q(\s2/m0_cyc_r ) );
  DFFX1 \s2/next_reg  ( .D(n18191), .CLK(clock), .Q(\s2/next ), .QN(n34667) );
  DFFX1 \s3/m7_cyc_r_reg  ( .D(m7s3_cyc), .CLK(clock), .Q(\s3/m7_cyc_r ) );
  DFFX1 \s3/m6_cyc_r_reg  ( .D(m6s3_cyc), .CLK(clock), .Q(\s3/m6_cyc_r ) );
  DFFX1 \s3/m5_cyc_r_reg  ( .D(m5s3_cyc), .CLK(clock), .Q(\s3/m5_cyc_r ) );
  DFFX1 \s3/m4_cyc_r_reg  ( .D(m4s3_cyc), .CLK(clock), .Q(\s3/m4_cyc_r ) );
  DFFX1 \s3/m3_cyc_r_reg  ( .D(m3s3_cyc), .CLK(clock), .Q(\s3/m3_cyc_r ) );
  DFFX1 \s3/m2_cyc_r_reg  ( .D(m2s3_cyc), .CLK(clock), .Q(\s3/m2_cyc_r ) );
  DFFX1 \s3/m1_cyc_r_reg  ( .D(m1s3_cyc), .CLK(clock), .Q(\s3/m1_cyc_r ) );
  DFFX1 \s3/m0_cyc_r_reg  ( .D(m0s3_cyc), .CLK(clock), .Q(\s3/m0_cyc_r ) );
  DFFX1 \s3/next_reg  ( .D(n18190), .CLK(clock), .Q(\s3/next ) );
  DFFX1 \s4/m7_cyc_r_reg  ( .D(m7s4_cyc), .CLK(clock), .Q(\s4/m7_cyc_r ) );
  DFFX1 \s4/m6_cyc_r_reg  ( .D(m6s4_cyc), .CLK(clock), .Q(\s4/m6_cyc_r ) );
  DFFX1 \s4/m5_cyc_r_reg  ( .D(m5s4_cyc), .CLK(clock), .Q(\s4/m5_cyc_r ) );
  DFFX1 \s4/m4_cyc_r_reg  ( .D(m4s4_cyc), .CLK(clock), .Q(\s4/m4_cyc_r ) );
  DFFX1 \s4/m3_cyc_r_reg  ( .D(m3s4_cyc), .CLK(clock), .Q(\s4/m3_cyc_r ) );
  DFFX1 \s4/m2_cyc_r_reg  ( .D(m2s4_cyc), .CLK(clock), .Q(\s4/m2_cyc_r ) );
  DFFX1 \s4/m1_cyc_r_reg  ( .D(m1s4_cyc), .CLK(clock), .Q(\s4/m1_cyc_r ) );
  DFFX1 \s4/m0_cyc_r_reg  ( .D(m0s4_cyc), .CLK(clock), .Q(\s4/m0_cyc_r ) );
  DFFX1 \s4/next_reg  ( .D(n18189), .CLK(clock), .Q(\s4/next ) );
  DFFX1 \s5/m7_cyc_r_reg  ( .D(m7s5_cyc), .CLK(clock), .Q(\s5/m7_cyc_r ) );
  DFFX1 \s5/m6_cyc_r_reg  ( .D(m6s5_cyc), .CLK(clock), .Q(\s5/m6_cyc_r ) );
  DFFX1 \s5/m5_cyc_r_reg  ( .D(m5s5_cyc), .CLK(clock), .Q(\s5/m5_cyc_r ) );
  DFFX1 \s5/m4_cyc_r_reg  ( .D(m4s5_cyc), .CLK(clock), .Q(\s5/m4_cyc_r ) );
  DFFX1 \s5/m3_cyc_r_reg  ( .D(m3s5_cyc), .CLK(clock), .Q(\s5/m3_cyc_r ) );
  DFFX1 \s5/m2_cyc_r_reg  ( .D(m2s5_cyc), .CLK(clock), .Q(\s5/m2_cyc_r ) );
  DFFX1 \s5/m1_cyc_r_reg  ( .D(m1s5_cyc), .CLK(clock), .Q(\s5/m1_cyc_r ) );
  DFFX1 \s5/m0_cyc_r_reg  ( .D(m0s5_cyc), .CLK(clock), .Q(\s5/m0_cyc_r ) );
  DFFX1 \s5/next_reg  ( .D(n18188), .CLK(clock), .Q(\s5/next ) );
  DFFX1 \s6/m7_cyc_r_reg  ( .D(m7s6_cyc), .CLK(clock), .Q(\s6/m7_cyc_r ) );
  DFFX1 \s6/m6_cyc_r_reg  ( .D(m6s6_cyc), .CLK(clock), .Q(\s6/m6_cyc_r ) );
  DFFX1 \s6/m5_cyc_r_reg  ( .D(m5s6_cyc), .CLK(clock), .Q(\s6/m5_cyc_r ) );
  DFFX1 \s6/m4_cyc_r_reg  ( .D(m4s6_cyc), .CLK(clock), .Q(\s6/m4_cyc_r ) );
  DFFX1 \s6/m3_cyc_r_reg  ( .D(m3s6_cyc), .CLK(clock), .Q(\s6/m3_cyc_r ) );
  DFFX1 \s6/m2_cyc_r_reg  ( .D(m2s6_cyc), .CLK(clock), .Q(\s6/m2_cyc_r ) );
  DFFX1 \s6/m1_cyc_r_reg  ( .D(m1s6_cyc), .CLK(clock), .Q(\s6/m1_cyc_r ) );
  DFFX1 \s6/m0_cyc_r_reg  ( .D(m0s6_cyc), .CLK(clock), .Q(\s6/m0_cyc_r ) );
  DFFX1 \s6/next_reg  ( .D(n18187), .CLK(clock), .Q(\s6/next ) );
  DFFX1 \s7/m7_cyc_r_reg  ( .D(m7s7_cyc), .CLK(clock), .Q(\s7/m7_cyc_r ) );
  DFFX1 \s7/m6_cyc_r_reg  ( .D(m6s7_cyc), .CLK(clock), .Q(\s7/m6_cyc_r ) );
  DFFX1 \s7/m5_cyc_r_reg  ( .D(m5s7_cyc), .CLK(clock), .Q(\s7/m5_cyc_r ) );
  DFFX1 \s7/m4_cyc_r_reg  ( .D(m4s7_cyc), .CLK(clock), .Q(\s7/m4_cyc_r ) );
  DFFX1 \s7/m3_cyc_r_reg  ( .D(m3s7_cyc), .CLK(clock), .Q(\s7/m3_cyc_r ) );
  DFFX1 \s7/m2_cyc_r_reg  ( .D(m2s7_cyc), .CLK(clock), .Q(\s7/m2_cyc_r ) );
  DFFX1 \s7/m1_cyc_r_reg  ( .D(m1s7_cyc), .CLK(clock), .Q(\s7/m1_cyc_r ) );
  DFFX1 \s7/m0_cyc_r_reg  ( .D(m0s7_cyc), .CLK(clock), .Q(\s7/m0_cyc_r ) );
  DFFX1 \s7/next_reg  ( .D(n18186), .CLK(clock), .Q(\s7/next ), .QN(n34377) );
  DFFX1 \s8/m7_cyc_r_reg  ( .D(m7s8_cyc), .CLK(clock), .Q(\s8/m7_cyc_r ) );
  DFFX1 \s8/m6_cyc_r_reg  ( .D(m6s8_cyc), .CLK(clock), .Q(\s8/m6_cyc_r ) );
  DFFX1 \s8/m5_cyc_r_reg  ( .D(m5s8_cyc), .CLK(clock), .Q(\s8/m5_cyc_r ) );
  DFFX1 \s8/m4_cyc_r_reg  ( .D(m4s8_cyc), .CLK(clock), .Q(\s8/m4_cyc_r ) );
  DFFX1 \s8/m3_cyc_r_reg  ( .D(m3s8_cyc), .CLK(clock), .Q(\s8/m3_cyc_r ) );
  DFFX1 \s8/m2_cyc_r_reg  ( .D(m2s8_cyc), .CLK(clock), .Q(\s8/m2_cyc_r ) );
  DFFX1 \s8/m1_cyc_r_reg  ( .D(m1s8_cyc), .CLK(clock), .Q(\s8/m1_cyc_r ) );
  DFFX1 \s8/m0_cyc_r_reg  ( .D(m0s8_cyc), .CLK(clock), .Q(\s8/m0_cyc_r ) );
  DFFX1 \s8/next_reg  ( .D(n18185), .CLK(clock), .Q(\s8/next ), .QN(n34674) );
  DFFX1 \s9/m7_cyc_r_reg  ( .D(m7s9_cyc), .CLK(clock), .Q(\s9/m7_cyc_r ) );
  DFFX1 \s9/m6_cyc_r_reg  ( .D(m6s9_cyc), .CLK(clock), .Q(\s9/m6_cyc_r ) );
  DFFX1 \s9/m5_cyc_r_reg  ( .D(m5s9_cyc), .CLK(clock), .Q(\s9/m5_cyc_r ) );
  DFFX1 \s9/m4_cyc_r_reg  ( .D(m4s9_cyc), .CLK(clock), .Q(\s9/m4_cyc_r ) );
  DFFX1 \s9/m3_cyc_r_reg  ( .D(m3s9_cyc), .CLK(clock), .Q(\s9/m3_cyc_r ) );
  DFFX1 \s9/m2_cyc_r_reg  ( .D(m2s9_cyc), .CLK(clock), .Q(\s9/m2_cyc_r ) );
  DFFX1 \s9/m1_cyc_r_reg  ( .D(m1s9_cyc), .CLK(clock), .Q(\s9/m1_cyc_r ) );
  DFFX1 \s9/m0_cyc_r_reg  ( .D(m0s9_cyc), .CLK(clock), .Q(\s9/m0_cyc_r ) );
  DFFX1 \s9/next_reg  ( .D(n18184), .CLK(clock), .Q(\s9/next ) );
  DFFX1 \s10/m7_cyc_r_reg  ( .D(m7s10_cyc), .CLK(clock), .Q(\s10/m7_cyc_r ) );
  DFFX1 \s10/m6_cyc_r_reg  ( .D(m6s10_cyc), .CLK(clock), .Q(\s10/m6_cyc_r ) );
  DFFX1 \s10/m5_cyc_r_reg  ( .D(m5s10_cyc), .CLK(clock), .Q(\s10/m5_cyc_r ) );
  DFFX1 \s10/m4_cyc_r_reg  ( .D(m4s10_cyc), .CLK(clock), .Q(\s10/m4_cyc_r ) );
  DFFX1 \s10/m3_cyc_r_reg  ( .D(m3s10_cyc), .CLK(clock), .Q(\s10/m3_cyc_r ) );
  DFFX1 \s10/m2_cyc_r_reg  ( .D(m2s10_cyc), .CLK(clock), .Q(\s10/m2_cyc_r ) );
  DFFX1 \s10/m1_cyc_r_reg  ( .D(m1s10_cyc), .CLK(clock), .Q(\s10/m1_cyc_r ) );
  DFFX1 \s10/m0_cyc_r_reg  ( .D(m0s10_cyc), .CLK(clock), .Q(\s10/m0_cyc_r ) );
  DFFX1 \s10/next_reg  ( .D(n18183), .CLK(clock), .Q(\s10/next ), .QN(n34376)
         );
  DFFX1 \s11/m7_cyc_r_reg  ( .D(m7s11_cyc), .CLK(clock), .Q(\s11/m7_cyc_r ) );
  DFFX1 \s11/m6_cyc_r_reg  ( .D(m6s11_cyc), .CLK(clock), .Q(\s11/m6_cyc_r ) );
  DFFX1 \s11/m5_cyc_r_reg  ( .D(m5s11_cyc), .CLK(clock), .Q(\s11/m5_cyc_r ) );
  DFFX1 \s11/m4_cyc_r_reg  ( .D(m4s11_cyc), .CLK(clock), .Q(\s11/m4_cyc_r ) );
  DFFX1 \s11/m3_cyc_r_reg  ( .D(m3s11_cyc), .CLK(clock), .Q(\s11/m3_cyc_r ) );
  DFFX1 \s11/m2_cyc_r_reg  ( .D(m2s11_cyc), .CLK(clock), .Q(\s11/m2_cyc_r ) );
  DFFX1 \s11/m1_cyc_r_reg  ( .D(m1s11_cyc), .CLK(clock), .Q(\s11/m1_cyc_r ) );
  DFFX1 \s11/m0_cyc_r_reg  ( .D(m0s11_cyc), .CLK(clock), .Q(\s11/m0_cyc_r ) );
  DFFX1 \s11/next_reg  ( .D(n18182), .CLK(clock), .Q(\s11/next ) );
  DFFX1 \s12/m7_cyc_r_reg  ( .D(m7s12_cyc), .CLK(clock), .Q(\s12/m7_cyc_r ) );
  DFFX1 \s12/m6_cyc_r_reg  ( .D(m6s12_cyc), .CLK(clock), .Q(\s12/m6_cyc_r ) );
  DFFX1 \s12/m5_cyc_r_reg  ( .D(m5s12_cyc), .CLK(clock), .Q(\s12/m5_cyc_r ) );
  DFFX1 \s12/m4_cyc_r_reg  ( .D(m4s12_cyc), .CLK(clock), .Q(\s12/m4_cyc_r ) );
  DFFX1 \s12/m3_cyc_r_reg  ( .D(m3s12_cyc), .CLK(clock), .Q(\s12/m3_cyc_r ) );
  DFFX1 \s12/m2_cyc_r_reg  ( .D(m2s12_cyc), .CLK(clock), .Q(\s12/m2_cyc_r ) );
  DFFX1 \s12/m1_cyc_r_reg  ( .D(m1s12_cyc), .CLK(clock), .Q(\s12/m1_cyc_r ) );
  DFFX1 \s12/m0_cyc_r_reg  ( .D(m0s12_cyc), .CLK(clock), .Q(\s12/m0_cyc_r ) );
  DFFX1 \s12/next_reg  ( .D(n18181), .CLK(clock), .Q(\s12/next ) );
  DFFX1 \s13/m7_cyc_r_reg  ( .D(m7s13_cyc), .CLK(clock), .Q(\s13/m7_cyc_r ) );
  DFFX1 \s13/m6_cyc_r_reg  ( .D(m6s13_cyc), .CLK(clock), .Q(\s13/m6_cyc_r ) );
  DFFX1 \s13/m5_cyc_r_reg  ( .D(m5s13_cyc), .CLK(clock), .Q(\s13/m5_cyc_r ) );
  DFFX1 \s13/m4_cyc_r_reg  ( .D(m4s13_cyc), .CLK(clock), .Q(\s13/m4_cyc_r ) );
  DFFX1 \s13/m3_cyc_r_reg  ( .D(m3s13_cyc), .CLK(clock), .Q(\s13/m3_cyc_r ) );
  DFFX1 \s13/m2_cyc_r_reg  ( .D(m2s13_cyc), .CLK(clock), .Q(\s13/m2_cyc_r ) );
  DFFX1 \s13/m1_cyc_r_reg  ( .D(m1s13_cyc), .CLK(clock), .Q(\s13/m1_cyc_r ) );
  DFFX1 \s13/m0_cyc_r_reg  ( .D(m0s13_cyc), .CLK(clock), .Q(\s13/m0_cyc_r ) );
  DFFX1 \s13/next_reg  ( .D(n18180), .CLK(clock), .Q(\s13/next ) );
  DFFX1 \s14/m7_cyc_r_reg  ( .D(m7s14_cyc), .CLK(clock), .Q(\s14/m7_cyc_r ) );
  DFFX1 \s14/m6_cyc_r_reg  ( .D(m6s14_cyc), .CLK(clock), .Q(\s14/m6_cyc_r ) );
  DFFX1 \s14/m5_cyc_r_reg  ( .D(m5s14_cyc), .CLK(clock), .Q(\s14/m5_cyc_r ) );
  DFFX1 \s14/m4_cyc_r_reg  ( .D(m4s14_cyc), .CLK(clock), .Q(\s14/m4_cyc_r ) );
  DFFX1 \s14/m3_cyc_r_reg  ( .D(m3s14_cyc), .CLK(clock), .Q(\s14/m3_cyc_r ) );
  DFFX1 \s14/m2_cyc_r_reg  ( .D(m2s14_cyc), .CLK(clock), .Q(\s14/m2_cyc_r ) );
  DFFX1 \s14/m1_cyc_r_reg  ( .D(m1s14_cyc), .CLK(clock), .Q(\s14/m1_cyc_r ) );
  DFFX1 \s14/m0_cyc_r_reg  ( .D(m0s14_cyc), .CLK(clock), .Q(\s14/m0_cyc_r ) );
  DFFX1 \s14/next_reg  ( .D(n18179), .CLK(clock), .Q(\s14/next ) );
  DFFX1 \s15/m7_cyc_r_reg  ( .D(m7s15_cyc), .CLK(clock), .Q(\s15/m7_cyc_r ) );
  DFFX1 \s15/m6_cyc_r_reg  ( .D(m6s15_cyc), .CLK(clock), .Q(\s15/m6_cyc_r ) );
  DFFX1 \s15/m5_cyc_r_reg  ( .D(m5s15_cyc), .CLK(clock), .Q(\s15/m5_cyc_r ) );
  DFFX1 \s15/m4_cyc_r_reg  ( .D(m4s15_cyc), .CLK(clock), .Q(\s15/m4_cyc_r ) );
  DFFX1 \s15/m3_cyc_r_reg  ( .D(m3s15_cyc), .CLK(clock), .Q(\s15/m3_cyc_r ) );
  DFFX1 \s15/m2_cyc_r_reg  ( .D(m2s15_cyc), .CLK(clock), .Q(\s15/m2_cyc_r ) );
  DFFX1 \s15/m1_cyc_r_reg  ( .D(m1s15_cyc), .CLK(clock), .Q(\s15/m1_cyc_r ) );
  DFFX1 \s15/m0_cyc_r_reg  ( .D(m0s15_cyc), .CLK(clock), .Q(\s15/m0_cyc_r ) );
  DFFX1 \s15/next_reg  ( .D(n18178), .CLK(clock), .Q(\s15/next ) );
  DFFX1 \rf/rf_dout_reg[0]  ( .D(\rf/N115 ), .CLK(clock), .Q(\rf/rf_dout [0])
         );
  DFFX1 \rf/rf_dout_reg[1]  ( .D(\rf/N116 ), .CLK(clock), .Q(\rf/rf_dout [1])
         );
  DFFX1 \rf/rf_dout_reg[2]  ( .D(\rf/N117 ), .CLK(clock), .Q(\rf/rf_dout [2])
         );
  DFFX1 \rf/rf_dout_reg[3]  ( .D(\rf/N118 ), .CLK(clock), .Q(\rf/rf_dout [3])
         );
  DFFX1 \rf/rf_dout_reg[4]  ( .D(\rf/N119 ), .CLK(clock), .Q(\rf/rf_dout [4])
         );
  DFFX1 \rf/rf_dout_reg[5]  ( .D(\rf/N120 ), .CLK(clock), .Q(\rf/rf_dout [5])
         );
  DFFX1 \rf/rf_dout_reg[6]  ( .D(\rf/N121 ), .CLK(clock), .Q(\rf/rf_dout [6])
         );
  DFFX1 \rf/rf_dout_reg[7]  ( .D(\rf/N122 ), .CLK(clock), .Q(\rf/rf_dout [7])
         );
  DFFX1 \rf/rf_dout_reg[8]  ( .D(\rf/N123 ), .CLK(clock), .Q(\rf/rf_dout [8])
         );
  DFFX1 \rf/rf_dout_reg[9]  ( .D(\rf/N124 ), .CLK(clock), .Q(\rf/rf_dout [9])
         );
  DFFX1 \rf/rf_dout_reg[10]  ( .D(\rf/N125 ), .CLK(clock), .Q(\rf/rf_dout [10]) );
  DFFX1 \rf/rf_dout_reg[11]  ( .D(\rf/N126 ), .CLK(clock), .Q(\rf/rf_dout [11]) );
  DFFX1 \rf/rf_dout_reg[12]  ( .D(\rf/N127 ), .CLK(clock), .Q(\rf/rf_dout [12]) );
  DFFX1 \rf/rf_dout_reg[13]  ( .D(\rf/N128 ), .CLK(clock), .Q(\rf/rf_dout [13]) );
  DFFX1 \rf/rf_dout_reg[14]  ( .D(\rf/N129 ), .CLK(clock), .Q(\rf/rf_dout [14]) );
  DFFX1 \rf/rf_dout_reg[15]  ( .D(\rf/N130 ), .CLK(clock), .Q(\rf/rf_dout [15]) );
  DFFX1 \rf/rf_ack_reg  ( .D(\rf/N19 ), .CLK(clock), .Q(\rf/rf_ack ) );
  DFFX1 \rf/rf_we_reg  ( .D(\rf/N18 ), .CLK(clock), .QN(n34379) );
  DFFX1 \s0/msel/pri_out_reg[0]  ( .D(n17599), .CLK(clock), .Q(
        \s0/msel/pri_out [0]) );
  DFFX1 \s0/msel/pri_out_reg[1]  ( .D(n17598), .CLK(clock), .Q(
        \s0/msel/pri_out [1]) );
  DFFX1 \s1/msel/pri_out_reg[0]  ( .D(n17597), .CLK(clock), .Q(
        \s1/msel/pri_out [0]) );
  DFFX1 \s1/msel/pri_out_reg[1]  ( .D(n17596), .CLK(clock), .Q(
        \s1/msel/pri_out [1]) );
  DFFX1 \s2/msel/pri_out_reg[0]  ( .D(n17595), .CLK(clock), .Q(
        \s2/msel/pri_out [0]) );
  DFFX1 \s2/msel/pri_out_reg[1]  ( .D(n17594), .CLK(clock), .Q(
        \s2/msel/pri_out [1]) );
  DFFX1 \s3/msel/pri_out_reg[0]  ( .D(n17593), .CLK(clock), .Q(
        \s3/msel/pri_out [0]) );
  DFFX1 \s3/msel/pri_out_reg[1]  ( .D(n17592), .CLK(clock), .Q(
        \s3/msel/pri_out [1]) );
  DFFX1 \s4/msel/pri_out_reg[0]  ( .D(n17591), .CLK(clock), .Q(
        \s4/msel/pri_out [0]) );
  DFFX1 \s4/msel/pri_out_reg[1]  ( .D(n17590), .CLK(clock), .Q(
        \s4/msel/pri_out [1]) );
  DFFX1 \s5/msel/pri_out_reg[0]  ( .D(n17589), .CLK(clock), .Q(
        \s5/msel/pri_out [0]) );
  DFFX1 \s5/msel/pri_out_reg[1]  ( .D(n17588), .CLK(clock), .Q(
        \s5/msel/pri_out [1]) );
  DFFX1 \s6/msel/pri_out_reg[0]  ( .D(n17587), .CLK(clock), .Q(
        \s6/msel/pri_out [0]) );
  DFFX1 \s6/msel/pri_out_reg[1]  ( .D(n17586), .CLK(clock), .Q(
        \s6/msel/pri_out [1]) );
  DFFX1 \s7/msel/pri_out_reg[0]  ( .D(n17585), .CLK(clock), .Q(
        \s7/msel/pri_out [0]), .QN(n34676) );
  DFFX1 \s7/msel/pri_out_reg[1]  ( .D(n17584), .CLK(clock), .Q(
        \s7/msel/pri_out [1]) );
  DFFX1 \s8/msel/pri_out_reg[0]  ( .D(n17583), .CLK(clock), .Q(
        \s8/msel/pri_out [0]) );
  DFFX1 \s8/msel/pri_out_reg[1]  ( .D(n17582), .CLK(clock), .Q(
        \s8/msel/pri_out [1]) );
  DFFX1 \s9/msel/pri_out_reg[0]  ( .D(n17581), .CLK(clock), .Q(
        \s9/msel/pri_out [0]) );
  DFFX1 \s9/msel/pri_out_reg[1]  ( .D(n17580), .CLK(clock), .Q(
        \s9/msel/pri_out [1]) );
  DFFX1 \s10/msel/pri_out_reg[0]  ( .D(n17579), .CLK(clock), .Q(
        \s10/msel/pri_out [0]) );
  DFFX1 \s10/msel/pri_out_reg[1]  ( .D(n17578), .CLK(clock), .Q(
        \s10/msel/pri_out [1]), .QN(n34672) );
  DFFX1 \s11/msel/pri_out_reg[0]  ( .D(n17577), .CLK(clock), .Q(
        \s11/msel/pri_out [0]) );
  DFFX1 \s11/msel/pri_out_reg[1]  ( .D(n17576), .CLK(clock), .Q(
        \s11/msel/pri_out [1]) );
  DFFX1 \s12/msel/pri_out_reg[0]  ( .D(n17575), .CLK(clock), .Q(
        \s12/msel/pri_out [0]) );
  DFFX1 \s12/msel/pri_out_reg[1]  ( .D(n17574), .CLK(clock), .Q(
        \s12/msel/pri_out [1]) );
  DFFX1 \s13/msel/pri_out_reg[0]  ( .D(n17573), .CLK(clock), .Q(
        \s13/msel/pri_out [0]) );
  DFFX1 \s13/msel/pri_out_reg[1]  ( .D(n17572), .CLK(clock), .Q(
        \s13/msel/pri_out [1]) );
  DFFX1 \s14/msel/pri_out_reg[0]  ( .D(n17571), .CLK(clock), .Q(
        \s14/msel/pri_out [0]) );
  DFFX1 \s14/msel/pri_out_reg[1]  ( .D(n17570), .CLK(clock), .Q(
        \s14/msel/pri_out [1]) );
  DFFX1 \s15/msel/pri_out_reg[0]  ( .D(n17569), .CLK(clock), .Q(
        \s15/msel/pri_out [0]) );
  DFFX1 \s15/msel/pri_out_reg[1]  ( .D(n17568), .CLK(clock), .Q(
        \s15/msel/pri_out [1]) );
  DFFARX1 \rf/conf15_reg[15]  ( .D(n17614), .CLK(clock), .RSTB(n34689), .Q(
        n34518), .QN(n13485) );
  DFFARX1 \rf/conf15_reg[14]  ( .D(n17615), .CLK(clock), .RSTB(n34695), .Q(
        n34301), .QN(n13538) );
  DFFARX1 \rf/conf15_reg[13]  ( .D(n17616), .CLK(clock), .RSTB(n34688), .Q(
        n34598), .QN(n13564) );
  DFFARX1 \rf/conf15_reg[0]  ( .D(n17629), .CLK(clock), .RSTB(n34685), .Q(
        n34298), .QN(n13914) );
  DFFARX1 \rf/conf15_reg[1]  ( .D(n17628), .CLK(clock), .RSTB(n34687), .Q(
        n34482), .QN(n13876) );
  DFFARX1 \rf/conf15_reg[2]  ( .D(n17627), .CLK(clock), .RSTB(n34694), .Q(
        n34302), .QN(n13850) );
  DFFARX1 \rf/conf15_reg[3]  ( .D(n17626), .CLK(clock), .RSTB(n34691), .Q(
        n34514), .QN(n13824) );
  DFFARX1 \rf/conf15_reg[4]  ( .D(n17625), .CLK(clock), .RSTB(n34693), .Q(
        n34359), .QN(n13798) );
  DFFARX1 \rf/conf15_reg[5]  ( .D(n17624), .CLK(clock), .RSTB(n34684), .Q(
        n34602), .QN(n13772) );
  DFFARX1 \rf/conf15_reg[6]  ( .D(n17623), .CLK(clock), .RSTB(n34694), .Q(
        n34303), .QN(n13746) );
  DFFARX1 \rf/conf15_reg[7]  ( .D(n17622), .CLK(clock), .RSTB(n34682), .Q(
        n34515), .QN(n13720) );
  DFFARX1 \rf/conf15_reg[8]  ( .D(n17621), .CLK(clock), .RSTB(n34680), .Q(
        n34299), .QN(n13694) );
  DFFARX1 \rf/conf15_reg[9]  ( .D(n17620), .CLK(clock), .RSTB(n34691), .Q(
        n34516), .QN(n13668) );
  DFFARX1 \rf/conf15_reg[10]  ( .D(n17619), .CLK(clock), .RSTB(n34689), .Q(
        n34300), .QN(n13642) );
  DFFARX1 \rf/conf15_reg[11]  ( .D(n17618), .CLK(clock), .RSTB(n34681), .Q(
        n34517), .QN(n13616) );
  DFFARX1 \rf/conf15_reg[12]  ( .D(n17617), .CLK(clock), .RSTB(n34693), .Q(
        n34360), .QN(n13590) );
  DFFARX1 \rf/conf14_reg[0]  ( .D(n17657), .CLK(clock), .RSTB(n34697), .Q(
        n34367), .QN(n13912) );
  DFFARX1 \rf/conf14_reg[1]  ( .D(n17656), .CLK(clock), .RSTB(n34696), .Q(
        n34604), .QN(n13875) );
  DFFARX1 \rf/conf14_reg[2]  ( .D(n17655), .CLK(clock), .RSTB(n34695), .Q(
        n34334), .QN(n13849) );
  DFFARX1 \rf/conf14_reg[3]  ( .D(n17654), .CLK(clock), .RSTB(n34679), .Q(
        n34512), .QN(n13823) );
  DFFARX1 \rf/conf14_reg[4]  ( .D(n17653), .CLK(clock), .RSTB(n34694), .Q(
        n34477), .QN(n13797) );
  DFFARX1 \rf/conf14_reg[5]  ( .D(n17652), .CLK(clock), .RSTB(n34688), .Q(
        n34646), .QN(n13771) );
  DFFARX1 \rf/conf14_reg[6]  ( .D(n17651), .CLK(clock), .RSTB(n34692), .Q(
        n34481), .QN(n13745) );
  DFFARX1 \rf/conf14_reg[7]  ( .D(n17650), .CLK(clock), .RSTB(n34692), .Q(
        n34648), .QN(n13719) );
  DFFARX1 \rf/conf14_reg[8]  ( .D(n17649), .CLK(clock), .RSTB(n34692), .Q(
        n34635), .QN(n13693) );
  DFFARX1 \rf/conf14_reg[9]  ( .D(n17648), .CLK(clock), .RSTB(n34692), .Q(
        n34571), .QN(n13667) );
  DFFARX1 \rf/conf14_reg[10]  ( .D(n17647), .CLK(clock), .RSTB(n34692), .Q(
        n34547), .QN(n13641) );
  DFFARX1 \rf/conf14_reg[11]  ( .D(n17646), .CLK(clock), .RSTB(n34692), .Q(
        n34652), .QN(n13615) );
  DFFARX1 \rf/conf14_reg[12]  ( .D(n17645), .CLK(clock), .RSTB(n34692), .Q(
        n34357), .QN(n13589) );
  DFFARX1 \rf/conf14_reg[13]  ( .D(n17644), .CLK(clock), .RSTB(n34692), .Q(
        n34544), .QN(n13563) );
  DFFARX1 \rf/conf14_reg[14]  ( .D(n17643), .CLK(clock), .RSTB(n34692), .Q(
        n34358), .QN(n13537) );
  DFFARX1 \rf/conf14_reg[15]  ( .D(n17642), .CLK(clock), .RSTB(n34692), .Q(
        n34513), .QN(n13484) );
  DFFARX1 \rf/conf13_reg[0]  ( .D(n17685), .CLK(clock), .RSTB(n34692), .Q(
        n34356), .QN(n13910) );
  DFFARX1 \rf/conf13_reg[1]  ( .D(n17684), .CLK(clock), .RSTB(n34692), .Q(
        n34542), .QN(n13874) );
  DFFARX1 \rf/conf13_reg[2]  ( .D(n17683), .CLK(clock), .RSTB(n34692), .Q(
        n34332), .QN(n13848) );
  DFFARX1 \rf/conf13_reg[3]  ( .D(n17682), .CLK(clock), .RSTB(n34677), .Q(
        n34510), .QN(n13822) );
  DFFARX1 \rf/conf13_reg[4]  ( .D(n17681), .CLK(clock), .RSTB(n34678), .Q(
        n34480), .QN(n13796) );
  DFFARX1 \rf/conf13_reg[5]  ( .D(n17680), .CLK(clock), .RSTB(n34685), .Q(
        n34645), .QN(n13770) );
  DFFARX1 \rf/conf13_reg[6]  ( .D(n17679), .CLK(clock), .RSTB(n34684), .Q(
        n34546), .QN(n13744) );
  DFFARX1 \rf/conf13_reg[7]  ( .D(n17678), .CLK(clock), .RSTB(n34682), .Q(
        n34651), .QN(n13718) );
  DFFARX1 \rf/conf13_reg[8]  ( .D(n17677), .CLK(clock), .RSTB(n34680), .Q(
        n34333), .QN(n13692) );
  DFFARX1 \rf/conf13_reg[9]  ( .D(n17676), .CLK(clock), .RSTB(n34691), .Q(
        n34543), .QN(n13666) );
  DFFARX1 \rf/conf13_reg[10]  ( .D(n17675), .CLK(clock), .RSTB(n34689), .Q(
        n34476), .QN(n13640) );
  DFFARX1 \rf/conf13_reg[11]  ( .D(n17674), .CLK(clock), .RSTB(n34681), .Q(
        n34644), .QN(n13614) );
  DFFARX1 \rf/conf13_reg[12]  ( .D(n17673), .CLK(clock), .RSTB(n34693), .Q(
        n34331), .QN(n13588) );
  DFFARX1 \rf/conf13_reg[13]  ( .D(n17672), .CLK(clock), .RSTB(n34697), .Q(
        n34511), .QN(n13562) );
  DFFARX1 \rf/conf13_reg[14]  ( .D(n17671), .CLK(clock), .RSTB(n34677), .Q(
        n34634), .QN(n13536) );
  DFFARX1 \rf/conf13_reg[15]  ( .D(n17670), .CLK(clock), .RSTB(n34693), .Q(
        n34586), .QN(n13482) );
  DFFARX1 \rf/conf12_reg[0]  ( .D(n17713), .CLK(clock), .RSTB(n34684), .Q(
        n34354), .QN(n13908) );
  DFFARX1 \rf/conf12_reg[1]  ( .D(n17712), .CLK(clock), .RSTB(n34688), .Q(
        n34509), .QN(n13873) );
  DFFARX1 \rf/conf12_reg[2]  ( .D(n17711), .CLK(clock), .RSTB(n34681), .Q(
        n34355), .QN(n13847) );
  DFFARX1 \rf/conf12_reg[3]  ( .D(n17710), .CLK(clock), .RSTB(n34682), .Q(
        n34508), .QN(n13821) );
  DFFARX1 \rf/conf12_reg[4]  ( .D(n17709), .CLK(clock), .RSTB(n34697), .Q(
        n34329), .QN(n13795) );
  DFFARX1 \rf/conf12_reg[5]  ( .D(n17708), .CLK(clock), .RSTB(n34677), .Q(
        n34541), .QN(n13769) );
  DFFARX1 \rf/conf12_reg[6]  ( .D(n17707), .CLK(clock), .RSTB(n34696), .Q(
        n34330), .QN(n13743) );
  DFFARX1 \rf/conf12_reg[7]  ( .D(n17706), .CLK(clock), .RSTB(n34695), .Q(
        n34507), .QN(n13717) );
  DFFARX1 \rf/conf12_reg[8]  ( .D(n17705), .CLK(clock), .RSTB(n34679), .Q(
        n34475), .QN(n13691) );
  DFFARX1 \rf/conf12_reg[9]  ( .D(n17704), .CLK(clock), .RSTB(n34693), .Q(
        n34642), .QN(n13665) );
  DFFARX1 \rf/conf12_reg[10]  ( .D(n17703), .CLK(clock), .RSTB(n34693), .Q(
        n34328), .QN(n13639) );
  DFFARX1 \rf/conf12_reg[11]  ( .D(n17702), .CLK(clock), .RSTB(n34693), .Q(
        n34506), .QN(n13613) );
  DFFARX1 \rf/conf12_reg[12]  ( .D(n17701), .CLK(clock), .RSTB(n34693), .Q(
        n34327), .QN(n13587) );
  DFFARX1 \rf/conf12_reg[13]  ( .D(n17700), .CLK(clock), .RSTB(n34693), .Q(
        n34540), .QN(n13561) );
  DFFARX1 \rf/conf12_reg[14]  ( .D(n17699), .CLK(clock), .RSTB(n34693), .Q(
        n34474), .QN(n13535) );
  DFFARX1 \rf/conf12_reg[15]  ( .D(n17698), .CLK(clock), .RSTB(n34693), .Q(
        n34643), .QN(n13481) );
  DFFARX1 \rf/conf11_reg[0]  ( .D(n17741), .CLK(clock), .RSTB(n34693), .Q(
        n34621), .QN(n13922) );
  DFFARX1 \rf/conf11_reg[1]  ( .D(n17740), .CLK(clock), .RSTB(n34693), .Q(
        n34584), .QN(n13880) );
  DFFARX1 \rf/conf11_reg[2]  ( .D(n17739), .CLK(clock), .RSTB(n34693), .Q(
        n34326), .QN(n13854) );
  DFFARX1 \rf/conf11_reg[3]  ( .D(n17738), .CLK(clock), .RSTB(n34693), .Q(
        n34537), .QN(n13828) );
  DFFARX1 \rf/conf11_reg[4]  ( .D(n17737), .CLK(clock), .RSTB(n34693), .Q(
        n34325), .QN(n13802) );
  DFFARX1 \rf/conf11_reg[5]  ( .D(n17736), .CLK(clock), .RSTB(n34694), .Q(
        n34538), .QN(n13776) );
  DFFARX1 \rf/conf11_reg[6]  ( .D(n17735), .CLK(clock), .RSTB(n34694), .Q(
        n34365), .QN(n13750) );
  DFFARX1 \rf/conf11_reg[7]  ( .D(n17734), .CLK(clock), .RSTB(n34694), .Q(
        n34601), .QN(n13724) );
  DFFARX1 \rf/conf11_reg[8]  ( .D(n17733), .CLK(clock), .RSTB(n34694), .Q(
        n34622), .QN(n13698) );
  DFFARX1 \rf/conf11_reg[9]  ( .D(n17732), .CLK(clock), .RSTB(n34694), .Q(
        n34569), .QN(n13672) );
  DFFARX1 \rf/conf11_reg[10]  ( .D(n17731), .CLK(clock), .RSTB(n34694), .Q(
        n34375), .QN(n13646) );
  DFFARX1 \rf/conf11_reg[11]  ( .D(n17730), .CLK(clock), .RSTB(n34694), .Q(
        n34585), .QN(n13620) );
  DFFARX1 \rf/conf11_reg[12]  ( .D(n17729), .CLK(clock), .RSTB(n34694), .Q(
        n34633), .QN(n13594) );
  DFFARX1 \rf/conf11_reg[13]  ( .D(n17728), .CLK(clock), .RSTB(n34694), .Q(
        n34570), .QN(n13568) );
  DFFARX1 \rf/conf11_reg[14]  ( .D(n17727), .CLK(clock), .RSTB(n34694), .Q(
        n34324), .QN(n13542) );
  DFFARX1 \rf/conf11_reg[15]  ( .D(n17726), .CLK(clock), .RSTB(n34694), .Q(
        n34539), .QN(n13495) );
  DFFARX1 \rf/conf10_reg[0]  ( .D(n17769), .CLK(clock), .RSTB(n34694), .Q(
        n34619), .QN(n13920) );
  DFFARX1 \rf/conf10_reg[1]  ( .D(n17768), .CLK(clock), .RSTB(n34695), .Q(
        n34582), .QN(n13879) );
  DFFARX1 \rf/conf10_reg[2]  ( .D(n17767), .CLK(clock), .RSTB(n34695), .Q(
        n34638), .QN(n13853) );
  DFFARX1 \rf/conf10_reg[3]  ( .D(n17766), .CLK(clock), .RSTB(n34695), .Q(
        n34611), .QN(n13827) );
  DFFARX1 \rf/conf10_reg[4]  ( .D(n17765), .CLK(clock), .RSTB(n34695), .Q(
        n34322), .QN(n13801) );
  DFFARX1 \rf/conf10_reg[5]  ( .D(n17764), .CLK(clock), .RSTB(n34695), .Q(
        n34503), .QN(n13775) );
  DFFARX1 \rf/conf10_reg[6]  ( .D(n17763), .CLK(clock), .RSTB(n34695), .Q(
        n34606), .QN(n13749) );
  DFFARX1 \rf/conf10_reg[7]  ( .D(n17762), .CLK(clock), .RSTB(n34695), .Q(
        n34372), .QN(n13723) );
  DFFARX1 \rf/conf10_reg[8]  ( .D(n17761), .CLK(clock), .RSTB(n34695), .Q(
        n34620), .QN(n13697) );
  DFFARX1 \rf/conf10_reg[9]  ( .D(n17760), .CLK(clock), .RSTB(n34695), .Q(
        n34583), .QN(n13671) );
  DFFARX1 \rf/conf10_reg[10]  ( .D(n17759), .CLK(clock), .RSTB(n34695), .Q(
        n34323), .QN(n13645) );
  DFFARX1 \rf/conf10_reg[11]  ( .D(n17758), .CLK(clock), .RSTB(n34695), .Q(
        n34504), .QN(n13619) );
  DFFARX1 \rf/conf10_reg[12]  ( .D(n17757), .CLK(clock), .RSTB(n34695), .Q(
        n34632), .QN(n13593) );
  DFFARX1 \rf/conf10_reg[13]  ( .D(n17756), .CLK(clock), .RSTB(n34696), .Q(
        n34568), .QN(n13567) );
  DFFARX1 \rf/conf10_reg[14]  ( .D(n17755), .CLK(clock), .RSTB(n34696), .Q(
        n34353), .QN(n13541) );
  DFFARX1 \rf/conf10_reg[15]  ( .D(n17754), .CLK(clock), .RSTB(n34696), .Q(
        n34505), .QN(n13494) );
  DFFARX1 \rf/conf9_reg[0]  ( .D(n17797), .CLK(clock), .RSTB(n34696), .Q(
        n34321), .QN(n13918) );
  DFFARX1 \rf/conf9_reg[1]  ( .D(n17796), .CLK(clock), .RSTB(n34696), .Q(
        n34502), .QN(n13878) );
  DFFARX1 \rf/conf9_reg[2]  ( .D(n17795), .CLK(clock), .RSTB(n34696), .Q(
        n34618), .QN(n13852) );
  DFFARX1 \rf/conf9_reg[3]  ( .D(n17794), .CLK(clock), .RSTB(n34696), .Q(
        n34581), .QN(n13826) );
  DFFARX1 \rf/conf9_reg[4]  ( .D(n17793), .CLK(clock), .RSTB(n34696), .Q(
        n34352), .QN(n13800) );
  DFFARX1 \rf/conf9_reg[5]  ( .D(n17792), .CLK(clock), .RSTB(n34696), .Q(
        n34535), .QN(n13774) );
  DFFARX1 \rf/conf9_reg[6]  ( .D(n17791), .CLK(clock), .RSTB(n34696), .Q(
        n34636), .QN(n13748) );
  DFFARX1 \rf/conf9_reg[7]  ( .D(n17790), .CLK(clock), .RSTB(n34696), .Q(
        n34596), .QN(n13722) );
  DFFARX1 \rf/conf9_reg[8]  ( .D(n17789), .CLK(clock), .RSTB(n34696), .Q(
        n34319), .QN(n13696) );
  DFFARX1 \rf/conf9_reg[9]  ( .D(n17788), .CLK(clock), .RSTB(n34697), .Q(
        n34536), .QN(n13670) );
  DFFARX1 \rf/conf9_reg[10]  ( .D(n17787), .CLK(clock), .RSTB(n34697), .Q(
        n34351), .QN(n13644) );
  DFFARX1 \rf/conf9_reg[11]  ( .D(n17786), .CLK(clock), .RSTB(n34697), .Q(
        n34501), .QN(n13618) );
  DFFARX1 \rf/conf9_reg[12]  ( .D(n17785), .CLK(clock), .RSTB(n34697), .Q(
        n34320), .QN(n13592) );
  DFFARX1 \rf/conf9_reg[13]  ( .D(n17784), .CLK(clock), .RSTB(n34697), .Q(
        n34500), .QN(n13566) );
  DFFARX1 \rf/conf9_reg[14]  ( .D(n17783), .CLK(clock), .RSTB(n34697), .Q(
        n34364), .QN(n13540) );
  DFFARX1 \rf/conf9_reg[15]  ( .D(n17782), .CLK(clock), .RSTB(n34697), .Q(
        n34603), .QN(n13490) );
  DFFARX1 \rf/conf8_reg[0]  ( .D(n17825), .CLK(clock), .RSTB(n34697), .Q(
        n34659), .QN(n13916) );
  DFFARX1 \rf/conf8_reg[1]  ( .D(n17824), .CLK(clock), .RSTB(n34697), .Q(
        n34589), .QN(n13877) );
  DFFARX1 \rf/conf8_reg[2]  ( .D(n17823), .CLK(clock), .RSTB(n34697), .Q(
        n34660), .QN(n13851) );
  DFFARX1 \rf/conf8_reg[3]  ( .D(n17822), .CLK(clock), .RSTB(n34697), .Q(
        n34593), .QN(n13825) );
  DFFARX1 \rf/conf8_reg[4]  ( .D(n17821), .CLK(clock), .RSTB(n34697), .Q(
        n34662), .QN(n13799) );
  DFFARX1 \rf/conf8_reg[5]  ( .D(n17820), .CLK(clock), .RSTB(n34686), .Q(
        n34591), .QN(n13773) );
  DFFARX1 \rf/conf8_reg[6]  ( .D(n17819), .CLK(clock), .RSTB(n34680), .Q(
        n34663), .QN(n13747) );
  DFFARX1 \rf/conf8_reg[7]  ( .D(n17818), .CLK(clock), .RSTB(n34680), .Q(
        n34590), .QN(n13721) );
  DFFARX1 \rf/conf8_reg[8]  ( .D(n17817), .CLK(clock), .RSTB(n34680), .Q(
        n34238), .QN(n13695) );
  DFFARX1 \rf/conf8_reg[9]  ( .D(n17816), .CLK(clock), .RSTB(n34681), .Q(
        n34369), .QN(n13669) );
  DFFARX1 \rf/conf8_reg[10]  ( .D(n17815), .CLK(clock), .RSTB(n34681), .Q(
        n34588), .QN(n13643) );
  DFFARX1 \rf/conf8_reg[11]  ( .D(n17814), .CLK(clock), .RSTB(n34681), .Q(
        n34239), .QN(n13617) );
  DFFARX1 \rf/conf8_reg[12]  ( .D(n17813), .CLK(clock), .RSTB(n34681), .Q(
        n34631), .QN(n13591) );
  DFFARX1 \rf/conf8_reg[13]  ( .D(n17812), .CLK(clock), .RSTB(n34681), .Q(
        n34580), .QN(n13565) );
  DFFARX1 \rf/conf8_reg[14]  ( .D(n17811), .CLK(clock), .RSTB(n34681), .Q(
        n34661), .QN(n13539) );
  DFFARX1 \rf/conf8_reg[15]  ( .D(n17810), .CLK(clock), .RSTB(n34681), .Q(
        n34592), .QN(n13489) );
  DFFARX1 \rf/conf7_reg[0]  ( .D(n17853), .CLK(clock), .RSTB(n34681), .Q(
        n34349), .QN(n13894) );
  DFFARX1 \rf/conf7_reg[1]  ( .D(n17852), .CLK(clock), .RSTB(n34681), .Q(
        n34497), .QN(n13864) );
  DFFARX1 \rf/conf7_reg[2]  ( .D(n17851), .CLK(clock), .RSTB(n34681), .Q(
        n34348), .QN(n13838) );
  DFFARX1 \rf/conf7_reg[3]  ( .D(n17850), .CLK(clock), .RSTB(n34681), .Q(
        n34533), .QN(n13812) );
  DFFARX1 \rf/conf7_reg[4]  ( .D(n17849), .CLK(clock), .RSTB(n34681), .Q(
        n34363), .QN(n13786) );
  DFFARX1 \rf/conf7_reg[5]  ( .D(n17848), .CLK(clock), .RSTB(n34682), .Q(
        n34600), .QN(n13760) );
  DFFARX1 \rf/conf7_reg[6]  ( .D(n17847), .CLK(clock), .RSTB(n34682), .Q(
        n34318), .QN(n13734) );
  DFFARX1 \rf/conf7_reg[7]  ( .D(n17846), .CLK(clock), .RSTB(n34682), .Q(
        n34498), .QN(n13708) );
  DFFARX1 \rf/conf7_reg[8]  ( .D(n17845), .CLK(clock), .RSTB(n34682), .Q(
        n34649), .QN(n13682) );
  DFFARX1 \rf/conf7_reg[9]  ( .D(n17844), .CLK(clock), .RSTB(n34682), .Q(
        n34594), .QN(n13656) );
  DFFARX1 \rf/conf7_reg[10]  ( .D(n17843), .CLK(clock), .RSTB(n34682), .Q(
        n34350), .QN(n13630) );
  DFFARX1 \rf/conf7_reg[11]  ( .D(n17842), .CLK(clock), .RSTB(n34682), .Q(
        n34534), .QN(n13604) );
  DFFARX1 \rf/conf7_reg[12]  ( .D(n17841), .CLK(clock), .RSTB(n34682), .Q(
        n34374), .QN(n13578) );
  DFFARX1 \rf/conf7_reg[13]  ( .D(n17840), .CLK(clock), .RSTB(n34682), .Q(
        n34567), .QN(n13552) );
  DFFARX1 \rf/conf7_reg[14]  ( .D(n17839), .CLK(clock), .RSTB(n34682), .Q(
        n34347), .QN(n13526) );
  DFFARX1 \rf/conf7_reg[15]  ( .D(n17838), .CLK(clock), .RSTB(n34682), .Q(
        n34499), .QN(n13470) );
  DFFARX1 \rf/conf6_reg[0]  ( .D(n17881), .CLK(clock), .RSTB(n34682), .Q(
        n34629), .QN(n13892) );
  DFFARX1 \rf/conf6_reg[1]  ( .D(n17880), .CLK(clock), .RSTB(n34683), .Q(
        n34579), .QN(n13863) );
  DFFARX1 \rf/conf6_reg[2]  ( .D(n17879), .CLK(clock), .RSTB(n34683), .Q(
        n34237), .QN(n13837) );
  DFFARX1 \rf/conf6_reg[3]  ( .D(n17878), .CLK(clock), .RSTB(n34683), .Q(
        n34368), .QN(n13811) );
  DFFARX1 \rf/conf6_reg[4]  ( .D(n17877), .CLK(clock), .RSTB(n34683), .Q(
        n34362), .QN(n13785) );
  DFFARX1 \rf/conf6_reg[5]  ( .D(n17876), .CLK(clock), .RSTB(n34683), .Q(
        n34552), .QN(n13759) );
  DFFARX1 \rf/conf6_reg[6]  ( .D(n17875), .CLK(clock), .RSTB(n34683), .Q(
        n34346), .QN(n13733) );
  DFFARX1 \rf/conf6_reg[7]  ( .D(n17874), .CLK(clock), .RSTB(n34683), .Q(
        n34532), .QN(n13707) );
  DFFARX1 \rf/conf6_reg[8]  ( .D(n17873), .CLK(clock), .RSTB(n34683), .Q(
        n34630), .QN(n13681) );
  DFFARX1 \rf/conf6_reg[9]  ( .D(n17872), .CLK(clock), .RSTB(n34683), .Q(
        n34566), .QN(n13655) );
  DFFARX1 \rf/conf6_reg[10]  ( .D(n17871), .CLK(clock), .RSTB(n34683), .Q(
        n34345), .QN(n13629) );
  DFFARX1 \rf/conf6_reg[11]  ( .D(n17870), .CLK(clock), .RSTB(n34683), .Q(
        n34531), .QN(n13603) );
  DFFARX1 \rf/conf6_reg[12]  ( .D(n17869), .CLK(clock), .RSTB(n34683), .Q(
        n34366), .QN(n13577) );
  DFFARX1 \rf/conf6_reg[13]  ( .D(n17868), .CLK(clock), .RSTB(n34684), .Q(
        n34599), .QN(n13551) );
  DFFARX1 \rf/conf6_reg[14]  ( .D(n17867), .CLK(clock), .RSTB(n34684), .Q(
        n34628), .QN(n13525) );
  DFFARX1 \rf/conf6_reg[15]  ( .D(n17866), .CLK(clock), .RSTB(n34684), .Q(
        n34565), .QN(n13469) );
  DFFARX1 \rf/conf5_reg[0]  ( .D(n17909), .CLK(clock), .RSTB(n34684), .Q(
        n34344), .QN(n13890) );
  DFFARX1 \rf/conf5_reg[1]  ( .D(n17908), .CLK(clock), .RSTB(n34684), .Q(
        n34493), .QN(n13862) );
  DFFARX1 \rf/conf5_reg[2]  ( .D(n17907), .CLK(clock), .RSTB(n34684), .Q(
        n34343), .QN(n13836) );
  DFFARX1 \rf/conf5_reg[3]  ( .D(n17906), .CLK(clock), .RSTB(n34684), .Q(
        n34494), .QN(n13810) );
  DFFARX1 \rf/conf5_reg[4]  ( .D(n17905), .CLK(clock), .RSTB(n34684), .Q(
        n34587), .QN(n13784) );
  DFFARX1 \rf/conf5_reg[5]  ( .D(n17904), .CLK(clock), .RSTB(n34684), .Q(
        n34370), .QN(n13758) );
  DFFARX1 \rf/conf5_reg[6]  ( .D(n17903), .CLK(clock), .RSTB(n34684), .Q(
        n34317), .QN(n13732) );
  DFFARX1 \rf/conf5_reg[7]  ( .D(n17902), .CLK(clock), .RSTB(n34684), .Q(
        n34495), .QN(n13706) );
  DFFARX1 \rf/conf5_reg[8]  ( .D(n17901), .CLK(clock), .RSTB(n34684), .Q(
        n34235), .QN(n13680) );
  DFFARX1 \rf/conf5_reg[9]  ( .D(n17900), .CLK(clock), .RSTB(n34685), .Q(
        n34496), .QN(n13654) );
  DFFARX1 \rf/conf5_reg[10]  ( .D(n17899), .CLK(clock), .RSTB(n34685), .Q(
        n34342), .QN(n13628) );
  DFFARX1 \rf/conf5_reg[11]  ( .D(n17898), .CLK(clock), .RSTB(n34685), .Q(
        n34528), .QN(n13602) );
  DFFARX1 \rf/conf5_reg[12]  ( .D(n17897), .CLK(clock), .RSTB(n34685), .Q(
        n34341), .QN(n13576) );
  DFFARX1 \rf/conf5_reg[13]  ( .D(n17896), .CLK(clock), .RSTB(n34685), .Q(
        n34529), .QN(n13550) );
  DFFARX1 \rf/conf5_reg[14]  ( .D(n17895), .CLK(clock), .RSTB(n34685), .Q(
        n34316), .QN(n13524) );
  DFFARX1 \rf/conf5_reg[15]  ( .D(n17894), .CLK(clock), .RSTB(n34685), .Q(
        n34530), .QN(n13465) );
  DFFARX1 \rf/conf4_reg[0]  ( .D(n17937), .CLK(clock), .RSTB(n34685), .Q(
        n34340), .QN(n13888) );
  DFFARX1 \rf/conf4_reg[1]  ( .D(n17936), .CLK(clock), .RSTB(n34685), .Q(
        n34490), .QN(n13861) );
  DFFARX1 \rf/conf4_reg[2]  ( .D(n17935), .CLK(clock), .RSTB(n34685), .Q(
        n34315), .QN(n13835) );
  DFFARX1 \rf/conf4_reg[3]  ( .D(n17934), .CLK(clock), .RSTB(n34685), .Q(
        n34491), .QN(n13809) );
  DFFARX1 \rf/conf4_reg[4]  ( .D(n17933), .CLK(clock), .RSTB(n34685), .Q(
        n34627), .QN(n13783) );
  DFFARX1 \rf/conf4_reg[5]  ( .D(n17932), .CLK(clock), .RSTB(n34686), .Q(
        n34577), .QN(n13757) );
  DFFARX1 \rf/conf4_reg[6]  ( .D(n17931), .CLK(clock), .RSTB(n34686), .Q(
        n34617), .QN(n13731) );
  DFFARX1 \rf/conf4_reg[7]  ( .D(n17930), .CLK(clock), .RSTB(n34686), .Q(
        n34578), .QN(n13705) );
  DFFARX1 \rf/conf4_reg[8]  ( .D(n17929), .CLK(clock), .RSTB(n34686), .Q(
        n34338), .QN(n13679) );
  DFFARX1 \rf/conf4_reg[9]  ( .D(n17928), .CLK(clock), .RSTB(n34686), .Q(
        n34525), .QN(n13653) );
  DFFARX1 \rf/conf4_reg[10]  ( .D(n17927), .CLK(clock), .RSTB(n34686), .Q(
        n34313), .QN(n13627) );
  DFFARX1 \rf/conf4_reg[11]  ( .D(n17926), .CLK(clock), .RSTB(n34686), .Q(
        n34492), .QN(n13601) );
  DFFARX1 \rf/conf4_reg[12]  ( .D(n17925), .CLK(clock), .RSTB(n34686), .Q(
        n34339), .QN(n13575) );
  DFFARX1 \rf/conf4_reg[13]  ( .D(n17924), .CLK(clock), .RSTB(n34686), .Q(
        n34526), .QN(n13549) );
  DFFARX1 \rf/conf4_reg[14]  ( .D(n17923), .CLK(clock), .RSTB(n34686), .Q(
        n34314), .QN(n13523) );
  DFFARX1 \rf/conf4_reg[15]  ( .D(n17922), .CLK(clock), .RSTB(n34686), .Q(
        n34527), .QN(n13464) );
  DFFARX1 \rf/conf3_reg[0]  ( .D(n17965), .CLK(clock), .RSTB(n34687), .Q(
        n34309), .QN(n13902) );
  DFFARX1 \rf/conf3_reg[1]  ( .D(n17964), .CLK(clock), .RSTB(n34687), .Q(
        n34485), .QN(n13868) );
  DFFARX1 \rf/conf3_reg[2]  ( .D(n17963), .CLK(clock), .RSTB(n34687), .Q(
        n34310), .QN(n13842) );
  DFFARX1 \rf/conf3_reg[3]  ( .D(n17962), .CLK(clock), .RSTB(n34687), .Q(
        n34486), .QN(n13816) );
  DFFARX1 \rf/conf3_reg[4]  ( .D(n17961), .CLK(clock), .RSTB(n34687), .Q(
        n34637), .QN(n13790) );
  DFFARX1 \rf/conf3_reg[5]  ( .D(n17960), .CLK(clock), .RSTB(n34687), .Q(
        n34595), .QN(n13764) );
  DFFARX1 \rf/conf3_reg[6]  ( .D(n17959), .CLK(clock), .RSTB(n34687), .Q(
        n34616), .QN(n13738) );
  DFFARX1 \rf/conf3_reg[7]  ( .D(n17958), .CLK(clock), .RSTB(n34677), .Q(
        n34564), .QN(n13712) );
  DFFARX1 \rf/conf3_reg[8]  ( .D(n17957), .CLK(clock), .RSTB(n34687), .Q(
        n34236), .QN(n13686) );
  DFFARX1 \rf/conf3_reg[9]  ( .D(n17956), .CLK(clock), .RSTB(n34687), .Q(
        n34487), .QN(n13660) );
  DFFARX1 \rf/conf3_reg[10]  ( .D(n17955), .CLK(clock), .RSTB(n34687), .Q(
        n34361), .QN(n13634) );
  DFFARX1 \rf/conf3_reg[11]  ( .D(n17954), .CLK(clock), .RSTB(n34687), .Q(
        n34551), .QN(n13608) );
  DFFARX1 \rf/conf3_reg[12]  ( .D(n17953), .CLK(clock), .RSTB(n34687), .Q(
        n34311), .QN(n13582) );
  DFFARX1 \rf/conf3_reg[13]  ( .D(n17952), .CLK(clock), .RSTB(n34688), .Q(
        n34488), .QN(n13556) );
  DFFARX1 \rf/conf3_reg[14]  ( .D(n17951), .CLK(clock), .RSTB(n34688), .Q(
        n34312), .QN(n13530) );
  DFFARX1 \rf/conf3_reg[15]  ( .D(n17950), .CLK(clock), .RSTB(n34688), .Q(
        n34489), .QN(n13475) );
  DFFARX1 \rf/conf2_reg[0]  ( .D(n17993), .CLK(clock), .RSTB(n34688), .Q(
        n34308), .QN(n13900) );
  DFFARX1 \rf/conf2_reg[1]  ( .D(n17992), .CLK(clock), .RSTB(n34688), .Q(
        n34523), .QN(n13867) );
  DFFARX1 \rf/conf2_reg[2]  ( .D(n17991), .CLK(clock), .RSTB(n34688), .Q(
        n34337), .QN(n13841) );
  DFFARX1 \rf/conf2_reg[3]  ( .D(n17990), .CLK(clock), .RSTB(n34688), .Q(
        n34524), .QN(n13815) );
  DFFARX1 \rf/conf2_reg[4]  ( .D(n17989), .CLK(clock), .RSTB(n34688), .Q(
        n34626), .QN(n13789) );
  DFFARX1 \rf/conf2_reg[5]  ( .D(n17988), .CLK(clock), .RSTB(n34688), .Q(
        n34563), .QN(n13763) );
  DFFARX1 \rf/conf2_reg[6]  ( .D(n17987), .CLK(clock), .RSTB(n34688), .Q(
        n34479), .QN(n13737) );
  DFFARX1 \rf/conf2_reg[7]  ( .D(n17986), .CLK(clock), .RSTB(n34688), .Q(
        n34647), .QN(n13711) );
  DFFARX1 \rf/conf2_reg[8]  ( .D(n17985), .CLK(clock), .RSTB(n34688), .Q(
        n34605), .QN(n13685) );
  DFFARX1 \rf/conf2_reg[9]  ( .D(n17984), .CLK(clock), .RSTB(n34689), .Q(
        n34373), .QN(n13659) );
  DFFARX1 \rf/conf2_reg[10]  ( .D(n17983), .CLK(clock), .RSTB(n34689), .Q(
        n34307), .QN(n13633) );
  DFFARX1 \rf/conf2_reg[11]  ( .D(n17982), .CLK(clock), .RSTB(n34689), .Q(
        n34484), .QN(n13607) );
  DFFARX1 \rf/conf2_reg[12]  ( .D(n17981), .CLK(clock), .RSTB(n34689), .Q(
        n34615), .QN(n13581) );
  DFFARX1 \rf/conf2_reg[13]  ( .D(n17980), .CLK(clock), .RSTB(n34689), .Q(
        n34576), .QN(n13555) );
  DFFARX1 \rf/conf2_reg[14]  ( .D(n17979), .CLK(clock), .RSTB(n34689), .Q(
        n34478), .QN(n13529) );
  DFFARX1 \rf/conf2_reg[15]  ( .D(n17978), .CLK(clock), .RSTB(n34689), .Q(
        n34641), .QN(n13474) );
  DFFARX1 \rf/conf1_reg[0]  ( .D(n18021), .CLK(clock), .RSTB(n34689), .Q(
        n34294), .QN(n13898) );
  DFFARX1 \rf/conf1_reg[1]  ( .D(n18020), .CLK(clock), .RSTB(n34689), .Q(
        n34557), .QN(n13866) );
  DFFARX1 \rf/conf1_reg[2]  ( .D(n18019), .CLK(clock), .RSTB(n34689), .Q(
        n34293), .QN(n13840) );
  DFFARX1 \rf/conf1_reg[3]  ( .D(n18018), .CLK(clock), .RSTB(n34689), .Q(
        n34555), .QN(n13814) );
  DFFARX1 \rf/conf1_reg[4]  ( .D(n18017), .CLK(clock), .RSTB(n34689), .Q(
        n34297), .QN(n13788) );
  DFFARX1 \rf/conf1_reg[5]  ( .D(n18016), .CLK(clock), .RSTB(n34690), .Q(
        n34558), .QN(n13762) );
  DFFARX1 \rf/conf1_reg[6]  ( .D(n18015), .CLK(clock), .RSTB(n34690), .Q(
        n34335), .QN(n13736) );
  DFFARX1 \rf/conf1_reg[7]  ( .D(n18014), .CLK(clock), .RSTB(n34690), .Q(
        n34521), .QN(n13710) );
  DFFARX1 \rf/conf1_reg[8]  ( .D(n18013), .CLK(clock), .RSTB(n34690), .Q(
        n34336), .QN(n13684) );
  DFFARX1 \rf/conf1_reg[9]  ( .D(n18012), .CLK(clock), .RSTB(n34690), .Q(
        n34483), .QN(n13658) );
  DFFARX1 \rf/conf1_reg[10]  ( .D(n18011), .CLK(clock), .RSTB(n34690), .Q(
        n34295), .QN(n13632) );
  DFFARX1 \rf/conf1_reg[11]  ( .D(n18010), .CLK(clock), .RSTB(n34690), .Q(
        n34556), .QN(n13606) );
  DFFARX1 \rf/conf1_reg[12]  ( .D(n18009), .CLK(clock), .RSTB(n34690), .Q(
        n34306), .QN(n13580) );
  DFFARX1 \rf/conf1_reg[13]  ( .D(n18008), .CLK(clock), .RSTB(n34690), .Q(
        n34522), .QN(n13554) );
  DFFARX1 \rf/conf1_reg[14]  ( .D(n18007), .CLK(clock), .RSTB(n34690), .Q(
        n34296), .QN(n13528) );
  DFFARX1 \rf/conf1_reg[15]  ( .D(n18006), .CLK(clock), .RSTB(n34690), .Q(
        n34559), .QN(n13472) );
  DFFARX1 \rf/conf0_reg[0]  ( .D(n18049), .CLK(clock), .RSTB(n34690), .Q(
        n34623), .QN(n13896) );
  DFFARX1 \rf/conf0_reg[1]  ( .D(n18048), .CLK(clock), .RSTB(n34691), .Q(
        n34572), .QN(n13865) );
  DFFARX1 \rf/conf0_reg[2]  ( .D(n18047), .CLK(clock), .RSTB(n34691), .Q(
        n34624), .QN(n13839) );
  DFFARX1 \rf/conf0_reg[3]  ( .D(n18046), .CLK(clock), .RSTB(n34691), .Q(
        n34573), .QN(n13813) );
  DFFARX1 \rf/conf0_reg[4]  ( .D(n18045), .CLK(clock), .RSTB(n34691), .Q(
        n34612), .QN(n13787) );
  DFFARX1 \rf/conf0_reg[5]  ( .D(n18044), .CLK(clock), .RSTB(n34691), .Q(
        n34574), .QN(n13761) );
  DFFARX1 \rf/conf0_reg[6]  ( .D(n18043), .CLK(clock), .RSTB(n34691), .Q(
        n34613), .QN(n13735) );
  DFFARX1 \rf/conf0_reg[7]  ( .D(n18042), .CLK(clock), .RSTB(n34691), .Q(
        n34561), .QN(n13709) );
  DFFARX1 \rf/conf0_reg[8]  ( .D(n18041), .CLK(clock), .RSTB(n34691), .Q(
        n34304), .QN(n13683) );
  DFFARX1 \rf/conf0_reg[9]  ( .D(n18040), .CLK(clock), .RSTB(n34691), .Q(
        n34519), .QN(n13657) );
  DFFARX1 \rf/conf0_reg[10]  ( .D(n18039), .CLK(clock), .RSTB(n34691), .Q(
        n34305), .QN(n13631) );
  DFFARX1 \rf/conf0_reg[11]  ( .D(n18038), .CLK(clock), .RSTB(n34691), .Q(
        n34520), .QN(n13605) );
  DFFARX1 \rf/conf0_reg[12]  ( .D(n18037), .CLK(clock), .RSTB(n34691), .Q(
        n34614), .QN(n13579) );
  DFFARX1 \rf/conf0_reg[13]  ( .D(n18036), .CLK(clock), .RSTB(n34692), .Q(
        n34575), .QN(n13553) );
  DFFARX1 \rf/conf0_reg[14]  ( .D(n18035), .CLK(clock), .RSTB(n34687), .Q(
        n34625), .QN(n13527) );
  DFFARX1 \rf/conf0_reg[15]  ( .D(n18034), .CLK(clock), .RSTB(n34683), .Q(
        n34562), .QN(n13471) );
  NAND2X0 U19373 ( .IN1(n18209), .IN2(n18212), .QN(n18210) );
  NAND2X0 U19374 ( .IN1(n18209), .IN2(n18208), .QN(n18216) );
  NAND2X0 U19375 ( .IN1(n18213), .IN2(n18212), .QN(n18215) );
  INVX0 U19376 ( .INP(n32343), .ZN(n32324) );
  NOR2X0 U19377 ( .IN1(n34378), .IN2(n30857), .QN(n18203) );
  NAND2X0 U19378 ( .IN1(n18213), .IN2(n18208), .QN(n18211) );
  NAND2X0 U19379 ( .IN1(n18199), .IN2(n18200), .QN(n32889) );
  NOR2X0 U19380 ( .IN1(n34249), .IN2(n32886), .QN(n18199) );
  NAND2X0 U19381 ( .IN1(n32902), .IN2(n32911), .QN(n18200) );
  NAND2X0 U19382 ( .IN1(n18203), .IN2(n18204), .QN(n30862) );
  NAND2X0 U19383 ( .IN1(n30859), .IN2(n30858), .QN(n18204) );
  INVX0 U19384 ( .INP(n30560), .ZN(n30551) );
  NAND2X0 U19385 ( .IN1(n18206), .IN2(n18207), .QN(n29533) );
  NAND2X0 U19386 ( .IN1(n29530), .IN2(n29529), .QN(n18207) );
  NOR2X0 U19387 ( .IN1(n34250), .IN2(n29528), .QN(n18206) );
  INVX0 U19388 ( .INP(n32983), .ZN(n32946) );
  NOR2X0 U19389 ( .IN1(n31374), .IN2(n31435), .QN(n18201) );
  NAND2X0 U19390 ( .IN1(n31376), .IN2(n31375), .QN(n18202) );
  NAND2X0 U19391 ( .IN1(n18205), .IN2(\s2/msel/gnt_p1 [0]), .QN(n30157) );
  NOR2X0 U19392 ( .IN1(n30129), .IN2(n34383), .QN(n18205) );
  NAND2X0 U19393 ( .IN1(n18201), .IN2(n18202), .QN(n31377) );
  OR4X1 U19394 ( .IN1(n18904), .IN2(n34080), .IN3(n18903), .IN4(n30004), .Q(
        n18194) );
  OAI21X1 U19395 ( .IN1(n31673), .IN2(n31658), .IN3(n31657), .QN(n18195) );
  INVX0 U19396 ( .INP(n29661), .ZN(n29645) );
  OR2X1 U19397 ( .IN1(n31986), .IN2(n31985), .Q(n18196) );
  OR3X1 U19398 ( .IN1(n18883), .IN2(n32034), .IN3(n18882), .Q(n18197) );
  AND2X1 U19399 ( .IN1(n31187), .IN2(n31186), .Q(n18198) );
  INVX0 U19400 ( .INP(rst_i), .ZN(n34694) );
  INVX0 U19401 ( .INP(rst_i), .ZN(n34679) );
  INVX0 U19402 ( .INP(rst_i), .ZN(n34695) );
  INVX0 U19403 ( .INP(rst_i), .ZN(n34696) );
  INVX0 U19404 ( .INP(rst_i), .ZN(n34697) );
  INVX0 U19405 ( .INP(rst_i), .ZN(n34681) );
  INVX0 U19406 ( .INP(rst_i), .ZN(n34677) );
  INVX0 U19407 ( .INP(rst_i), .ZN(n34692) );
  INVX0 U19408 ( .INP(rst_i), .ZN(n34678) );
  INVX0 U19409 ( .INP(rst_i), .ZN(n34693) );
  INVX0 U19410 ( .INP(rst_i), .ZN(n34687) );
  INVX0 U19411 ( .INP(rst_i), .ZN(n34688) );
  INVX0 U19412 ( .INP(rst_i), .ZN(n34689) );
  INVX0 U19413 ( .INP(rst_i), .ZN(n34690) );
  INVX0 U19414 ( .INP(rst_i), .ZN(n34691) );
  INVX0 U19415 ( .INP(rst_i), .ZN(n34680) );
  INVX0 U19416 ( .INP(rst_i), .ZN(n34682) );
  INVX0 U19417 ( .INP(rst_i), .ZN(n34683) );
  INVX0 U19418 ( .INP(rst_i), .ZN(n34684) );
  INVX0 U19419 ( .INP(rst_i), .ZN(n34686) );
  INVX0 U19420 ( .INP(rst_i), .ZN(n34685) );
  MUX41X1 U19421 ( .IN1(\s15/msel/gnt_p0 [0]), .IN3(\s15/msel/gnt_p2 [0]), 
        .IN2(\s15/msel/gnt_p1 [0]), .IN4(\s15/msel/gnt_p3 [0]), .S0(
        \s15/msel/pri_out [1]), .S1(\s15/msel/pri_out [0]), .Q(n18217) );
  INVX0 U19422 ( .INP(n18217), .ZN(n18214) );
  MUX41X1 U19423 ( .IN1(\s15/msel/gnt_p0 [1]), .IN3(\s15/msel/gnt_p2 [1]), 
        .IN2(\s15/msel/gnt_p1 [1]), .IN4(\s15/msel/gnt_p3 [1]), .S0(
        \s15/msel/pri_out [1]), .S1(\s15/msel/pri_out [0]), .Q(n18209) );
  MUX41X1 U19424 ( .IN1(\s15/msel/gnt_p0 [2]), .IN3(\s15/msel/gnt_p2 [2]), 
        .IN2(\s15/msel/gnt_p1 [2]), .IN4(\s15/msel/gnt_p3 [2]), .S0(
        \s15/msel/pri_out [1]), .S1(\s15/msel/pri_out [0]), .Q(n18212) );
  INVX0 U19425 ( .INP(n18212), .ZN(n18208) );
  NOR2X0 U19426 ( .IN1(n18214), .IN2(n18216), .QN(n18239) );
  INVX0 U19427 ( .INP(n18239), .ZN(n23812) );
  INVX0 U19428 ( .INP(m3s0_addr[4]), .ZN(n28618) );
  INVX0 U19429 ( .INP(n18209), .ZN(n18213) );
  NOR2X0 U19430 ( .IN1(n18214), .IN2(n18211), .QN(n18246) );
  INVX0 U19431 ( .INP(n18246), .ZN(n23831) );
  INVX0 U19432 ( .INP(m1s0_addr[4]), .ZN(n28616) );
  OA22X1 U19433 ( .IN1(n23812), .IN2(n28618), .IN3(n23831), .IN4(n28616), .Q(
        n18221) );
  NOR2X0 U19434 ( .IN1(n18214), .IN2(n18210), .QN(n18230) );
  INVX0 U19435 ( .INP(n18230), .ZN(n23834) );
  INVX0 U19436 ( .INP(m7s0_addr[4]), .ZN(n28619) );
  NOR2X0 U19437 ( .IN1(n18217), .IN2(n18210), .QN(n18231) );
  INVX0 U19438 ( .INP(n18231), .ZN(n23833) );
  INVX0 U19439 ( .INP(m6s0_addr[4]), .ZN(n28620) );
  OA22X1 U19440 ( .IN1(n23834), .IN2(n28619), .IN3(n23833), .IN4(n28620), .Q(
        n18220) );
  NOR2X0 U19441 ( .IN1(n18217), .IN2(n18211), .QN(n18237) );
  INVX0 U19442 ( .INP(n18237), .ZN(n23823) );
  INVX0 U19443 ( .INP(m0s0_addr[4]), .ZN(n28617) );
  NOR2X0 U19444 ( .IN1(n18214), .IN2(n18215), .QN(n18247) );
  INVX0 U19445 ( .INP(n18247), .ZN(n23832) );
  INVX0 U19446 ( .INP(m5s0_addr[4]), .ZN(n28614) );
  OA22X1 U19447 ( .IN1(n23823), .IN2(n28617), .IN3(n23832), .IN4(n28614), .Q(
        n18219) );
  NOR2X0 U19448 ( .IN1(n18217), .IN2(n18215), .QN(n18238) );
  INVX0 U19449 ( .INP(n18238), .ZN(n23836) );
  INVX0 U19450 ( .INP(m4s0_addr[4]), .ZN(n28615) );
  NOR2X0 U19451 ( .IN1(n18217), .IN2(n18216), .QN(n18232) );
  INVX0 U19452 ( .INP(n18232), .ZN(n23817) );
  INVX0 U19453 ( .INP(m2s0_addr[4]), .ZN(n28613) );
  OA22X1 U19454 ( .IN1(n23836), .IN2(n28615), .IN3(n23817), .IN4(n28613), .Q(
        n18218) );
  NAND4X0 U19455 ( .IN1(n18221), .IN2(n18220), .IN3(n18219), .IN4(n18218), 
        .QN(s15_addr_o[4]) );
  INVX0 U19456 ( .INP(n18231), .ZN(n23799) );
  INVX0 U19457 ( .INP(m6s0_addr[5]), .ZN(n28628) );
  INVX0 U19458 ( .INP(m2s0_addr[5]), .ZN(n28632) );
  OA22X1 U19459 ( .IN1(n23799), .IN2(n28628), .IN3(n23817), .IN4(n28632), .Q(
        n18225) );
  INVX0 U19460 ( .INP(m5s0_addr[5]), .ZN(n28627) );
  INVX0 U19461 ( .INP(n18239), .ZN(n23835) );
  INVX0 U19462 ( .INP(m3s0_addr[5]), .ZN(n28626) );
  OA22X1 U19463 ( .IN1(n23832), .IN2(n28627), .IN3(n23835), .IN4(n28626), .Q(
        n18224) );
  INVX0 U19464 ( .INP(m4s0_addr[5]), .ZN(n28631) );
  INVX0 U19465 ( .INP(m1s0_addr[5]), .ZN(n28630) );
  OA22X1 U19466 ( .IN1(n23836), .IN2(n28631), .IN3(n23831), .IN4(n28630), .Q(
        n18223) );
  INVX0 U19467 ( .INP(n18237), .ZN(n23838) );
  INVX0 U19468 ( .INP(m0s0_addr[5]), .ZN(n28629) );
  INVX0 U19469 ( .INP(n18230), .ZN(n23824) );
  INVX0 U19470 ( .INP(m7s0_addr[5]), .ZN(n28625) );
  OA22X1 U19471 ( .IN1(n23838), .IN2(n28629), .IN3(n23824), .IN4(n28625), .Q(
        n18222) );
  NAND4X0 U19472 ( .IN1(n18225), .IN2(n18224), .IN3(n18223), .IN4(n18222), 
        .QN(s15_addr_o[5]) );
  INVX0 U19473 ( .INP(m5s0_addr[3]), .ZN(n28602) );
  INVX0 U19474 ( .INP(n18232), .ZN(n23837) );
  INVX0 U19475 ( .INP(m2s0_addr[3]), .ZN(n28604) );
  OA22X1 U19476 ( .IN1(n23832), .IN2(n28602), .IN3(n23837), .IN4(n28604), .Q(
        n18229) );
  INVX0 U19477 ( .INP(n18238), .ZN(n23825) );
  INVX0 U19478 ( .INP(m4s0_addr[3]), .ZN(n28606) );
  INVX0 U19479 ( .INP(m1s0_addr[3]), .ZN(n28605) );
  OA22X1 U19480 ( .IN1(n23825), .IN2(n28606), .IN3(n23831), .IN4(n28605), .Q(
        n18228) );
  INVX0 U19481 ( .INP(m0s0_addr[3]), .ZN(n28601) );
  INVX0 U19482 ( .INP(m6s0_addr[3]), .ZN(n28603) );
  OA22X1 U19483 ( .IN1(n23823), .IN2(n28601), .IN3(n23833), .IN4(n28603), .Q(
        n18227) );
  INVX0 U19484 ( .INP(m3s0_addr[3]), .ZN(n28607) );
  INVX0 U19485 ( .INP(m7s0_addr[3]), .ZN(n28608) );
  OA22X1 U19486 ( .IN1(n23835), .IN2(n28607), .IN3(n23824), .IN4(n28608), .Q(
        n18226) );
  NAND4X0 U19487 ( .IN1(n18229), .IN2(n18228), .IN3(n18227), .IN4(n18226), 
        .QN(s15_addr_o[3]) );
  NAND3X0 U19488 ( .IN1(m7s15_cyc), .IN2(n18230), .IN3(\s15/m7_cyc_r ), .QN(
        n18236) );
  NAND3X0 U19489 ( .IN1(m6s15_cyc), .IN2(n18231), .IN3(\s15/m6_cyc_r ), .QN(
        n18235) );
  NAND3X0 U19490 ( .IN1(m1s15_cyc), .IN2(n18246), .IN3(\s15/m1_cyc_r ), .QN(
        n18234) );
  NAND3X0 U19491 ( .IN1(m2s15_cyc), .IN2(n18232), .IN3(\s15/m2_cyc_r ), .QN(
        n18233) );
  NAND4X0 U19492 ( .IN1(n18236), .IN2(n18235), .IN3(n18234), .IN4(n18233), 
        .QN(n18245) );
  NAND3X0 U19493 ( .IN1(m0s15_cyc), .IN2(n18237), .IN3(\s15/m0_cyc_r ), .QN(
        n18243) );
  NAND3X0 U19494 ( .IN1(m4s15_cyc), .IN2(n18238), .IN3(\s15/m4_cyc_r ), .QN(
        n18242) );
  NAND3X0 U19495 ( .IN1(m5s15_cyc), .IN2(n18247), .IN3(\s15/m5_cyc_r ), .QN(
        n18241) );
  NAND3X0 U19496 ( .IN1(m3s15_cyc), .IN2(n18239), .IN3(\s15/m3_cyc_r ), .QN(
        n18240) );
  NAND4X0 U19497 ( .IN1(n18243), .IN2(n18242), .IN3(n18241), .IN4(n18240), 
        .QN(n18244) );
  NOR2X0 U19498 ( .IN1(n18245), .IN2(n18244), .QN(n18178) );
  INVX0 U19499 ( .INP(m0s0_data_o[0]), .ZN(n28134) );
  INVX0 U19500 ( .INP(m3s0_data_o[0]), .ZN(n28139) );
  OA22X1 U19501 ( .IN1(n23823), .IN2(n28134), .IN3(n23812), .IN4(n28139), .Q(
        n18251) );
  INVX0 U19502 ( .INP(m4s0_data_o[0]), .ZN(n28138) );
  INVX0 U19503 ( .INP(n18246), .ZN(n23818) );
  INVX0 U19504 ( .INP(m1s0_data_o[0]), .ZN(n28140) );
  OA22X1 U19505 ( .IN1(n23825), .IN2(n28138), .IN3(n23818), .IN4(n28140), .Q(
        n18250) );
  INVX0 U19506 ( .INP(m7s0_data_o[0]), .ZN(n28135) );
  INVX0 U19507 ( .INP(m6s0_data_o[0]), .ZN(n28137) );
  OA22X1 U19508 ( .IN1(n23824), .IN2(n28135), .IN3(n23833), .IN4(n28137), .Q(
        n18249) );
  INVX0 U19509 ( .INP(n18247), .ZN(n23826) );
  INVX0 U19510 ( .INP(m5s0_data_o[0]), .ZN(n28136) );
  INVX0 U19511 ( .INP(m2s0_data_o[0]), .ZN(n28133) );
  OA22X1 U19512 ( .IN1(n23826), .IN2(n28136), .IN3(n23837), .IN4(n28133), .Q(
        n18248) );
  NAND4X0 U19513 ( .IN1(n18251), .IN2(n18250), .IN3(n18249), .IN4(n18248), 
        .QN(s15_data_o[0]) );
  INVX0 U19514 ( .INP(m4s0_data_o[1]), .ZN(n28149) );
  INVX0 U19515 ( .INP(m5s0_data_o[1]), .ZN(n28152) );
  OA22X1 U19516 ( .IN1(n23836), .IN2(n28149), .IN3(n23826), .IN4(n28152), .Q(
        n18255) );
  INVX0 U19517 ( .INP(m0s0_data_o[1]), .ZN(n28150) );
  INVX0 U19518 ( .INP(m6s0_data_o[1]), .ZN(n28151) );
  OA22X1 U19519 ( .IN1(n23838), .IN2(n28150), .IN3(n23833), .IN4(n28151), .Q(
        n18254) );
  INVX0 U19520 ( .INP(m7s0_data_o[1]), .ZN(n28147) );
  INVX0 U19521 ( .INP(m1s0_data_o[1]), .ZN(n28146) );
  OA22X1 U19522 ( .IN1(n23834), .IN2(n28147), .IN3(n23831), .IN4(n28146), .Q(
        n18253) );
  INVX0 U19523 ( .INP(m3s0_data_o[1]), .ZN(n28145) );
  INVX0 U19524 ( .INP(m2s0_data_o[1]), .ZN(n28148) );
  OA22X1 U19525 ( .IN1(n23812), .IN2(n28145), .IN3(n23837), .IN4(n28148), .Q(
        n18252) );
  NAND4X0 U19526 ( .IN1(n18255), .IN2(n18254), .IN3(n18253), .IN4(n18252), 
        .QN(s15_data_o[1]) );
  INVX0 U19527 ( .INP(m0s0_data_o[2]), .ZN(n28160) );
  INVX0 U19528 ( .INP(m4s0_data_o[2]), .ZN(n28158) );
  OA22X1 U19529 ( .IN1(n23823), .IN2(n28160), .IN3(n23825), .IN4(n28158), .Q(
        n18259) );
  INVX0 U19530 ( .INP(m5s0_data_o[2]), .ZN(n28162) );
  INVX0 U19531 ( .INP(m6s0_data_o[2]), .ZN(n28157) );
  OA22X1 U19532 ( .IN1(n23832), .IN2(n28162), .IN3(n23833), .IN4(n28157), .Q(
        n18258) );
  INVX0 U19533 ( .INP(m3s0_data_o[2]), .ZN(n28159) );
  INVX0 U19534 ( .INP(m2s0_data_o[2]), .ZN(n28163) );
  OA22X1 U19535 ( .IN1(n23835), .IN2(n28159), .IN3(n23837), .IN4(n28163), .Q(
        n18257) );
  INVX0 U19536 ( .INP(m7s0_data_o[2]), .ZN(n28161) );
  INVX0 U19537 ( .INP(m1s0_data_o[2]), .ZN(n28164) );
  OA22X1 U19538 ( .IN1(n23824), .IN2(n28161), .IN3(n23818), .IN4(n28164), .Q(
        n18256) );
  NAND4X0 U19539 ( .IN1(n18259), .IN2(n18258), .IN3(n18257), .IN4(n18256), 
        .QN(s15_data_o[2]) );
  INVX0 U19540 ( .INP(m3s0_data_o[3]), .ZN(n28170) );
  INVX0 U19541 ( .INP(m1s0_data_o[3]), .ZN(n28174) );
  OA22X1 U19542 ( .IN1(n23812), .IN2(n28170), .IN3(n23818), .IN4(n28174), .Q(
        n18263) );
  INVX0 U19543 ( .INP(m0s0_data_o[3]), .ZN(n28172) );
  INVX0 U19544 ( .INP(m7s0_data_o[3]), .ZN(n28173) );
  OA22X1 U19545 ( .IN1(n23823), .IN2(n28172), .IN3(n23824), .IN4(n28173), .Q(
        n18262) );
  INVX0 U19546 ( .INP(m4s0_data_o[3]), .ZN(n28171) );
  INVX0 U19547 ( .INP(m6s0_data_o[3]), .ZN(n28169) );
  OA22X1 U19548 ( .IN1(n23825), .IN2(n28171), .IN3(n23833), .IN4(n28169), .Q(
        n18261) );
  INVX0 U19549 ( .INP(m5s0_data_o[3]), .ZN(n28175) );
  INVX0 U19550 ( .INP(m2s0_data_o[3]), .ZN(n28176) );
  OA22X1 U19551 ( .IN1(n23826), .IN2(n28175), .IN3(n23837), .IN4(n28176), .Q(
        n18260) );
  NAND4X0 U19552 ( .IN1(n18263), .IN2(n18262), .IN3(n18261), .IN4(n18260), 
        .QN(s15_data_o[3]) );
  INVX0 U19553 ( .INP(m0s0_data_o[4]), .ZN(n28182) );
  INVX0 U19554 ( .INP(m4s0_data_o[4]), .ZN(n28185) );
  OA22X1 U19555 ( .IN1(n23823), .IN2(n28182), .IN3(n23825), .IN4(n28185), .Q(
        n18267) );
  INVX0 U19556 ( .INP(m5s0_data_o[4]), .ZN(n28183) );
  INVX0 U19557 ( .INP(m7s0_data_o[4]), .ZN(n28181) );
  OA22X1 U19558 ( .IN1(n23832), .IN2(n28183), .IN3(n23824), .IN4(n28181), .Q(
        n18266) );
  INVX0 U19559 ( .INP(m3s0_data_o[4]), .ZN(n28188) );
  INVX0 U19560 ( .INP(m2s0_data_o[4]), .ZN(n28186) );
  OA22X1 U19561 ( .IN1(n23835), .IN2(n28188), .IN3(n23837), .IN4(n28186), .Q(
        n18265) );
  INVX0 U19562 ( .INP(m6s0_data_o[4]), .ZN(n28187) );
  INVX0 U19563 ( .INP(m1s0_data_o[4]), .ZN(n28184) );
  OA22X1 U19564 ( .IN1(n23799), .IN2(n28187), .IN3(n23831), .IN4(n28184), .Q(
        n18264) );
  NAND4X0 U19565 ( .IN1(n18267), .IN2(n18266), .IN3(n18265), .IN4(n18264), 
        .QN(s15_data_o[4]) );
  INVX0 U19566 ( .INP(m0s0_data_o[5]), .ZN(n28196) );
  INVX0 U19567 ( .INP(m7s0_data_o[5]), .ZN(n28199) );
  OA22X1 U19568 ( .IN1(n23838), .IN2(n28196), .IN3(n23834), .IN4(n28199), .Q(
        n18271) );
  INVX0 U19569 ( .INP(m3s0_data_o[5]), .ZN(n28193) );
  INVX0 U19570 ( .INP(m1s0_data_o[5]), .ZN(n28200) );
  OA22X1 U19571 ( .IN1(n23812), .IN2(n28193), .IN3(n23818), .IN4(n28200), .Q(
        n18270) );
  INVX0 U19572 ( .INP(m4s0_data_o[5]), .ZN(n28198) );
  INVX0 U19573 ( .INP(m6s0_data_o[5]), .ZN(n28195) );
  OA22X1 U19574 ( .IN1(n23836), .IN2(n28198), .IN3(n23833), .IN4(n28195), .Q(
        n18269) );
  INVX0 U19575 ( .INP(m5s0_data_o[5]), .ZN(n28197) );
  INVX0 U19576 ( .INP(m2s0_data_o[5]), .ZN(n28194) );
  OA22X1 U19577 ( .IN1(n23826), .IN2(n28197), .IN3(n23837), .IN4(n28194), .Q(
        n18268) );
  NAND4X0 U19578 ( .IN1(n18271), .IN2(n18270), .IN3(n18269), .IN4(n18268), 
        .QN(s15_data_o[5]) );
  INVX0 U19579 ( .INP(m3s0_data_o[6]), .ZN(n28212) );
  INVX0 U19580 ( .INP(m6s0_data_o[6]), .ZN(n28210) );
  OA22X1 U19581 ( .IN1(n23835), .IN2(n28212), .IN3(n23833), .IN4(n28210), .Q(
        n18275) );
  INVX0 U19582 ( .INP(m1s0_data_o[6]), .ZN(n28207) );
  INVX0 U19583 ( .INP(m2s0_data_o[6]), .ZN(n28206) );
  OA22X1 U19584 ( .IN1(n23818), .IN2(n28207), .IN3(n23837), .IN4(n28206), .Q(
        n18274) );
  INVX0 U19585 ( .INP(m5s0_data_o[6]), .ZN(n28205) );
  INVX0 U19586 ( .INP(m7s0_data_o[6]), .ZN(n28209) );
  OA22X1 U19587 ( .IN1(n23832), .IN2(n28205), .IN3(n23824), .IN4(n28209), .Q(
        n18273) );
  INVX0 U19588 ( .INP(m0s0_data_o[6]), .ZN(n28208) );
  INVX0 U19589 ( .INP(m4s0_data_o[6]), .ZN(n28211) );
  OA22X1 U19590 ( .IN1(n23823), .IN2(n28208), .IN3(n23825), .IN4(n28211), .Q(
        n18272) );
  NAND4X0 U19591 ( .IN1(n18275), .IN2(n18274), .IN3(n18273), .IN4(n18272), 
        .QN(s15_data_o[6]) );
  INVX0 U19592 ( .INP(m4s0_data_o[7]), .ZN(n28217) );
  INVX0 U19593 ( .INP(m2s0_data_o[7]), .ZN(n28224) );
  OA22X1 U19594 ( .IN1(n23825), .IN2(n28217), .IN3(n23837), .IN4(n28224), .Q(
        n18279) );
  INVX0 U19595 ( .INP(m0s0_data_o[7]), .ZN(n28220) );
  INVX0 U19596 ( .INP(m5s0_data_o[7]), .ZN(n28223) );
  OA22X1 U19597 ( .IN1(n23823), .IN2(n28220), .IN3(n23832), .IN4(n28223), .Q(
        n18278) );
  INVX0 U19598 ( .INP(m3s0_data_o[7]), .ZN(n28218) );
  INVX0 U19599 ( .INP(m6s0_data_o[7]), .ZN(n28222) );
  OA22X1 U19600 ( .IN1(n23812), .IN2(n28218), .IN3(n23833), .IN4(n28222), .Q(
        n18277) );
  INVX0 U19601 ( .INP(m7s0_data_o[7]), .ZN(n28221) );
  INVX0 U19602 ( .INP(m1s0_data_o[7]), .ZN(n28219) );
  OA22X1 U19603 ( .IN1(n23834), .IN2(n28221), .IN3(n23818), .IN4(n28219), .Q(
        n18276) );
  NAND4X0 U19604 ( .IN1(n18279), .IN2(n18278), .IN3(n18277), .IN4(n18276), 
        .QN(s15_data_o[7]) );
  INVX0 U19605 ( .INP(m6s0_data_o[8]), .ZN(n28233) );
  INVX0 U19606 ( .INP(m2s0_data_o[8]), .ZN(n28231) );
  OA22X1 U19607 ( .IN1(n23799), .IN2(n28233), .IN3(n23837), .IN4(n28231), .Q(
        n18283) );
  INVX0 U19608 ( .INP(m0s0_data_o[8]), .ZN(n28230) );
  INVX0 U19609 ( .INP(m5s0_data_o[8]), .ZN(n28229) );
  OA22X1 U19610 ( .IN1(n23823), .IN2(n28230), .IN3(n23832), .IN4(n28229), .Q(
        n18282) );
  INVX0 U19611 ( .INP(m7s0_data_o[8]), .ZN(n28235) );
  INVX0 U19612 ( .INP(m1s0_data_o[8]), .ZN(n28232) );
  OA22X1 U19613 ( .IN1(n23824), .IN2(n28235), .IN3(n23818), .IN4(n28232), .Q(
        n18281) );
  INVX0 U19614 ( .INP(m4s0_data_o[8]), .ZN(n28236) );
  INVX0 U19615 ( .INP(m3s0_data_o[8]), .ZN(n28234) );
  OA22X1 U19616 ( .IN1(n23836), .IN2(n28236), .IN3(n23835), .IN4(n28234), .Q(
        n18280) );
  NAND4X0 U19617 ( .IN1(n18283), .IN2(n18282), .IN3(n18281), .IN4(n18280), 
        .QN(s15_data_o[8]) );
  INVX0 U19618 ( .INP(m7s0_data_o[9]), .ZN(n28247) );
  INVX0 U19619 ( .INP(m6s0_data_o[9]), .ZN(n28243) );
  OA22X1 U19620 ( .IN1(n23834), .IN2(n28247), .IN3(n23833), .IN4(n28243), .Q(
        n18287) );
  INVX0 U19621 ( .INP(m3s0_data_o[9]), .ZN(n28248) );
  INVX0 U19622 ( .INP(m2s0_data_o[9]), .ZN(n28246) );
  OA22X1 U19623 ( .IN1(n23835), .IN2(n28248), .IN3(n23837), .IN4(n28246), .Q(
        n18286) );
  INVX0 U19624 ( .INP(m4s0_data_o[9]), .ZN(n28241) );
  INVX0 U19625 ( .INP(m5s0_data_o[9]), .ZN(n28245) );
  OA22X1 U19626 ( .IN1(n23825), .IN2(n28241), .IN3(n23832), .IN4(n28245), .Q(
        n18285) );
  INVX0 U19627 ( .INP(m0s0_data_o[9]), .ZN(n28242) );
  INVX0 U19628 ( .INP(m1s0_data_o[9]), .ZN(n28244) );
  OA22X1 U19629 ( .IN1(n23823), .IN2(n28242), .IN3(n23818), .IN4(n28244), .Q(
        n18284) );
  NAND4X0 U19630 ( .IN1(n18287), .IN2(n18286), .IN3(n18285), .IN4(n18284), 
        .QN(s15_data_o[9]) );
  INVX0 U19631 ( .INP(m4s0_data_o[10]), .ZN(n28254) );
  INVX0 U19632 ( .INP(m6s0_data_o[10]), .ZN(n28253) );
  OA22X1 U19633 ( .IN1(n23836), .IN2(n28254), .IN3(n23833), .IN4(n28253), .Q(
        n18291) );
  INVX0 U19634 ( .INP(m7s0_data_o[10]), .ZN(n28259) );
  INVX0 U19635 ( .INP(m1s0_data_o[10]), .ZN(n28257) );
  OA22X1 U19636 ( .IN1(n23824), .IN2(n28259), .IN3(n23818), .IN4(n28257), .Q(
        n18290) );
  INVX0 U19637 ( .INP(m3s0_data_o[10]), .ZN(n28256) );
  INVX0 U19638 ( .INP(m2s0_data_o[10]), .ZN(n28260) );
  OA22X1 U19639 ( .IN1(n23812), .IN2(n28256), .IN3(n23837), .IN4(n28260), .Q(
        n18289) );
  INVX0 U19640 ( .INP(m0s0_data_o[10]), .ZN(n28258) );
  INVX0 U19641 ( .INP(m5s0_data_o[10]), .ZN(n28255) );
  OA22X1 U19642 ( .IN1(n23823), .IN2(n28258), .IN3(n23832), .IN4(n28255), .Q(
        n18288) );
  NAND4X0 U19643 ( .IN1(n18291), .IN2(n18290), .IN3(n18289), .IN4(n18288), 
        .QN(s15_data_o[10]) );
  INVX0 U19644 ( .INP(m5s0_data_o[11]), .ZN(n28270) );
  INVX0 U19645 ( .INP(m3s0_data_o[11]), .ZN(n28271) );
  OA22X1 U19646 ( .IN1(n23826), .IN2(n28270), .IN3(n23835), .IN4(n28271), .Q(
        n18295) );
  INVX0 U19647 ( .INP(m0s0_data_o[11]), .ZN(n28266) );
  INVX0 U19648 ( .INP(m4s0_data_o[11]), .ZN(n28268) );
  OA22X1 U19649 ( .IN1(n23823), .IN2(n28266), .IN3(n23825), .IN4(n28268), .Q(
        n18294) );
  INVX0 U19650 ( .INP(m7s0_data_o[11]), .ZN(n28269) );
  INVX0 U19651 ( .INP(m6s0_data_o[11]), .ZN(n28267) );
  OA22X1 U19652 ( .IN1(n23834), .IN2(n28269), .IN3(n23833), .IN4(n28267), .Q(
        n18293) );
  INVX0 U19653 ( .INP(m1s0_data_o[11]), .ZN(n28272) );
  INVX0 U19654 ( .INP(m2s0_data_o[11]), .ZN(n28265) );
  OA22X1 U19655 ( .IN1(n23818), .IN2(n28272), .IN3(n23837), .IN4(n28265), .Q(
        n18292) );
  NAND4X0 U19656 ( .IN1(n18295), .IN2(n18294), .IN3(n18293), .IN4(n18292), 
        .QN(s15_data_o[11]) );
  INVX0 U19657 ( .INP(m7s0_data_o[12]), .ZN(n28277) );
  INVX0 U19658 ( .INP(m6s0_data_o[12]), .ZN(n28279) );
  OA22X1 U19659 ( .IN1(n23824), .IN2(n28277), .IN3(n23833), .IN4(n28279), .Q(
        n18299) );
  INVX0 U19660 ( .INP(m0s0_data_o[12]), .ZN(n28284) );
  INVX0 U19661 ( .INP(m1s0_data_o[12]), .ZN(n28278) );
  OA22X1 U19662 ( .IN1(n23823), .IN2(n28284), .IN3(n23818), .IN4(n28278), .Q(
        n18298) );
  INVX0 U19663 ( .INP(m5s0_data_o[12]), .ZN(n28281) );
  INVX0 U19664 ( .INP(m3s0_data_o[12]), .ZN(n28282) );
  OA22X1 U19665 ( .IN1(n23832), .IN2(n28281), .IN3(n23835), .IN4(n28282), .Q(
        n18297) );
  INVX0 U19666 ( .INP(m4s0_data_o[12]), .ZN(n28283) );
  INVX0 U19667 ( .INP(m2s0_data_o[12]), .ZN(n28280) );
  OA22X1 U19668 ( .IN1(n23825), .IN2(n28283), .IN3(n23837), .IN4(n28280), .Q(
        n18296) );
  NAND4X0 U19669 ( .IN1(n18299), .IN2(n18298), .IN3(n18297), .IN4(n18296), 
        .QN(s15_data_o[12]) );
  INVX0 U19670 ( .INP(m3s0_data_o[13]), .ZN(n28292) );
  INVX0 U19671 ( .INP(m7s0_data_o[13]), .ZN(n28295) );
  OA22X1 U19672 ( .IN1(n23835), .IN2(n28292), .IN3(n23824), .IN4(n28295), .Q(
        n18303) );
  INVX0 U19673 ( .INP(m5s0_data_o[13]), .ZN(n28293) );
  INVX0 U19674 ( .INP(m6s0_data_o[13]), .ZN(n28291) );
  OA22X1 U19675 ( .IN1(n23826), .IN2(n28293), .IN3(n23833), .IN4(n28291), .Q(
        n18302) );
  INVX0 U19676 ( .INP(m4s0_data_o[13]), .ZN(n28289) );
  INVX0 U19677 ( .INP(m1s0_data_o[13]), .ZN(n28294) );
  OA22X1 U19678 ( .IN1(n23836), .IN2(n28289), .IN3(n23831), .IN4(n28294), .Q(
        n18301) );
  INVX0 U19679 ( .INP(m0s0_data_o[13]), .ZN(n28290) );
  INVX0 U19680 ( .INP(m2s0_data_o[13]), .ZN(n28296) );
  OA22X1 U19681 ( .IN1(n23823), .IN2(n28290), .IN3(n23837), .IN4(n28296), .Q(
        n18300) );
  NAND4X0 U19682 ( .IN1(n18303), .IN2(n18302), .IN3(n18301), .IN4(n18300), 
        .QN(s15_data_o[13]) );
  INVX0 U19683 ( .INP(m3s0_data_o[14]), .ZN(n28305) );
  INVX0 U19684 ( .INP(m2s0_data_o[14]), .ZN(n28308) );
  OA22X1 U19685 ( .IN1(n23812), .IN2(n28305), .IN3(n23837), .IN4(n28308), .Q(
        n18307) );
  INVX0 U19686 ( .INP(m5s0_data_o[14]), .ZN(n28302) );
  INVX0 U19687 ( .INP(m1s0_data_o[14]), .ZN(n28304) );
  OA22X1 U19688 ( .IN1(n23832), .IN2(n28302), .IN3(n23818), .IN4(n28304), .Q(
        n18306) );
  INVX0 U19689 ( .INP(m4s0_data_o[14]), .ZN(n28307) );
  INVX0 U19690 ( .INP(m6s0_data_o[14]), .ZN(n28301) );
  OA22X1 U19691 ( .IN1(n23825), .IN2(n28307), .IN3(n23833), .IN4(n28301), .Q(
        n18305) );
  INVX0 U19692 ( .INP(m0s0_data_o[14]), .ZN(n28306) );
  INVX0 U19693 ( .INP(m7s0_data_o[14]), .ZN(n28303) );
  OA22X1 U19694 ( .IN1(n23823), .IN2(n28306), .IN3(n23824), .IN4(n28303), .Q(
        n18304) );
  NAND4X0 U19695 ( .IN1(n18307), .IN2(n18306), .IN3(n18305), .IN4(n18304), 
        .QN(s15_data_o[14]) );
  INVX0 U19696 ( .INP(m7s0_data_o[15]), .ZN(n28319) );
  INVX0 U19697 ( .INP(m1s0_data_o[15]), .ZN(n28315) );
  OA22X1 U19698 ( .IN1(n23834), .IN2(n28319), .IN3(n23831), .IN4(n28315), .Q(
        n18311) );
  INVX0 U19699 ( .INP(m4s0_data_o[15]), .ZN(n28320) );
  INVX0 U19700 ( .INP(m6s0_data_o[15]), .ZN(n28317) );
  OA22X1 U19701 ( .IN1(n23836), .IN2(n28320), .IN3(n23833), .IN4(n28317), .Q(
        n18310) );
  INVX0 U19702 ( .INP(m5s0_data_o[15]), .ZN(n28318) );
  INVX0 U19703 ( .INP(m2s0_data_o[15]), .ZN(n28314) );
  OA22X1 U19704 ( .IN1(n23832), .IN2(n28318), .IN3(n23837), .IN4(n28314), .Q(
        n18309) );
  INVX0 U19705 ( .INP(m0s0_data_o[15]), .ZN(n28316) );
  INVX0 U19706 ( .INP(m3s0_data_o[15]), .ZN(n28313) );
  OA22X1 U19707 ( .IN1(n23823), .IN2(n28316), .IN3(n23812), .IN4(n28313), .Q(
        n18308) );
  NAND4X0 U19708 ( .IN1(n18311), .IN2(n18310), .IN3(n18309), .IN4(n18308), 
        .QN(s15_data_o[15]) );
  NAND2X0 U19709 ( .IN1(n13825), .IN2(m1s8_cyc), .QN(n18312) );
  NOR2X0 U19710 ( .IN1(n13851), .IN2(n18312), .QN(n18709) );
  NAND2X0 U19711 ( .IN1(\s8/msel/gnt_p1 [0]), .IN2(n18709), .QN(n18712) );
  NOR2X0 U19712 ( .IN1(n18712), .IN2(\s8/msel/gnt_p1 [1]), .QN(n18346) );
  NAND2X0 U19713 ( .IN1(n13773), .IN2(m2s8_cyc), .QN(n18313) );
  NOR2X0 U19714 ( .IN1(n13799), .IN2(n18313), .QN(n18343) );
  NAND2X0 U19715 ( .IN1(n13877), .IN2(m0s8_cyc), .QN(n18314) );
  NOR2X0 U19716 ( .IN1(n13916), .IN2(n18314), .QN(n18701) );
  NOR2X0 U19717 ( .IN1(\s8/msel/gnt_p1 [0]), .IN2(\s8/msel/gnt_p1 [1]), .QN(
        n18327) );
  NAND3X0 U19718 ( .IN1(n13565), .IN2(m6s8_cyc), .IN3(n34631), .QN(n32008) );
  INVX0 U19719 ( .INP(n18343), .ZN(n18706) );
  INVX0 U19720 ( .INP(n18701), .ZN(n18713) );
  NAND2X0 U19721 ( .IN1(n18706), .IN2(n18713), .QN(n18319) );
  NOR2X0 U19722 ( .IN1(n34229), .IN2(n18319), .QN(n18320) );
  INVX0 U19723 ( .INP(n18709), .ZN(n31987) );
  NAND2X0 U19724 ( .IN1(n13489), .IN2(m7s8_cyc), .QN(n18315) );
  NOR2X0 U19725 ( .IN1(n13539), .IN2(n18315), .QN(n31993) );
  INVX0 U19726 ( .INP(n31993), .ZN(n32005) );
  OA21X1 U19727 ( .IN1(n31987), .IN2(n18701), .IN3(n32005), .Q(n18336) );
  INVX0 U19728 ( .INP(n18336), .ZN(n18316) );
  AND3X1 U19729 ( .IN1(n13617), .IN2(m5s8_cyc), .IN3(n34588), .Q(n32009) );
  AO221X1 U19730 ( .IN1(n32008), .IN2(n18320), .IN3(n32008), .IN4(n18316), 
        .IN5(n32009), .Q(n18331) );
  NAND2X0 U19731 ( .IN1(n18327), .IN2(n18331), .QN(n18325) );
  NAND2X0 U19732 ( .IN1(n13721), .IN2(m3s8_cyc), .QN(n18317) );
  NOR2X0 U19733 ( .IN1(n13747), .IN2(n18317), .QN(n18711) );
  INVX0 U19734 ( .INP(n18711), .ZN(n31988) );
  NAND3X0 U19735 ( .IN1(n13669), .IN2(m4s8_cyc), .IN3(n34238), .QN(n18330) );
  NAND2X0 U19736 ( .IN1(n32009), .IN2(n18330), .QN(n18318) );
  NAND2X0 U19737 ( .IN1(n31988), .IN2(n18318), .QN(n18332) );
  AO21X1 U19738 ( .IN1(n18706), .IN2(n18332), .IN3(n18709), .Q(n18326) );
  NAND3X0 U19739 ( .IN1(\s8/msel/gnt_p1 [1]), .IN2(n18326), .IN3(n18713), .QN(
        n18324) );
  OA21X1 U19740 ( .IN1(n31988), .IN2(n18319), .IN3(n18336), .Q(n18322) );
  INVX0 U19741 ( .INP(n18330), .ZN(n32011) );
  INVX0 U19742 ( .INP(n18320), .ZN(n18321) );
  INVX0 U19743 ( .INP(n32008), .ZN(n18347) );
  AO221X1 U19744 ( .IN1(n18322), .IN2(n32011), .IN3(n18322), .IN4(n18321), 
        .IN5(n18347), .Q(n18323) );
  NAND4X0 U19745 ( .IN1(\s8/msel/gnt_p1 [2]), .IN2(n18325), .IN3(n18324), 
        .IN4(n18323), .QN(n18342) );
  INVX0 U19746 ( .INP(n18326), .ZN(n18329) );
  NOR2X0 U19747 ( .IN1(n18347), .IN2(n32011), .QN(n18334) );
  NAND3X0 U19748 ( .IN1(n18334), .IN2(n31993), .IN3(n18706), .QN(n18328) );
  INVX0 U19749 ( .INP(n18327), .ZN(n31998) );
  AO21X1 U19750 ( .IN1(n18329), .IN2(n18328), .IN3(n31998), .Q(n18340) );
  NAND3X0 U19751 ( .IN1(\s8/msel/gnt_p1 [1]), .IN2(n18331), .IN3(n18330), .QN(
        n18339) );
  AND3X1 U19752 ( .IN1(n18713), .IN2(n18334), .IN3(\s8/msel/gnt_p1 [0]), .Q(
        n18333) );
  NOR2X0 U19753 ( .IN1(n18333), .IN2(n18332), .QN(n18337) );
  INVX0 U19754 ( .INP(n18334), .ZN(n18335) );
  NAND2X0 U19755 ( .IN1(\s8/msel/gnt_p1 [0]), .IN2(n34276), .QN(n31992) );
  NAND2X0 U19756 ( .IN1(\s8/msel/gnt_p1 [1]), .IN2(n34229), .QN(n32007) );
  OA21X1 U19757 ( .IN1(n18343), .IN2(n31992), .IN3(n32007), .Q(n18710) );
  AO221X1 U19758 ( .IN1(n18337), .IN2(n18336), .IN3(n18337), .IN4(n18335), 
        .IN5(n18710), .Q(n18338) );
  NAND4X0 U19759 ( .IN1(n34420), .IN2(n18340), .IN3(n18339), .IN4(n18338), 
        .QN(n18341) );
  NAND2X0 U19760 ( .IN1(n18342), .IN2(n18341), .QN(n18348) );
  AO221X1 U19761 ( .IN1(\s8/msel/gnt_p1 [1]), .IN2(n18343), .IN3(n34276), 
        .IN4(n18701), .IN5(n18348), .Q(n18344) );
  NOR2X0 U19762 ( .IN1(n34229), .IN2(n34276), .QN(n32004) );
  NAND2X0 U19763 ( .IN1(n18711), .IN2(n32004), .QN(n18707) );
  NAND2X0 U19764 ( .IN1(n18344), .IN2(n18707), .QN(n18345) );
  NOR2X0 U19765 ( .IN1(n18346), .IN2(n18345), .QN(n18350) );
  MUX21X1 U19766 ( .IN1(n32011), .IN2(n18347), .S(\s8/msel/gnt_p1 [1]), .Q(
        n18703) );
  OA21X1 U19767 ( .IN1(n34420), .IN2(n18703), .IN3(n34229), .Q(n18349) );
  OA22X1 U19768 ( .IN1(\s8/msel/gnt_p1 [2]), .IN2(n18350), .IN3(n18349), .IN4(
        n18348), .Q(n18351) );
  MUX21X1 U19769 ( .IN1(n32009), .IN2(n31993), .S(\s8/msel/gnt_p1 [1]), .Q(
        n18704) );
  NAND3X0 U19770 ( .IN1(\s8/msel/gnt_p1 [0]), .IN2(\s8/msel/gnt_p1 [2]), .IN3(
        n18704), .QN(n18719) );
  NAND2X0 U19771 ( .IN1(n18351), .IN2(n18719), .QN(n17804) );
  NAND3X0 U19772 ( .IN1(n13552), .IN2(m6s7_cyc), .IN3(n34374), .QN(n31710) );
  NAND3X0 U19773 ( .IN1(n13470), .IN2(m7s7_cyc), .IN3(n34347), .QN(n31720) );
  NAND2X0 U19774 ( .IN1(n31710), .IN2(n31720), .QN(n31701) );
  INVX0 U19775 ( .INP(n31701), .ZN(n34129) );
  NOR2X0 U19776 ( .IN1(\s7/msel/gnt_p1 [1]), .IN2(n34129), .QN(n31704) );
  NAND3X0 U19777 ( .IN1(n13812), .IN2(m1s7_cyc), .IN3(n34348), .QN(n31748) );
  NAND3X0 U19778 ( .IN1(n13864), .IN2(m0s7_cyc), .IN3(n34349), .QN(n31750) );
  NAND2X0 U19779 ( .IN1(n31748), .IN2(n31750), .QN(n31696) );
  NAND3X0 U19780 ( .IN1(n13760), .IN2(m2s7_cyc), .IN3(n34363), .QN(n31732) );
  NAND3X0 U19781 ( .IN1(n13708), .IN2(m3s7_cyc), .IN3(n34318), .QN(n31737) );
  NAND2X0 U19782 ( .IN1(n31732), .IN2(n31737), .QN(n31699) );
  NOR2X0 U19783 ( .IN1(n31696), .IN2(n31699), .QN(n34128) );
  NAND3X0 U19784 ( .IN1(n13604), .IN2(m5s7_cyc), .IN3(n34350), .QN(n31734) );
  INVX0 U19785 ( .INP(n31734), .ZN(n31712) );
  NAND2X0 U19786 ( .IN1(\s7/msel/gnt_p1 [1]), .IN2(n31720), .QN(n31697) );
  OA21X1 U19787 ( .IN1(\s7/msel/gnt_p1 [1]), .IN2(n31712), .IN3(n31697), .Q(
        n18363) );
  AND3X1 U19788 ( .IN1(n13656), .IN2(m4s7_cyc), .IN3(n34649), .Q(n31733) );
  INVX0 U19789 ( .INP(n31710), .ZN(n31742) );
  MUX21X1 U19790 ( .IN1(n31733), .IN2(n31742), .S(\s7/msel/gnt_p1 [1]), .Q(
        n31755) );
  OA21X1 U19791 ( .IN1(n18363), .IN2(n31755), .IN3(n34245), .Q(n18352) );
  NOR3X0 U19792 ( .IN1(n31704), .IN2(n34128), .IN3(n18352), .QN(n18362) );
  NAND2X0 U19793 ( .IN1(\s7/msel/gnt_p1 [0]), .IN2(\s7/msel/gnt_p1 [1]), .QN(
        n31729) );
  NOR2X0 U19794 ( .IN1(n31737), .IN2(n31729), .QN(n31752) );
  NOR2X0 U19795 ( .IN1(\s7/msel/gnt_p1 [2]), .IN2(n31752), .QN(n18354) );
  INVX0 U19796 ( .INP(n31732), .ZN(n31727) );
  NOR2X0 U19797 ( .IN1(\s7/msel/gnt_p1 [0]), .IN2(n34439), .QN(n31694) );
  NAND2X0 U19798 ( .IN1(n31727), .IN2(n31694), .QN(n18353) );
  NAND2X0 U19799 ( .IN1(n18354), .IN2(n18353), .QN(n31708) );
  INVX0 U19800 ( .INP(n31729), .ZN(n18358) );
  AND2X1 U19801 ( .IN1(n34439), .IN2(n31748), .Q(n31693) );
  NOR2X0 U19802 ( .IN1(n31693), .IN2(n31694), .QN(n18356) );
  NAND2X0 U19803 ( .IN1(n31737), .IN2(n31732), .QN(n18355) );
  NOR2X0 U19804 ( .IN1(n18356), .IN2(n18355), .QN(n18357) );
  OR2X1 U19805 ( .IN1(\s7/msel/gnt_p1 [0]), .IN2(n31750), .Q(n31709) );
  OA22X1 U19806 ( .IN1(n18358), .IN2(n18357), .IN3(\s7/msel/gnt_p1 [1]), .IN4(
        n31709), .Q(n18360) );
  NOR2X0 U19807 ( .IN1(n31733), .IN2(n31712), .QN(n34130) );
  NAND2X0 U19808 ( .IN1(n34130), .IN2(n34129), .QN(n18359) );
  NAND2X0 U19809 ( .IN1(n18360), .IN2(n18359), .QN(n18361) );
  OA22X1 U19810 ( .IN1(n18362), .IN2(n34424), .IN3(n31708), .IN4(n18361), .Q(
        n18364) );
  NAND3X0 U19811 ( .IN1(\s7/msel/gnt_p1 [0]), .IN2(\s7/msel/gnt_p1 [2]), .IN3(
        n18363), .QN(n31757) );
  NAND2X0 U19812 ( .IN1(n18364), .IN2(n31757), .QN(n17834) );
  NAND3X0 U19813 ( .IN1(m6s12_cyc), .IN2(n34327), .IN3(n34540), .QN(n32976) );
  NAND2X0 U19814 ( .IN1(m7s12_cyc), .IN2(n34643), .QN(n19156) );
  NOR2X0 U19815 ( .IN1(n13535), .IN2(n19156), .QN(n18380) );
  INVX0 U19816 ( .INP(n18380), .ZN(n32978) );
  NAND2X0 U19817 ( .IN1(n32976), .IN2(n32978), .QN(n32952) );
  NAND2X0 U19818 ( .IN1(n34230), .IN2(n32952), .QN(n32958) );
  NAND3X0 U19819 ( .IN1(m2s12_cyc), .IN2(n34329), .IN3(n34541), .QN(n32968) );
  INVX0 U19820 ( .INP(n32968), .ZN(n33005) );
  NAND3X0 U19821 ( .IN1(m3s12_cyc), .IN2(n34330), .IN3(n34507), .QN(n32980) );
  INVX0 U19822 ( .INP(n32980), .ZN(n32965) );
  NOR2X0 U19823 ( .IN1(n33005), .IN2(n32965), .QN(n34183) );
  NAND3X0 U19824 ( .IN1(m0s12_cyc), .IN2(n34354), .IN3(n34509), .QN(n32969) );
  NAND3X0 U19825 ( .IN1(m1s12_cyc), .IN2(n34355), .IN3(n34508), .QN(n33003) );
  NAND2X0 U19826 ( .IN1(n32969), .IN2(n33003), .QN(n18373) );
  NAND3X0 U19827 ( .IN1(m5s12_cyc), .IN2(n34328), .IN3(n34506), .QN(n32979) );
  INVX0 U19828 ( .INP(n32979), .ZN(n18381) );
  AO221X1 U19829 ( .IN1(n32958), .IN2(n34183), .IN3(n32958), .IN4(n18373), 
        .IN5(n18381), .Q(n18368) );
  NAND2X0 U19830 ( .IN1(\s12/msel/gnt_p3 [1]), .IN2(n34269), .QN(n32983) );
  OR2X1 U19831 ( .IN1(n32978), .IN2(n32983), .Q(n18367) );
  NAND2X0 U19832 ( .IN1(n34269), .IN2(n34230), .QN(n32988) );
  NAND2X0 U19833 ( .IN1(m4s12_cyc), .IN2(n34642), .QN(n19157) );
  NOR2X0 U19834 ( .IN1(n13691), .IN2(n19157), .QN(n32962) );
  INVX0 U19835 ( .INP(n32962), .ZN(n32994) );
  NAND3X0 U19836 ( .IN1(\s12/msel/gnt_p3 [1]), .IN2(n32994), .IN3(n32979), 
        .QN(n18365) );
  NAND2X0 U19837 ( .IN1(n34183), .IN2(n18365), .QN(n18369) );
  NAND4X0 U19838 ( .IN1(n32969), .IN2(n33003), .IN3(n32988), .IN4(n18369), 
        .QN(n18366) );
  NAND4X0 U19839 ( .IN1(\s12/msel/gnt_p3 [2]), .IN2(n18368), .IN3(n18367), 
        .IN4(n18366), .QN(n18378) );
  NAND3X0 U19840 ( .IN1(n32994), .IN2(n32979), .IN3(n32952), .QN(n18372) );
  INVX0 U19841 ( .INP(n18369), .ZN(n18371) );
  INVX0 U19842 ( .INP(n32988), .ZN(n18370) );
  INVX0 U19843 ( .INP(n33003), .ZN(n32967) );
  AO222X1 U19844 ( .IN1(n18372), .IN2(n18371), .IN3(n18372), .IN4(n32988), 
        .IN5(n18370), .IN6(n32967), .Q(n18376) );
  INVX0 U19845 ( .INP(n18373), .ZN(n34184) );
  NAND4X0 U19846 ( .IN1(\s12/msel/gnt_p3 [1]), .IN2(n34184), .IN3(n32979), 
        .IN4(n32994), .QN(n18375) );
  NAND2X0 U19847 ( .IN1(n34230), .IN2(\s12/msel/gnt_p3 [0]), .QN(n33002) );
  AO21X1 U19848 ( .IN1(n32983), .IN2(n33002), .IN3(n34183), .Q(n18374) );
  NAND4X0 U19849 ( .IN1(n18376), .IN2(n34450), .IN3(n18375), .IN4(n18374), 
        .QN(n18377) );
  NAND2X0 U19850 ( .IN1(n18378), .IN2(n18377), .QN(n18382) );
  INVX0 U19851 ( .INP(n32969), .ZN(n33004) );
  MUX21X1 U19852 ( .IN1(n33004), .IN2(n32967), .S(\s12/msel/gnt_p3 [0]), .Q(
        n32949) );
  NOR2X0 U19853 ( .IN1(n34269), .IN2(n34230), .QN(n32948) );
  NAND2X0 U19854 ( .IN1(n32965), .IN2(n32948), .QN(n33007) );
  OA21X1 U19855 ( .IN1(n18382), .IN2(n32949), .IN3(n33007), .Q(n18379) );
  OA22X1 U19856 ( .IN1(\s12/msel/gnt_p3 [2]), .IN2(n18379), .IN3(n34230), 
        .IN4(n18382), .Q(n18386) );
  NAND2X0 U19857 ( .IN1(\s12/msel/gnt_p3 [1]), .IN2(n18380), .QN(n32956) );
  OA21X1 U19858 ( .IN1(n18381), .IN2(n18382), .IN3(n32956), .Q(n18384) );
  OA22X1 U19859 ( .IN1(n32962), .IN2(n18382), .IN3(n34230), .IN4(n32976), .Q(
        n18383) );
  AO221X1 U19860 ( .IN1(\s12/msel/gnt_p3 [0]), .IN2(n18384), .IN3(n34269), 
        .IN4(n18383), .IN5(n34450), .Q(n18385) );
  NAND2X0 U19861 ( .IN1(n18386), .IN2(n18385), .QN(n17696) );
  NAND3X0 U19862 ( .IN1(m3s7_cyc), .IN2(n34318), .IN3(n34498), .QN(n31644) );
  NAND2X0 U19863 ( .IN1(\s7/msel/gnt_p3 [0]), .IN2(\s7/msel/gnt_p3 [1]), .QN(
        n31671) );
  NAND2X0 U19864 ( .IN1(m6s7_cyc), .IN2(n34567), .QN(n18387) );
  NOR2X0 U19865 ( .IN1(n13578), .IN2(n18387), .QN(n31643) );
  INVX0 U19866 ( .INP(n31643), .ZN(n31676) );
  NAND3X0 U19867 ( .IN1(m7s7_cyc), .IN2(n34347), .IN3(n34499), .QN(n31657) );
  NAND2X0 U19868 ( .IN1(n31676), .IN2(n31657), .QN(n31635) );
  INVX0 U19869 ( .INP(n31635), .ZN(n18394) );
  NAND3X0 U19870 ( .IN1(m2s7_cyc), .IN2(n34363), .IN3(n34600), .QN(n31680) );
  NAND3X0 U19871 ( .IN1(m0s7_cyc), .IN2(n34349), .IN3(n34497), .QN(n31681) );
  NAND3X0 U19872 ( .IN1(m1s7_cyc), .IN2(n34348), .IN3(n34533), .QN(n31658) );
  NAND2X0 U19873 ( .IN1(n31681), .IN2(n31658), .QN(n18398) );
  NAND3X0 U19874 ( .IN1(m5s7_cyc), .IN2(n34350), .IN3(n34534), .QN(n31642) );
  NAND2X0 U19875 ( .IN1(n34410), .IN2(n31642), .QN(n31669) );
  AO221X1 U19876 ( .IN1(n18394), .IN2(n31680), .IN3(n18394), .IN4(n18398), 
        .IN5(n31669), .Q(n18393) );
  NAND2X0 U19877 ( .IN1(m4s7_cyc), .IN2(n34594), .QN(n18388) );
  NOR2X0 U19878 ( .IN1(n13682), .IN2(n18388), .QN(n31645) );
  INVX0 U19879 ( .INP(n31645), .ZN(n31670) );
  NAND2X0 U19880 ( .IN1(n31670), .IN2(n31642), .QN(n31630) );
  NOR2X0 U19881 ( .IN1(n34262), .IN2(n31630), .QN(n18389) );
  NAND2X0 U19882 ( .IN1(n31680), .IN2(n31644), .QN(n31629) );
  NOR2X0 U19883 ( .IN1(n18389), .IN2(n31629), .QN(n18396) );
  AND2X1 U19884 ( .IN1(n31644), .IN2(n18396), .Q(n18391) );
  NAND2X0 U19885 ( .IN1(\s7/msel/gnt_p3 [1]), .IN2(n34410), .QN(n31652) );
  NAND2X0 U19886 ( .IN1(\s7/msel/gnt_p3 [0]), .IN2(n34262), .QN(n31648) );
  NAND2X0 U19887 ( .IN1(n31652), .IN2(n31648), .QN(n18399) );
  INVX0 U19888 ( .INP(n18399), .ZN(n18390) );
  OA22X1 U19889 ( .IN1(n18391), .IN2(n18398), .IN3(n18394), .IN4(n18390), .Q(
        n18392) );
  NAND3X0 U19890 ( .IN1(n18393), .IN2(n18392), .IN3(\s7/msel/gnt_p3 [2]), .QN(
        n18404) );
  OR2X1 U19891 ( .IN1(n31630), .IN2(n18394), .Q(n18397) );
  NAND2X0 U19892 ( .IN1(n34410), .IN2(n34262), .QN(n31655) );
  INVX0 U19893 ( .INP(n31655), .ZN(n18395) );
  INVX0 U19894 ( .INP(n31658), .ZN(n31683) );
  AO222X1 U19895 ( .IN1(n18397), .IN2(n18396), .IN3(n18397), .IN4(n31655), 
        .IN5(n18395), .IN6(n31683), .Q(n18402) );
  INVX0 U19896 ( .INP(n18398), .ZN(n21783) );
  NAND4X0 U19897 ( .IN1(\s7/msel/gnt_p3 [1]), .IN2(n21783), .IN3(n31642), 
        .IN4(n31670), .QN(n18401) );
  NAND2X0 U19898 ( .IN1(n31629), .IN2(n18399), .QN(n18400) );
  NAND4X0 U19899 ( .IN1(n18402), .IN2(n34380), .IN3(n18401), .IN4(n18400), 
        .QN(n18403) );
  NAND2X0 U19900 ( .IN1(n18404), .IN2(n18403), .QN(n18407) );
  INVX0 U19901 ( .INP(n31681), .ZN(n31673) );
  MUX21X1 U19902 ( .IN1(n31673), .IN2(n31683), .S(\s7/msel/gnt_p3 [0]), .Q(
        n31633) );
  OA22X1 U19903 ( .IN1(n31644), .IN2(n31671), .IN3(n18407), .IN4(n31633), .Q(
        n18405) );
  OA22X1 U19904 ( .IN1(\s7/msel/gnt_p3 [2]), .IN2(n18405), .IN3(n18407), .IN4(
        n34262), .Q(n18412) );
  INVX0 U19905 ( .INP(n31642), .ZN(n31661) );
  OR2X1 U19906 ( .IN1(n34262), .IN2(n31657), .Q(n31634) );
  OA21X1 U19907 ( .IN1(n31661), .IN2(n18407), .IN3(n31634), .Q(n18406) );
  NOR2X0 U19908 ( .IN1(n18406), .IN2(n34380), .QN(n18410) );
  OR2X1 U19909 ( .IN1(n18407), .IN2(n31645), .Q(n18408) );
  NAND2X0 U19910 ( .IN1(n34410), .IN2(n18408), .QN(n18409) );
  NAND2X0 U19911 ( .IN1(n18410), .IN2(n18409), .QN(n18411) );
  NAND2X0 U19912 ( .IN1(n18412), .IN2(n18411), .QN(n17836) );
  NAND3X0 U19913 ( .IN1(n13619), .IN2(m5s10_cyc), .IN3(n34323), .QN(n32581) );
  INVX0 U19914 ( .INP(n32581), .ZN(n18414) );
  NAND3X0 U19915 ( .IN1(n13494), .IN2(m7s10_cyc), .IN3(n34353), .QN(n32577) );
  NAND2X0 U19916 ( .IN1(\s10/msel/gnt_p1 [1]), .IN2(n32577), .QN(n32591) );
  OA21X1 U19917 ( .IN1(\s10/msel/gnt_p1 [1]), .IN2(n18414), .IN3(n32591), .Q(
        n32560) );
  NAND3X0 U19918 ( .IN1(\s10/msel/gnt_p1 [0]), .IN2(n32560), .IN3(
        \s10/msel/gnt_p1 [2]), .QN(n18435) );
  NAND3X0 U19919 ( .IN1(n13671), .IN2(m4s10_cyc), .IN3(n34620), .QN(n32583) );
  NAND3X0 U19920 ( .IN1(n13567), .IN2(m6s10_cyc), .IN3(n34632), .QN(n32578) );
  OA221X1 U19921 ( .IN1(\s10/msel/gnt_p1 [1]), .IN2(n32583), .IN3(n34253), 
        .IN4(n32578), .IN5(\s10/msel/gnt_p1 [2]), .Q(n18413) );
  NOR2X0 U19922 ( .IN1(\s10/msel/gnt_p1 [0]), .IN2(n18413), .QN(n32574) );
  NAND3X0 U19923 ( .IN1(n13775), .IN2(m2s10_cyc), .IN3(n34322), .QN(n32576) );
  INVX0 U19924 ( .INP(n32576), .ZN(n32567) );
  NAND3X0 U19925 ( .IN1(n13723), .IN2(m3s10_cyc), .IN3(n34606), .QN(n32586) );
  NAND2X0 U19926 ( .IN1(n18414), .IN2(n32583), .QN(n18415) );
  AND2X1 U19927 ( .IN1(n32586), .IN2(n18415), .Q(n18423) );
  NAND3X0 U19928 ( .IN1(n13827), .IN2(m1s10_cyc), .IN3(n34638), .QN(n32565) );
  OAI21X1 U19929 ( .IN1(n32567), .IN2(n18423), .IN3(n32565), .QN(n18425) );
  NAND3X0 U19930 ( .IN1(n13879), .IN2(m0s10_cyc), .IN3(n34619), .QN(n32566) );
  NAND3X0 U19931 ( .IN1(\s10/msel/gnt_p1 [1]), .IN2(n18425), .IN3(n32566), 
        .QN(n18420) );
  INVX0 U19932 ( .INP(n32578), .ZN(n32598) );
  INVX0 U19933 ( .INP(n32566), .ZN(n18431) );
  OA21X1 U19934 ( .IN1(n18431), .IN2(n32565), .IN3(n32577), .Q(n18421) );
  OA21X1 U19935 ( .IN1(n32598), .IN2(n18421), .IN3(n32581), .Q(n18424) );
  NAND2X0 U19936 ( .IN1(n32566), .IN2(n32576), .QN(n18417) );
  NAND2X0 U19937 ( .IN1(\s10/msel/gnt_p1 [0]), .IN2(n32583), .QN(n18416) );
  OA221X1 U19938 ( .IN1(n18417), .IN2(n32586), .IN3(n18417), .IN4(n18416), 
        .IN5(n18421), .Q(n18418) );
  OA22X1 U19939 ( .IN1(\s10/msel/gnt_p1 [1]), .IN2(n18424), .IN3(n32598), 
        .IN4(n18418), .Q(n18419) );
  NAND3X0 U19940 ( .IN1(\s10/msel/gnt_p1 [2]), .IN2(n18420), .IN3(n18419), 
        .QN(n18430) );
  INVX0 U19941 ( .INP(n32583), .ZN(n32595) );
  AO221X1 U19942 ( .IN1(n18421), .IN2(n18431), .IN3(n18421), .IN4(n34434), 
        .IN5(n32595), .Q(n18422) );
  AO221X1 U19943 ( .IN1(n18423), .IN2(n32598), .IN3(n18423), .IN4(n18422), 
        .IN5(n32567), .Q(n18428) );
  OR4X1 U19944 ( .IN1(n34253), .IN2(n34434), .IN3(n32595), .IN4(n18424), .Q(
        n18427) );
  NAND2X0 U19945 ( .IN1(n34253), .IN2(n18425), .QN(n18426) );
  NAND4X0 U19946 ( .IN1(n34610), .IN2(n18428), .IN3(n18427), .IN4(n18426), 
        .QN(n18429) );
  NAND2X0 U19947 ( .IN1(n18430), .IN2(n18429), .QN(n18433) );
  INVX0 U19948 ( .INP(n32586), .ZN(n21772) );
  NOR2X0 U19949 ( .IN1(n34434), .IN2(n34253), .QN(n32564) );
  NAND2X0 U19950 ( .IN1(n21772), .IN2(n32564), .QN(n32568) );
  OA221X1 U19951 ( .IN1(n18433), .IN2(n18431), .IN3(n18433), .IN4(n34253), 
        .IN5(n32568), .Q(n18432) );
  OA22X1 U19952 ( .IN1(n32574), .IN2(n18433), .IN3(\s10/msel/gnt_p1 [2]), 
        .IN4(n18432), .Q(n18434) );
  NAND2X0 U19953 ( .IN1(n18435), .IN2(n18434), .QN(n17748) );
  NAND3X0 U19954 ( .IN1(n13670), .IN2(m4s9_cyc), .IN3(n34319), .QN(n32242) );
  INVX0 U19955 ( .INP(n32242), .ZN(n32269) );
  NAND3X0 U19956 ( .IN1(n13566), .IN2(m6s9_cyc), .IN3(n34320), .QN(n32265) );
  INVX0 U19957 ( .INP(n32265), .ZN(n32233) );
  MUX21X1 U19958 ( .IN1(n32269), .IN2(n32233), .S(\s9/msel/gnt_p1 [1]), .Q(
        n32231) );
  OA21X1 U19959 ( .IN1(n34442), .IN2(n32231), .IN3(n34260), .Q(n18456) );
  NAND3X0 U19960 ( .IN1(n13774), .IN2(m2s9_cyc), .IN3(n34352), .QN(n32237) );
  INVX0 U19961 ( .INP(n32237), .ZN(n18443) );
  NAND3X0 U19962 ( .IN1(n13618), .IN2(m5s9_cyc), .IN3(n34351), .QN(n32241) );
  NAND3X0 U19963 ( .IN1(n13722), .IN2(m3s9_cyc), .IN3(n34636), .QN(n32250) );
  OA21X1 U19964 ( .IN1(n32269), .IN2(n32241), .IN3(n32250), .Q(n18441) );
  NAND3X0 U19965 ( .IN1(n13826), .IN2(m1s9_cyc), .IN3(n34618), .QN(n32239) );
  OA21X1 U19966 ( .IN1(n18443), .IN2(n18441), .IN3(n32239), .Q(n18445) );
  NAND3X0 U19967 ( .IN1(n13878), .IN2(m0s9_cyc), .IN3(n34321), .QN(n32238) );
  INVX0 U19968 ( .INP(n32238), .ZN(n18446) );
  NAND3X0 U19969 ( .IN1(n13490), .IN2(m7s9_cyc), .IN3(n34364), .QN(n18457) );
  OA21X1 U19970 ( .IN1(n32239), .IN2(n18446), .IN3(n18457), .Q(n18444) );
  AO221X1 U19971 ( .IN1(n18444), .IN2(n18446), .IN3(n18444), .IN4(n34260), 
        .IN5(n32269), .Q(n18436) );
  OA21X1 U19972 ( .IN1(n32233), .IN2(n18436), .IN3(n18441), .Q(n18437) );
  OA22X1 U19973 ( .IN1(\s9/msel/gnt_p1 [1]), .IN2(n18445), .IN3(n18443), .IN4(
        n18437), .Q(n18439) );
  OAI21X1 U19974 ( .IN1(n32233), .IN2(n18444), .IN3(n32241), .QN(n18440) );
  NAND4X0 U19975 ( .IN1(\s9/msel/gnt_p1 [1]), .IN2(\s9/msel/gnt_p1 [0]), .IN3(
        n32242), .IN4(n18440), .QN(n18438) );
  NAND3X0 U19976 ( .IN1(n34442), .IN2(n18439), .IN3(n18438), .QN(n18451) );
  NAND2X0 U19977 ( .IN1(n34400), .IN2(n18440), .QN(n18449) );
  AO221X1 U19978 ( .IN1(n18441), .IN2(n32269), .IN3(n18441), .IN4(n34260), 
        .IN5(n18446), .Q(n18442) );
  AO221X1 U19979 ( .IN1(n18444), .IN2(n18443), .IN3(n18444), .IN4(n18442), 
        .IN5(n32233), .Q(n18448) );
  OR3X1 U19980 ( .IN1(n34400), .IN2(n18446), .IN3(n18445), .Q(n18447) );
  NAND4X0 U19981 ( .IN1(\s9/msel/gnt_p1 [2]), .IN2(n18449), .IN3(n18448), 
        .IN4(n18447), .QN(n18450) );
  NAND2X0 U19982 ( .IN1(n18451), .IN2(n18450), .QN(n18455) );
  NOR2X0 U19983 ( .IN1(\s9/msel/gnt_p1 [1]), .IN2(n32238), .QN(n18453) );
  NAND2X0 U19984 ( .IN1(\s9/msel/gnt_p1 [0]), .IN2(\s9/msel/gnt_p1 [1]), .QN(
        n18452) );
  OA22X1 U19985 ( .IN1(n18453), .IN2(n18455), .IN3(n32250), .IN4(n18452), .Q(
        n18454) );
  OA22X1 U19986 ( .IN1(n18456), .IN2(n18455), .IN3(\s9/msel/gnt_p1 [2]), .IN4(
        n18454), .Q(n18459) );
  INVX0 U19987 ( .INP(n18457), .ZN(n32232) );
  NOR2X0 U19988 ( .IN1(n32232), .IN2(n34400), .QN(n32256) );
  INVX0 U19989 ( .INP(n32241), .ZN(n32268) );
  NOR2X0 U19990 ( .IN1(\s9/msel/gnt_p1 [1]), .IN2(n32268), .QN(n32234) );
  OR4X1 U19991 ( .IN1(n32256), .IN2(n32234), .IN3(n34442), .IN4(n34260), .Q(
        n18458) );
  NAND2X0 U19992 ( .IN1(n18459), .IN2(n18458), .QN(n17776) );
  AND3X1 U19993 ( .IN1(n13641), .IN2(n13615), .IN3(m5s14_cyc), .Q(n33684) );
  NAND3X0 U19994 ( .IN1(n13537), .IN2(n13484), .IN3(m7s14_cyc), .QN(n33676) );
  INVX0 U19995 ( .INP(n33676), .ZN(n33667) );
  OA221X1 U19996 ( .IN1(\s14/msel/gnt_p0 [1]), .IN2(n33684), .IN3(n34247), 
        .IN4(n33667), .IN5(\s14/msel/gnt_p0 [2]), .Q(n33696) );
  NAND3X0 U19997 ( .IN1(n13745), .IN2(n13719), .IN3(m3s14_cyc), .QN(n18461) );
  INVX0 U19998 ( .INP(n18461), .ZN(n33668) );
  NAND3X0 U19999 ( .IN1(n13849), .IN2(n13823), .IN3(m1s14_cyc), .QN(n33672) );
  NAND3X0 U20000 ( .IN1(n13797), .IN2(n13771), .IN3(m2s14_cyc), .QN(n33669) );
  INVX0 U20001 ( .INP(n33669), .ZN(n33682) );
  NOR2X0 U20002 ( .IN1(n33668), .IN2(n33682), .QN(n33654) );
  NAND2X0 U20003 ( .IN1(n33672), .IN2(n33654), .QN(n18460) );
  OA21X1 U20004 ( .IN1(n33668), .IN2(n34247), .IN3(n18460), .Q(n18467) );
  NAND2X0 U20005 ( .IN1(\s14/msel/gnt_p0 [0]), .IN2(\s14/msel/gnt_p0 [1]), 
        .QN(n33673) );
  NOR2X0 U20006 ( .IN1(n18461), .IN2(n33673), .QN(n33700) );
  NOR2X0 U20007 ( .IN1(\s14/msel/gnt_p0 [2]), .IN2(n33700), .QN(n18463) );
  NOR2X0 U20008 ( .IN1(\s14/msel/gnt_p0 [0]), .IN2(n34247), .QN(n33659) );
  NAND2X0 U20009 ( .IN1(n33682), .IN2(n33659), .QN(n18462) );
  NAND2X0 U20010 ( .IN1(n18463), .IN2(n18462), .QN(n33663) );
  NAND3X0 U20011 ( .IN1(n13693), .IN2(n13667), .IN3(m4s14_cyc), .QN(n33688) );
  INVX0 U20012 ( .INP(n33688), .ZN(n18469) );
  NOR2X0 U20013 ( .IN1(n18469), .IN2(n33684), .QN(n33643) );
  NAND3X0 U20014 ( .IN1(n13589), .IN2(n13563), .IN3(m6s14_cyc), .QN(n33686) );
  NAND2X0 U20015 ( .IN1(n33686), .IN2(n33676), .QN(n33644) );
  INVX0 U20016 ( .INP(n33644), .ZN(n18465) );
  NAND3X0 U20017 ( .IN1(n13912), .IN2(n13875), .IN3(m0s14_cyc), .QN(n33694) );
  NOR2X0 U20018 ( .IN1(\s14/msel/gnt_p0 [0]), .IN2(n33694), .QN(n18464) );
  AO22X1 U20019 ( .IN1(n33643), .IN2(n18465), .IN3(n18464), .IN4(n34247), .Q(
        n18466) );
  NOR3X0 U20020 ( .IN1(n18467), .IN2(n33663), .IN3(n18466), .QN(n18468) );
  NOR2X0 U20021 ( .IN1(n33696), .IN2(n18468), .QN(n18472) );
  INVX0 U20022 ( .INP(n33686), .ZN(n33660) );
  MUX21X1 U20023 ( .IN1(n18469), .IN2(n33660), .S(\s14/msel/gnt_p0 [1]), .Q(
        n33695) );
  AND2X1 U20024 ( .IN1(n33694), .IN2(n33672), .Q(n33649) );
  AO222X1 U20025 ( .IN1(n34639), .IN2(n33695), .IN3(n34247), .IN4(n33644), 
        .IN5(n33649), .IN6(n33654), .Q(n18470) );
  NAND2X0 U20026 ( .IN1(\s14/msel/gnt_p0 [2]), .IN2(n18470), .QN(n18471) );
  NAND2X0 U20027 ( .IN1(n18472), .IN2(n18471), .QN(n17635) );
  NOR2X0 U20028 ( .IN1(n34280), .IN2(n34428), .QN(n29801) );
  NAND3X0 U20029 ( .IN1(m2s1_cyc), .IN2(n34297), .IN3(n34558), .QN(n29789) );
  NAND2X0 U20030 ( .IN1(\s1/msel/gnt_p3 [1]), .IN2(n34280), .QN(n29734) );
  NAND3X0 U20031 ( .IN1(m7s1_cyc), .IN2(n34296), .IN3(n34559), .QN(n29758) );
  OA21X1 U20032 ( .IN1(n29758), .IN2(n29734), .IN3(\s1/msel/gnt_p3 [2]), .Q(
        n18477) );
  NAND3X0 U20033 ( .IN1(m5s1_cyc), .IN2(n34295), .IN3(n34556), .QN(n29750) );
  INVX0 U20034 ( .INP(n29750), .ZN(n29754) );
  NOR2X0 U20035 ( .IN1(\s1/msel/gnt_p3 [0]), .IN2(\s1/msel/gnt_p3 [1]), .QN(
        n29763) );
  INVX0 U20036 ( .INP(n29789), .ZN(n29773) );
  NAND3X0 U20037 ( .IN1(m3s1_cyc), .IN2(n34335), .IN3(n34521), .QN(n29749) );
  INVX0 U20038 ( .INP(n29749), .ZN(n29791) );
  NOR2X0 U20039 ( .IN1(n29773), .IN2(n29791), .QN(n18481) );
  NAND2X0 U20040 ( .IN1(\s1/msel/gnt_p3 [0]), .IN2(\s1/msel/gnt_p3 [1]), .QN(
        n29752) );
  INVX0 U20041 ( .INP(n29752), .ZN(n29777) );
  NAND3X0 U20042 ( .IN1(m4s1_cyc), .IN2(n34336), .IN3(n34483), .QN(n29776) );
  INVX0 U20043 ( .INP(n29776), .ZN(n29765) );
  NOR2X0 U20044 ( .IN1(n29765), .IN2(n29754), .QN(n18480) );
  NAND2X0 U20045 ( .IN1(n29777), .IN2(n18480), .QN(n18473) );
  AO22X1 U20046 ( .IN1(n29754), .IN2(n29763), .IN3(n18481), .IN4(n18473), .Q(
        n18474) );
  INVX0 U20047 ( .INP(n18480), .ZN(n29732) );
  NAND3X0 U20048 ( .IN1(m0s1_cyc), .IN2(n34294), .IN3(n34557), .QN(n29790) );
  NAND3X0 U20049 ( .IN1(m1s1_cyc), .IN2(n34293), .IN3(n34555), .QN(n29751) );
  NAND2X0 U20050 ( .IN1(n29790), .IN2(n29751), .QN(n29742) );
  AO221X1 U20051 ( .IN1(n18474), .IN2(n29732), .IN3(n18474), .IN4(n29734), 
        .IN5(n29742), .Q(n18476) );
  NAND3X0 U20052 ( .IN1(m6s1_cyc), .IN2(n34306), .IN3(n34522), .QN(n29756) );
  NAND2X0 U20053 ( .IN1(n29758), .IN2(n29756), .QN(n29731) );
  NAND3X0 U20054 ( .IN1(n29750), .IN2(n29731), .IN3(n34427), .QN(n18475) );
  NAND3X0 U20055 ( .IN1(n18477), .IN2(n18476), .IN3(n18475), .QN(n18486) );
  NOR2X0 U20056 ( .IN1(\s1/msel/gnt_p3 [1]), .IN2(n34280), .QN(n29733) );
  INVX0 U20057 ( .INP(n18481), .ZN(n29741) );
  INVX0 U20058 ( .INP(n29758), .ZN(n29771) );
  INVX0 U20059 ( .INP(n29763), .ZN(n29772) );
  INVX0 U20060 ( .INP(n29742), .ZN(n18478) );
  AO222X1 U20061 ( .IN1(n29751), .IN2(n29771), .IN3(n29772), .IN4(n29731), 
        .IN5(n18478), .IN6(\s1/msel/gnt_p3 [1]), .Q(n18479) );
  AOI22X1 U20062 ( .IN1(n29733), .IN2(n29741), .IN3(n18480), .IN4(n18479), 
        .QN(n18484) );
  NAND2X0 U20063 ( .IN1(n29763), .IN2(n29751), .QN(n29736) );
  AO221X1 U20064 ( .IN1(n18481), .IN2(n29732), .IN3(n18481), .IN4(n29756), 
        .IN5(n29736), .Q(n18483) );
  INVX0 U20065 ( .INP(n29734), .ZN(n29768) );
  NAND2X0 U20066 ( .IN1(n29791), .IN2(n29768), .QN(n18482) );
  NAND4X0 U20067 ( .IN1(n18484), .IN2(n34428), .IN3(n18483), .IN4(n18482), 
        .QN(n18485) );
  NAND2X0 U20068 ( .IN1(n18486), .IN2(n18485), .QN(n18491) );
  INVX0 U20069 ( .INP(n29790), .ZN(n29753) );
  INVX0 U20070 ( .INP(n29751), .ZN(n29792) );
  MUX21X1 U20071 ( .IN1(n29753), .IN2(n29792), .S(\s1/msel/gnt_p3 [0]), .Q(
        n29737) );
  OA22X1 U20072 ( .IN1(n29789), .IN2(n29734), .IN3(n18491), .IN4(n29737), .Q(
        n18488) );
  NAND2X0 U20073 ( .IN1(n29791), .IN2(n29777), .QN(n18487) );
  AND3X1 U20074 ( .IN1(n18488), .IN2(n34428), .IN3(n18487), .Q(n18490) );
  OA21X1 U20075 ( .IN1(n34427), .IN2(n29756), .IN3(\s1/msel/gnt_p3 [2]), .Q(
        n29793) );
  OA21X1 U20076 ( .IN1(n29765), .IN2(n18491), .IN3(n29793), .Q(n18489) );
  NOR3X0 U20077 ( .IN1(n29801), .IN2(n18490), .IN3(n18489), .QN(n18493) );
  NOR2X0 U20078 ( .IN1(n34427), .IN2(n29758), .QN(n29800) );
  INVX0 U20079 ( .INP(n18491), .ZN(n18494) );
  OA221X1 U20080 ( .IN1(n29800), .IN2(n18494), .IN3(n29800), .IN4(n29750), 
        .IN5(n29801), .Q(n18492) );
  NOR2X0 U20081 ( .IN1(n18493), .IN2(n18492), .QN(n18496) );
  NAND2X0 U20082 ( .IN1(n18494), .IN2(\s1/msel/gnt_p3 [1]), .QN(n18495) );
  NAND2X0 U20083 ( .IN1(n18496), .IN2(n18495), .QN(n18004) );
  NAND3X0 U20084 ( .IN1(n13601), .IN2(m5s4_cyc), .IN3(n34313), .QN(n30754) );
  INVX0 U20085 ( .INP(n30754), .ZN(n18497) );
  NAND3X0 U20086 ( .IN1(n13464), .IN2(m7s4_cyc), .IN3(n34314), .QN(n30752) );
  NAND2X0 U20087 ( .IN1(\s4/msel/gnt_p1 [1]), .IN2(n30752), .QN(n30729) );
  OA21X1 U20088 ( .IN1(\s4/msel/gnt_p1 [1]), .IN2(n18497), .IN3(n30729), .Q(
        n18508) );
  NAND3X0 U20089 ( .IN1(n13653), .IN2(m4s4_cyc), .IN3(n34338), .QN(n30725) );
  INVX0 U20090 ( .INP(n30725), .ZN(n30762) );
  NAND3X0 U20091 ( .IN1(n13549), .IN2(m6s4_cyc), .IN3(n34339), .QN(n30742) );
  INVX0 U20092 ( .INP(n30742), .ZN(n30766) );
  MUX21X1 U20093 ( .IN1(n30762), .IN2(n30766), .S(\s4/msel/gnt_p1 [1]), .Q(
        n30781) );
  NOR2X0 U20094 ( .IN1(n18508), .IN2(n30781), .QN(n18498) );
  NOR2X0 U20095 ( .IN1(n18498), .IN2(\s4/msel/gnt_p1 [0]), .QN(n18500) );
  NAND2X0 U20096 ( .IN1(n30742), .IN2(n30752), .QN(n30723) );
  NAND2X0 U20097 ( .IN1(n34389), .IN2(n30723), .QN(n30733) );
  NAND3X0 U20098 ( .IN1(n13861), .IN2(m0s4_cyc), .IN3(n34340), .QN(n30751) );
  INVX0 U20099 ( .INP(n30751), .ZN(n30777) );
  NAND3X0 U20100 ( .IN1(n13809), .IN2(m1s4_cyc), .IN3(n34315), .QN(n30753) );
  INVX0 U20101 ( .INP(n30753), .ZN(n18502) );
  NOR2X0 U20102 ( .IN1(n30777), .IN2(n18502), .QN(n30724) );
  NAND3X0 U20103 ( .IN1(n13757), .IN2(m2s4_cyc), .IN3(n34627), .QN(n30750) );
  INVX0 U20104 ( .INP(n30750), .ZN(n30764) );
  NAND3X0 U20105 ( .IN1(n13705), .IN2(m3s4_cyc), .IN3(n34617), .QN(n30749) );
  INVX0 U20106 ( .INP(n30749), .ZN(n30717) );
  NOR2X0 U20107 ( .IN1(n30764), .IN2(n30717), .QN(n30721) );
  NAND2X0 U20108 ( .IN1(n30724), .IN2(n30721), .QN(n34099) );
  NAND2X0 U20109 ( .IN1(n30733), .IN2(n34099), .QN(n18499) );
  NOR2X0 U20110 ( .IN1(n18500), .IN2(n18499), .QN(n18507) );
  NOR2X0 U20111 ( .IN1(\s4/msel/gnt_p1 [0]), .IN2(n34389), .QN(n30718) );
  NAND2X0 U20112 ( .IN1(n30718), .IN2(n30764), .QN(n18501) );
  NOR2X0 U20113 ( .IN1(n34246), .IN2(n34389), .QN(n18504) );
  NAND2X0 U20114 ( .IN1(n30717), .IN2(n18504), .QN(n30778) );
  NAND3X0 U20115 ( .IN1(n18501), .IN2(n30778), .IN3(n34459), .QN(n30740) );
  AND2X1 U20116 ( .IN1(n34389), .IN2(n30753), .Q(n30722) );
  AO22X1 U20117 ( .IN1(n30721), .IN2(n30722), .IN3(n30718), .IN4(n30749), .Q(
        n18503) );
  NAND2X0 U20118 ( .IN1(\s4/msel/gnt_p1 [0]), .IN2(n18502), .QN(n30776) );
  OA21X1 U20119 ( .IN1(\s4/msel/gnt_p1 [0]), .IN2(n30751), .IN3(n30776), .Q(
        n30741) );
  OA22X1 U20120 ( .IN1(n18504), .IN2(n18503), .IN3(\s4/msel/gnt_p1 [1]), .IN4(
        n30741), .Q(n18505) );
  NAND2X0 U20121 ( .IN1(n30754), .IN2(n30725), .QN(n30720) );
  OR2X1 U20122 ( .IN1(n30723), .IN2(n30720), .Q(n34098) );
  NAND2X0 U20123 ( .IN1(n18505), .IN2(n34098), .QN(n18506) );
  OA22X1 U20124 ( .IN1(n18507), .IN2(n34459), .IN3(n30740), .IN4(n18506), .Q(
        n18509) );
  NAND3X0 U20125 ( .IN1(\s4/msel/gnt_p1 [0]), .IN2(\s4/msel/gnt_p1 [2]), .IN3(
        n18508), .QN(n30782) );
  NAND2X0 U20126 ( .IN1(n18509), .IN2(n30782), .QN(n17918) );
  NAND3X0 U20127 ( .IN1(n13645), .IN2(m5s10_cyc), .IN3(n34504), .QN(n32701) );
  INVX0 U20128 ( .INP(n32701), .ZN(n18578) );
  NAND2X0 U20129 ( .IN1(\s10/msel/gnt_p2 [0]), .IN2(\s10/msel/gnt_p2 [2]), 
        .QN(n18527) );
  NAND2X0 U20130 ( .IN1(\s10/msel/gnt_p2 [1]), .IN2(n34463), .QN(n18524) );
  NAND3X0 U20131 ( .IN1(n13541), .IN2(m7s10_cyc), .IN3(n34505), .QN(n18555) );
  INVX0 U20132 ( .INP(n18555), .ZN(n32696) );
  NAND3X0 U20133 ( .IN1(n13593), .IN2(m6s10_cyc), .IN3(n34568), .QN(n18550) );
  INVX0 U20134 ( .INP(n18550), .ZN(n18528) );
  NOR2X0 U20135 ( .IN1(n32696), .IN2(n18528), .QN(n32702) );
  NAND3X0 U20136 ( .IN1(n13697), .IN2(m4s10_cyc), .IN3(n34583), .QN(n18564) );
  NAND2X0 U20137 ( .IN1(n18564), .IN2(n32701), .QN(n18510) );
  NAND3X0 U20138 ( .IN1(n13749), .IN2(m3s10_cyc), .IN3(n34372), .QN(n18547) );
  OA21X1 U20139 ( .IN1(n32702), .IN2(n18510), .IN3(n18547), .Q(n18514) );
  NAND3X0 U20140 ( .IN1(n13920), .IN2(m0s10_cyc), .IN3(n34582), .QN(n18561) );
  INVX0 U20141 ( .INP(n18561), .ZN(n18584) );
  AND3X1 U20142 ( .IN1(n13853), .IN2(m1s10_cyc), .IN3(n34611), .Q(n18582) );
  NOR2X0 U20143 ( .IN1(n18584), .IN2(n18582), .QN(n18515) );
  INVX0 U20144 ( .INP(n18510), .ZN(n21771) );
  NAND2X0 U20145 ( .IN1(n18515), .IN2(n21771), .QN(n18518) );
  MUX21X1 U20146 ( .IN1(n18582), .IN2(\s10/msel/gnt_p2 [1]), .S(
        \s10/msel/gnt_p2 [0]), .Q(n32705) );
  NAND3X0 U20147 ( .IN1(n13801), .IN2(m2s10_cyc), .IN3(n34503), .QN(n18574) );
  NOR2X0 U20148 ( .IN1(n34463), .IN2(n34255), .QN(n18562) );
  INVX0 U20149 ( .INP(n18515), .ZN(n21770) );
  NAND2X0 U20150 ( .IN1(n32702), .IN2(n21770), .QN(n18511) );
  NAND4X0 U20151 ( .IN1(n18562), .IN2(n18564), .IN3(n32701), .IN4(n18511), 
        .QN(n18512) );
  OA221X1 U20152 ( .IN1(n32705), .IN2(n18514), .IN3(n32705), .IN4(n18574), 
        .IN5(n18512), .Q(n18513) );
  OA221X1 U20153 ( .IN1(n18524), .IN2(n18514), .IN3(n18524), .IN4(n18518), 
        .IN5(n18513), .Q(n18523) );
  NOR2X0 U20154 ( .IN1(\s10/msel/gnt_p2 [0]), .IN2(\s10/msel/gnt_p2 [1]), .QN(
        n18559) );
  NAND2X0 U20155 ( .IN1(n18547), .IN2(n18574), .QN(n32704) );
  NAND2X0 U20156 ( .IN1(n18515), .IN2(n32704), .QN(n18521) );
  INVX0 U20157 ( .INP(n18524), .ZN(n18516) );
  NOR2X0 U20158 ( .IN1(\s10/msel/gnt_p2 [1]), .IN2(n18528), .QN(n18517) );
  NOR2X0 U20159 ( .IN1(n18516), .IN2(n18517), .QN(n18566) );
  NOR2X0 U20160 ( .IN1(n32696), .IN2(n18566), .QN(n18519) );
  AO222X1 U20161 ( .IN1(n18519), .IN2(n18518), .IN3(n18519), .IN4(n18517), 
        .IN5(n18518), .IN6(n18562), .Q(n18520) );
  AO22X1 U20162 ( .IN1(n18559), .IN2(n18578), .IN3(n18521), .IN4(n18520), .Q(
        n18522) );
  MUX21X1 U20163 ( .IN1(n18523), .IN2(n18522), .S(\s10/msel/gnt_p2 [2]), .Q(
        n18532) );
  AO221X1 U20164 ( .IN1(n34255), .IN2(n18578), .IN3(n34255), .IN4(n18527), 
        .IN5(n18532), .Q(n18534) );
  NOR2X0 U20165 ( .IN1(n18524), .IN2(n18574), .QN(n18526) );
  INVX0 U20166 ( .INP(n18547), .ZN(n32706) );
  NAND2X0 U20167 ( .IN1(n32706), .IN2(n18562), .QN(n18586) );
  NAND2X0 U20168 ( .IN1(n18586), .IN2(n34405), .QN(n18525) );
  NOR2X0 U20169 ( .IN1(n18526), .IN2(n18525), .QN(n32708) );
  MUX21X1 U20170 ( .IN1(n18584), .IN2(n18582), .S(\s10/msel/gnt_p2 [0]), .Q(
        n32707) );
  INVX0 U20171 ( .INP(n18527), .ZN(n18577) );
  INVX0 U20172 ( .INP(n18564), .ZN(n18548) );
  NAND2X0 U20173 ( .IN1(\s10/msel/gnt_p2 [1]), .IN2(n18528), .QN(n32699) );
  AND2X1 U20174 ( .IN1(n32699), .IN2(\s10/msel/gnt_p2 [2]), .Q(n18576) );
  OA21X1 U20175 ( .IN1(n18548), .IN2(n18532), .IN3(n18576), .Q(n18530) );
  INVX0 U20176 ( .INP(n18562), .ZN(n18529) );
  OA22X1 U20177 ( .IN1(n18577), .IN2(n18530), .IN3(n18555), .IN4(n18529), .Q(
        n18531) );
  AO221X1 U20178 ( .IN1(n32708), .IN2(n18532), .IN3(n32708), .IN4(n32707), 
        .IN5(n18531), .Q(n18533) );
  NAND2X0 U20179 ( .IN1(n18534), .IN2(n18533), .QN(n17743) );
  NAND3X0 U20180 ( .IN1(n13556), .IN2(m6s3_cyc), .IN3(n34311), .QN(n19092) );
  NAND3X0 U20181 ( .IN1(n13475), .IN2(m7s3_cyc), .IN3(n34312), .QN(n18535) );
  NAND2X0 U20182 ( .IN1(n19092), .IN2(n18535), .QN(n30435) );
  AND2X1 U20183 ( .IN1(n34388), .IN2(n30435), .Q(n30429) );
  NAND3X0 U20184 ( .IN1(n13868), .IN2(m0s3_cyc), .IN3(n34309), .QN(n19091) );
  NAND3X0 U20185 ( .IN1(n13816), .IN2(m1s3_cyc), .IN3(n34310), .QN(n19078) );
  AND2X1 U20186 ( .IN1(n19091), .IN2(n19078), .Q(n30427) );
  NAND3X0 U20187 ( .IN1(n13764), .IN2(m2s3_cyc), .IN3(n34637), .QN(n19077) );
  INVX0 U20188 ( .INP(n19077), .ZN(n19106) );
  NAND3X0 U20189 ( .IN1(n13712), .IN2(m3s3_cyc), .IN3(n34616), .QN(n19076) );
  INVX0 U20190 ( .INP(n19076), .ZN(n30425) );
  NOR2X0 U20191 ( .IN1(n19106), .IN2(n30425), .QN(n30434) );
  NAND2X0 U20192 ( .IN1(n30427), .IN2(n30434), .QN(n21801) );
  INVX0 U20193 ( .INP(n21801), .ZN(n18537) );
  NAND3X0 U20194 ( .IN1(n13608), .IN2(m5s3_cyc), .IN3(n34361), .QN(n19079) );
  INVX0 U20195 ( .INP(n19079), .ZN(n30445) );
  INVX0 U20196 ( .INP(n18535), .ZN(n30440) );
  MUX21X1 U20197 ( .IN1(n30445), .IN2(n30440), .S(\s3/msel/gnt_p1 [1]), .Q(
        n18545) );
  NAND3X0 U20198 ( .IN1(n13660), .IN2(m4s3_cyc), .IN3(n34236), .QN(n19090) );
  INVX0 U20199 ( .INP(n19090), .ZN(n30446) );
  INVX0 U20200 ( .INP(n19092), .ZN(n30442) );
  MUX21X1 U20201 ( .IN1(n30446), .IN2(n30442), .S(\s3/msel/gnt_p1 [1]), .Q(
        n19111) );
  OA21X1 U20202 ( .IN1(n18545), .IN2(n19111), .IN3(n34658), .Q(n18536) );
  NOR3X0 U20203 ( .IN1(n30429), .IN2(n18537), .IN3(n18536), .QN(n18544) );
  NOR2X0 U20204 ( .IN1(\s3/msel/gnt_p1 [0]), .IN2(n34388), .QN(n30441) );
  NAND2X0 U20205 ( .IN1(n30441), .IN2(n19106), .QN(n18538) );
  NOR2X0 U20206 ( .IN1(n34658), .IN2(n34388), .QN(n30439) );
  NAND2X0 U20207 ( .IN1(n30425), .IN2(n30439), .QN(n19108) );
  NAND3X0 U20208 ( .IN1(n18538), .IN2(n19108), .IN3(n34418), .QN(n30437) );
  NOR2X0 U20209 ( .IN1(\s3/msel/gnt_p1 [1]), .IN2(n34658), .QN(n19075) );
  AO21X1 U20210 ( .IN1(n19075), .IN2(n19077), .IN3(n30441), .Q(n19097) );
  NAND2X0 U20211 ( .IN1(n34658), .IN2(n34388), .QN(n30430) );
  INVX0 U20212 ( .INP(n30430), .ZN(n18539) );
  NAND2X0 U20213 ( .IN1(n18539), .IN2(n19078), .QN(n30422) );
  NOR2X0 U20214 ( .IN1(n19106), .IN2(n30422), .QN(n18540) );
  OA21X1 U20215 ( .IN1(n19097), .IN2(n18540), .IN3(n19076), .Q(n18541) );
  MUX21X1 U20216 ( .IN1(n19091), .IN2(n19078), .S(\s3/msel/gnt_p1 [0]), .Q(
        n30438) );
  OA22X1 U20217 ( .IN1(n30439), .IN2(n18541), .IN3(\s3/msel/gnt_p1 [1]), .IN4(
        n30438), .Q(n18542) );
  NAND2X0 U20218 ( .IN1(n19079), .IN2(n19090), .QN(n30421) );
  OR2X1 U20219 ( .IN1(n30435), .IN2(n30421), .Q(n21800) );
  NAND2X0 U20220 ( .IN1(n18542), .IN2(n21800), .QN(n18543) );
  OA22X1 U20221 ( .IN1(n18544), .IN2(n34418), .IN3(n30437), .IN4(n18543), .Q(
        n18546) );
  NAND3X0 U20222 ( .IN1(\s3/msel/gnt_p1 [0]), .IN2(\s3/msel/gnt_p1 [2]), .IN3(
        n18545), .QN(n19115) );
  NAND2X0 U20223 ( .IN1(n18546), .IN2(n19115), .QN(n17946) );
  NAND2X0 U20224 ( .IN1(n18548), .IN2(n34255), .QN(n32698) );
  NAND2X0 U20225 ( .IN1(n18550), .IN2(n18564), .QN(n18553) );
  NOR2X0 U20226 ( .IN1(n34463), .IN2(n18553), .QN(n18549) );
  OA21X1 U20227 ( .IN1(n32701), .IN2(n18548), .IN3(n18547), .Q(n18557) );
  INVX0 U20228 ( .INP(n18557), .ZN(n18565) );
  AO221X1 U20229 ( .IN1(n18574), .IN2(n18549), .IN3(n18574), .IN4(n18565), 
        .IN5(n18582), .Q(n18560) );
  NAND2X0 U20230 ( .IN1(n18559), .IN2(n18560), .QN(n18552) );
  AO21X1 U20231 ( .IN1(n18582), .IN2(n18561), .IN3(n32696), .Q(n18563) );
  AO21X1 U20232 ( .IN1(n18550), .IN2(n18563), .IN3(n18578), .Q(n18558) );
  NAND3X0 U20233 ( .IN1(n18562), .IN2(n18564), .IN3(n18558), .QN(n18551) );
  NAND3X0 U20234 ( .IN1(n18552), .IN2(n34405), .IN3(n18551), .QN(n18575) );
  NOR2X0 U20235 ( .IN1(\s10/msel/gnt_p2 [0]), .IN2(n18582), .QN(n18554) );
  AO221X1 U20236 ( .IN1(n18555), .IN2(n18584), .IN3(n18555), .IN4(n18554), 
        .IN5(n18553), .Q(n18556) );
  NAND2X0 U20237 ( .IN1(n18557), .IN2(n18556), .QN(n18573) );
  NAND2X0 U20238 ( .IN1(n18559), .IN2(n18558), .QN(n18571) );
  NAND3X0 U20239 ( .IN1(n18562), .IN2(n18561), .IN3(n18560), .QN(n18570) );
  INVX0 U20240 ( .INP(n18563), .ZN(n18568) );
  OAI221X1 U20241 ( .IN1(n18565), .IN2(n18564), .IN3(n18565), .IN4(
        \s10/msel/gnt_p2 [0]), .IN5(n18574), .QN(n18567) );
  AO221X1 U20242 ( .IN1(n18568), .IN2(n18584), .IN3(n18568), .IN4(n18567), 
        .IN5(n18566), .Q(n18569) );
  NAND4X0 U20243 ( .IN1(\s10/msel/gnt_p2 [2]), .IN2(n18571), .IN3(n18570), 
        .IN4(n18569), .QN(n18572) );
  OA221X1 U20244 ( .IN1(n18575), .IN2(n18574), .IN3(n18575), .IN4(n18573), 
        .IN5(n18572), .Q(n18581) );
  OA221X1 U20245 ( .IN1(\s10/msel/gnt_p2 [0]), .IN2(n18576), .IN3(
        \s10/msel/gnt_p2 [0]), .IN4(n32698), .IN5(n18581), .Q(n18580) );
  OA221X1 U20246 ( .IN1(\s10/msel/gnt_p2 [1]), .IN2(n18578), .IN3(n34255), 
        .IN4(n32696), .IN5(n18577), .Q(n18579) );
  NOR2X0 U20247 ( .IN1(n18580), .IN2(n18579), .QN(n18590) );
  INVX0 U20248 ( .INP(n18581), .ZN(n18585) );
  NAND2X0 U20249 ( .IN1(\s10/msel/gnt_p2 [0]), .IN2(n18582), .QN(n18583) );
  OA222X1 U20250 ( .IN1(n18585), .IN2(n18584), .IN3(n18585), .IN4(n34255), 
        .IN5(\s10/msel/gnt_p2 [1]), .IN6(n18583), .Q(n18587) );
  NAND2X0 U20251 ( .IN1(n18587), .IN2(n18586), .QN(n18588) );
  NAND2X0 U20252 ( .IN1(n34405), .IN2(n18588), .QN(n18589) );
  NAND2X0 U20253 ( .IN1(n18590), .IN2(n18589), .QN(n17742) );
  NAND2X0 U20254 ( .IN1(m5s14_cyc), .IN2(n34652), .QN(n18757) );
  NOR2X0 U20255 ( .IN1(n34547), .IN2(n18757), .QN(n33718) );
  NAND2X0 U20256 ( .IN1(\s14/msel/gnt_p2 [0]), .IN2(\s14/msel/gnt_p2 [2]), 
        .QN(n33754) );
  NOR2X0 U20257 ( .IN1(n34271), .IN2(n34381), .QN(n18609) );
  NAND3X0 U20258 ( .IN1(n13693), .IN2(m4s14_cyc), .IN3(n34571), .QN(n33735) );
  NAND2X0 U20259 ( .IN1(n18609), .IN2(n33735), .QN(n33721) );
  NAND3X0 U20260 ( .IN1(n13589), .IN2(m6s14_cyc), .IN3(n34544), .QN(n33730) );
  INVX0 U20261 ( .INP(n33730), .ZN(n33717) );
  NAND3X0 U20262 ( .IN1(n13537), .IN2(m7s14_cyc), .IN3(n34513), .QN(n33756) );
  INVX0 U20263 ( .INP(n33756), .ZN(n18610) );
  NOR2X0 U20264 ( .IN1(n33717), .IN2(n18610), .QN(n33707) );
  AND3X1 U20265 ( .IN1(n13912), .IN2(m0s14_cyc), .IN3(n34604), .Q(n33751) );
  NAND3X0 U20266 ( .IN1(n13849), .IN2(m1s14_cyc), .IN3(n34512), .QN(n33719) );
  INVX0 U20267 ( .INP(n33719), .ZN(n33749) );
  NOR2X0 U20268 ( .IN1(n33751), .IN2(n33749), .QN(n18597) );
  INVX0 U20269 ( .INP(n18597), .ZN(n21766) );
  AO221X1 U20270 ( .IN1(n33707), .IN2(n34381), .IN3(n33707), .IN4(n21766), 
        .IN5(n33718), .Q(n18595) );
  NOR2X0 U20271 ( .IN1(\s14/msel/gnt_p2 [0]), .IN2(n34381), .QN(n18611) );
  INVX0 U20272 ( .INP(n18611), .ZN(n18594) );
  NAND2X0 U20273 ( .IN1(m3s14_cyc), .IN2(n34648), .QN(n18755) );
  NOR2X0 U20274 ( .IN1(n34481), .IN2(n18755), .QN(n33731) );
  INVX0 U20275 ( .INP(n33718), .ZN(n33755) );
  NAND2X0 U20276 ( .IN1(n33755), .IN2(n33735), .QN(n21765) );
  NOR2X0 U20277 ( .IN1(n21766), .IN2(n21765), .QN(n18599) );
  NOR2X0 U20278 ( .IN1(n33707), .IN2(n21765), .QN(n18591) );
  NOR3X0 U20279 ( .IN1(n33731), .IN2(n18599), .IN3(n18591), .QN(n18593) );
  NAND2X0 U20280 ( .IN1(m2s14_cyc), .IN2(n34646), .QN(n18756) );
  NOR2X0 U20281 ( .IN1(n34477), .IN2(n18756), .QN(n33729) );
  OR2X1 U20282 ( .IN1(n33729), .IN2(n33731), .Q(n33705) );
  NOR2X0 U20283 ( .IN1(n18591), .IN2(n33705), .QN(n18592) );
  NAND2X0 U20284 ( .IN1(n34271), .IN2(n34381), .QN(n33732) );
  NAND2X0 U20285 ( .IN1(\s14/msel/gnt_p2 [0]), .IN2(n34381), .QN(n18598) );
  OA21X1 U20286 ( .IN1(n33749), .IN2(n33732), .IN3(n18598), .Q(n33706) );
  OA222X1 U20287 ( .IN1(n33721), .IN2(n18595), .IN3(n18594), .IN4(n18593), 
        .IN5(n18592), .IN6(n33706), .Q(n18607) );
  INVX0 U20288 ( .INP(n18595), .ZN(n18596) );
  NOR2X0 U20289 ( .IN1(n18596), .IN2(n33732), .QN(n18605) );
  NAND2X0 U20290 ( .IN1(n18597), .IN2(n33705), .QN(n18604) );
  NOR2X0 U20291 ( .IN1(n33717), .IN2(n18598), .QN(n18600) );
  NOR2X0 U20292 ( .IN1(n18611), .IN2(n18600), .QN(n33740) );
  NOR2X0 U20293 ( .IN1(n18610), .IN2(n33740), .QN(n18602) );
  INVX0 U20294 ( .INP(n18599), .ZN(n18601) );
  AO222X1 U20295 ( .IN1(n18602), .IN2(n18601), .IN3(n18602), .IN4(n18600), 
        .IN5(n18601), .IN6(n18609), .Q(n18603) );
  AO222X1 U20296 ( .IN1(n18605), .IN2(n18604), .IN3(n18605), .IN4(n33718), 
        .IN5(n18604), .IN6(n18603), .Q(n18606) );
  MUX21X1 U20297 ( .IN1(n18607), .IN2(n18606), .S(\s14/msel/gnt_p2 [2]), .Q(
        n18615) );
  AO221X1 U20298 ( .IN1(n34381), .IN2(n33718), .IN3(n34381), .IN4(n33754), 
        .IN5(n18615), .Q(n18617) );
  NAND2X0 U20299 ( .IN1(n33731), .IN2(n18609), .QN(n33752) );
  NAND2X0 U20300 ( .IN1(n33729), .IN2(n18611), .QN(n18608) );
  AND3X1 U20301 ( .IN1(n34460), .IN2(n33752), .IN3(n18608), .Q(n33713) );
  MUX21X1 U20302 ( .IN1(n33751), .IN2(n33749), .S(\s14/msel/gnt_p2 [0]), .Q(
        n33709) );
  INVX0 U20303 ( .INP(n33735), .ZN(n33702) );
  NOR3X0 U20304 ( .IN1(\s14/msel/gnt_p2 [0]), .IN2(n33702), .IN3(n18615), .QN(
        n18613) );
  AO22X1 U20305 ( .IN1(n33717), .IN2(n18611), .IN3(n18610), .IN4(n18609), .Q(
        n18612) );
  NOR3X0 U20306 ( .IN1(n18613), .IN2(n34460), .IN3(n18612), .QN(n18614) );
  AO221X1 U20307 ( .IN1(n33713), .IN2(n18615), .IN3(n33713), .IN4(n33709), 
        .IN5(n18614), .Q(n18616) );
  NAND2X0 U20308 ( .IN1(n18617), .IN2(n18616), .QN(n17631) );
  NAND3X0 U20309 ( .IN1(n13848), .IN2(n13822), .IN3(m1s13_cyc), .QN(n18620) );
  INVX0 U20310 ( .INP(n18620), .ZN(n33395) );
  NAND2X0 U20311 ( .IN1(\s13/msel/gnt_p0 [0]), .IN2(n33395), .QN(n33397) );
  NOR2X0 U20312 ( .IN1(n33397), .IN2(\s13/msel/gnt_p0 [1]), .QN(n18649) );
  NAND3X0 U20313 ( .IN1(n13796), .IN2(n13770), .IN3(m2s13_cyc), .QN(n18619) );
  INVX0 U20314 ( .INP(n18619), .ZN(n33392) );
  NAND3X0 U20315 ( .IN1(n13910), .IN2(n13874), .IN3(m0s13_cyc), .QN(n33398) );
  INVX0 U20316 ( .INP(n33398), .ZN(n33388) );
  NAND3X0 U20317 ( .IN1(n13588), .IN2(n13562), .IN3(m6s13_cyc), .QN(n33383) );
  INVX0 U20318 ( .INP(n33383), .ZN(n33442) );
  NAND3X0 U20319 ( .IN1(n13692), .IN2(n13666), .IN3(m4s13_cyc), .QN(n33412) );
  INVX0 U20320 ( .INP(n33412), .ZN(n33439) );
  NOR2X0 U20321 ( .IN1(n33442), .IN2(n33439), .QN(n18634) );
  NAND3X0 U20322 ( .IN1(n13640), .IN2(n13614), .IN3(m5s13_cyc), .QN(n33411) );
  INVX0 U20323 ( .INP(n33411), .ZN(n33438) );
  AND3X1 U20324 ( .IN1(n13744), .IN2(n13718), .IN3(m3s13_cyc), .Q(n33409) );
  AO21X1 U20325 ( .IN1(n33438), .IN2(n33412), .IN3(n33409), .Q(n18635) );
  AO21X1 U20326 ( .IN1(\s13/msel/gnt_p0 [0]), .IN2(n18634), .IN3(n18635), .Q(
        n18618) );
  AO21X1 U20327 ( .IN1(n18619), .IN2(n18618), .IN3(n33395), .Q(n18631) );
  NAND3X0 U20328 ( .IN1(\s13/msel/gnt_p0 [1]), .IN2(n18631), .IN3(n33398), 
        .QN(n18630) );
  NAND2X0 U20329 ( .IN1(n18619), .IN2(n33398), .QN(n18622) );
  NAND3X0 U20330 ( .IN1(n13536), .IN2(n13482), .IN3(m7s13_cyc), .QN(n33385) );
  OA21X1 U20331 ( .IN1(n33388), .IN2(n18620), .IN3(n33385), .Q(n18639) );
  OA21X1 U20332 ( .IN1(n34653), .IN2(n18622), .IN3(n18639), .Q(n18621) );
  OA21X1 U20333 ( .IN1(n33442), .IN2(n18621), .IN3(n33411), .Q(n18641) );
  INVX0 U20334 ( .INP(n18622), .ZN(n18625) );
  NAND3X0 U20335 ( .IN1(n18625), .IN2(n33409), .IN3(n33383), .QN(n18623) );
  NAND2X0 U20336 ( .IN1(n34653), .IN2(n34264), .QN(n33424) );
  AO21X1 U20337 ( .IN1(n18641), .IN2(n18623), .IN3(n33424), .Q(n18629) );
  NOR2X0 U20338 ( .IN1(\s13/msel/gnt_p0 [0]), .IN2(n34264), .QN(n33408) );
  NAND2X0 U20339 ( .IN1(\s13/msel/gnt_p0 [0]), .IN2(n34264), .QN(n33414) );
  NOR2X0 U20340 ( .IN1(n33442), .IN2(n33414), .QN(n33386) );
  NAND3X0 U20341 ( .IN1(n18625), .IN2(\s13/msel/gnt_p0 [0]), .IN3(n33412), 
        .QN(n18624) );
  NAND2X0 U20342 ( .IN1(n18624), .IN2(n18639), .QN(n18627) );
  AND2X1 U20343 ( .IN1(n18635), .IN2(n18625), .Q(n18626) );
  OAI22X1 U20344 ( .IN1(n33408), .IN2(n33386), .IN3(n18627), .IN4(n18626), 
        .QN(n18628) );
  NAND4X0 U20345 ( .IN1(\s13/msel/gnt_p0 [2]), .IN2(n18630), .IN3(n18629), 
        .IN4(n18628), .QN(n18646) );
  INVX0 U20346 ( .INP(n18631), .ZN(n18633) );
  INVX0 U20347 ( .INP(n18634), .ZN(n18638) );
  OR3X1 U20348 ( .IN1(n33385), .IN2(n18638), .IN3(n33392), .Q(n18632) );
  AO21X1 U20349 ( .IN1(n18633), .IN2(n18632), .IN3(n33424), .Q(n18644) );
  AND3X1 U20350 ( .IN1(n33398), .IN2(n18634), .IN3(\s13/msel/gnt_p0 [0]), .Q(
        n18636) );
  NOR2X0 U20351 ( .IN1(n18636), .IN2(n18635), .QN(n18640) );
  INVX0 U20352 ( .INP(n33408), .ZN(n18637) );
  OA21X1 U20353 ( .IN1(n33392), .IN2(n33414), .IN3(n18637), .Q(n33396) );
  AO221X1 U20354 ( .IN1(n18640), .IN2(n18639), .IN3(n18640), .IN4(n18638), 
        .IN5(n33396), .Q(n18643) );
  OR3X1 U20355 ( .IN1(n34264), .IN2(n18641), .IN3(n33439), .Q(n18642) );
  NAND4X0 U20356 ( .IN1(n34292), .IN2(n18644), .IN3(n18643), .IN4(n18642), 
        .QN(n18645) );
  NAND2X0 U20357 ( .IN1(n18646), .IN2(n18645), .QN(n18650) );
  AO221X1 U20358 ( .IN1(\s13/msel/gnt_p0 [1]), .IN2(n33392), .IN3(n34264), 
        .IN4(n33388), .IN5(n18650), .Q(n18647) );
  NOR2X0 U20359 ( .IN1(n34653), .IN2(n34264), .QN(n33400) );
  NAND2X0 U20360 ( .IN1(n33409), .IN2(n33400), .QN(n33393) );
  NAND2X0 U20361 ( .IN1(n18647), .IN2(n33393), .QN(n18648) );
  NOR2X0 U20362 ( .IN1(n18649), .IN2(n18648), .QN(n18652) );
  MUX21X1 U20363 ( .IN1(n33439), .IN2(n33442), .S(\s13/msel/gnt_p0 [1]), .Q(
        n33389) );
  OA21X1 U20364 ( .IN1(n34292), .IN2(n33389), .IN3(n34653), .Q(n18651) );
  OA22X1 U20365 ( .IN1(\s13/msel/gnt_p0 [2]), .IN2(n18652), .IN3(n18651), 
        .IN4(n18650), .Q(n18653) );
  NAND2X0 U20366 ( .IN1(\s13/msel/gnt_p0 [1]), .IN2(n33385), .QN(n33387) );
  NAND2X0 U20367 ( .IN1(n34264), .IN2(n33411), .QN(n33384) );
  NAND4X0 U20368 ( .IN1(\s13/msel/gnt_p0 [2]), .IN2(\s13/msel/gnt_p0 [0]), 
        .IN3(n33387), .IN4(n33384), .QN(n33406) );
  NAND2X0 U20369 ( .IN1(n18653), .IN2(n33406), .QN(n17661) );
  NAND3X0 U20370 ( .IN1(n13771), .IN2(m2s14_cyc), .IN3(n34477), .QN(n18843) );
  NAND3X0 U20371 ( .IN1(n13719), .IN2(m3s14_cyc), .IN3(n34481), .QN(n33625) );
  NAND2X0 U20372 ( .IN1(n18843), .IN2(n33625), .QN(n33612) );
  NAND3X0 U20373 ( .IN1(n13875), .IN2(m0s14_cyc), .IN3(n34367), .QN(n18842) );
  NAND3X0 U20374 ( .IN1(n13823), .IN2(m1s14_cyc), .IN3(n34334), .QN(n18864) );
  NAND2X0 U20375 ( .IN1(n18842), .IN2(n18864), .QN(n33613) );
  NOR2X0 U20376 ( .IN1(n33612), .IN2(n33613), .QN(n34213) );
  NAND3X0 U20377 ( .IN1(n13563), .IN2(m6s14_cyc), .IN3(n34357), .QN(n18841) );
  NAND3X0 U20378 ( .IN1(n13484), .IN2(m7s14_cyc), .IN3(n34358), .QN(n18844) );
  NAND2X0 U20379 ( .IN1(n18841), .IN2(n18844), .QN(n33614) );
  NAND3X0 U20380 ( .IN1(n13615), .IN2(m5s14_cyc), .IN3(n34547), .QN(n33632) );
  NAND2X0 U20381 ( .IN1(n34242), .IN2(n33632), .QN(n18662) );
  NAND2X0 U20382 ( .IN1(\s14/msel/gnt_p1 [1]), .IN2(n18844), .QN(n18663) );
  OA21X1 U20383 ( .IN1(n33614), .IN2(n34394), .IN3(n18663), .Q(n33617) );
  OA21X1 U20384 ( .IN1(n33614), .IN2(n18662), .IN3(n33617), .Q(n18654) );
  NOR3X0 U20385 ( .IN1(n34213), .IN2(n18654), .IN3(n34386), .QN(n18661) );
  NAND3X0 U20386 ( .IN1(n13667), .IN2(m4s14_cyc), .IN3(n34635), .QN(n33631) );
  OA221X1 U20387 ( .IN1(\s14/msel/gnt_p1 [1]), .IN2(n33631), .IN3(n34242), 
        .IN4(n18841), .IN5(\s14/msel/gnt_p1 [2]), .Q(n18655) );
  NOR2X0 U20388 ( .IN1(\s14/msel/gnt_p1 [0]), .IN2(n18655), .QN(n18868) );
  INVX0 U20389 ( .INP(n18868), .ZN(n18660) );
  AO221X1 U20390 ( .IN1(n34394), .IN2(n18843), .IN3(\s14/msel/gnt_p1 [0]), 
        .IN4(n33625), .IN5(n34242), .Q(n33636) );
  OA21X1 U20391 ( .IN1(\s14/msel/gnt_p1 [0]), .IN2(n18842), .IN3(n18864), .Q(
        n33638) );
  INVX0 U20392 ( .INP(n33612), .ZN(n33626) );
  NOR2X0 U20393 ( .IN1(n34394), .IN2(n34242), .QN(n18656) );
  OA22X1 U20394 ( .IN1(\s14/msel/gnt_p1 [1]), .IN2(n33638), .IN3(n33626), 
        .IN4(n18656), .Q(n18658) );
  INVX0 U20395 ( .INP(n33614), .ZN(n34215) );
  AND2X1 U20396 ( .IN1(n33632), .IN2(n33631), .Q(n34214) );
  NAND2X0 U20397 ( .IN1(n34215), .IN2(n34214), .QN(n18657) );
  NAND3X0 U20398 ( .IN1(n33636), .IN2(n18658), .IN3(n18657), .QN(n18659) );
  AO22X1 U20399 ( .IN1(n18661), .IN2(n18660), .IN3(n18659), .IN4(n34386), .Q(
        n18664) );
  NAND4X0 U20400 ( .IN1(\s14/msel/gnt_p1 [2]), .IN2(\s14/msel/gnt_p1 [0]), 
        .IN3(n18663), .IN4(n18662), .QN(n18870) );
  NAND2X0 U20401 ( .IN1(n18664), .IN2(n18870), .QN(n17638) );
  NAND3X0 U20402 ( .IN1(n13724), .IN2(m3s11_cyc), .IN3(n34365), .QN(n32811) );
  NAND2X0 U20403 ( .IN1(\s11/msel/gnt_p1 [0]), .IN2(\s11/msel/gnt_p1 [1]), 
        .QN(n18697) );
  NOR2X0 U20404 ( .IN1(n32811), .IN2(n18697), .QN(n32800) );
  NAND3X0 U20405 ( .IN1(n13776), .IN2(m2s11_cyc), .IN3(n34325), .QN(n18680) );
  INVX0 U20406 ( .INP(n18680), .ZN(n32801) );
  NAND3X0 U20407 ( .IN1(n13620), .IN2(m5s11_cyc), .IN3(n34375), .QN(n32797) );
  INVX0 U20408 ( .INP(n32797), .ZN(n32835) );
  NAND3X0 U20409 ( .IN1(n13672), .IN2(m4s11_cyc), .IN3(n34622), .QN(n32836) );
  NAND2X0 U20410 ( .IN1(n32835), .IN2(n32836), .QN(n18673) );
  NAND2X0 U20411 ( .IN1(n32811), .IN2(n18673), .QN(n18667) );
  NAND3X0 U20412 ( .IN1(n13568), .IN2(m6s11_cyc), .IN3(n34633), .QN(n32788) );
  INVX0 U20413 ( .INP(n32788), .ZN(n32832) );
  NAND3X0 U20414 ( .IN1(n13880), .IN2(m0s11_cyc), .IN3(n34621), .QN(n32799) );
  INVX0 U20415 ( .INP(n32799), .ZN(n32791) );
  NAND3X0 U20416 ( .IN1(n13828), .IN2(m1s11_cyc), .IN3(n34326), .QN(n32798) );
  NAND3X0 U20417 ( .IN1(n13495), .IN2(m7s11_cyc), .IN3(n34324), .QN(n32789) );
  OA21X1 U20418 ( .IN1(n32791), .IN2(n32798), .IN3(n32789), .Q(n18677) );
  NOR2X0 U20419 ( .IN1(n32832), .IN2(n18677), .QN(n18671) );
  NAND2X0 U20420 ( .IN1(\s11/msel/gnt_p1 [0]), .IN2(n32836), .QN(n18672) );
  NOR2X0 U20421 ( .IN1(n32832), .IN2(n18672), .QN(n18666) );
  AO22X1 U20422 ( .IN1(n18671), .IN2(n32836), .IN3(n18666), .IN4(n32799), .Q(
        n18665) );
  NOR2X0 U20423 ( .IN1(n18667), .IN2(n18665), .QN(n18669) );
  INVX0 U20424 ( .INP(n32798), .ZN(n32790) );
  AO221X1 U20425 ( .IN1(n18680), .IN2(n18667), .IN3(n18680), .IN4(n18666), 
        .IN5(n32790), .Q(n18679) );
  INVX0 U20426 ( .INP(n18679), .ZN(n18668) );
  NAND2X0 U20427 ( .IN1(n34655), .IN2(n34390), .QN(n32824) );
  OA22X1 U20428 ( .IN1(n32801), .IN2(n18669), .IN3(n18668), .IN4(n32824), .Q(
        n18670) );
  NAND2X0 U20429 ( .IN1(n18670), .IN2(n34425), .QN(n18688) );
  NOR2X0 U20430 ( .IN1(n34390), .IN2(n18672), .QN(n32814) );
  NOR2X0 U20431 ( .IN1(n32835), .IN2(n18671), .QN(n18682) );
  INVX0 U20432 ( .INP(n18682), .ZN(n18687) );
  NAND3X0 U20433 ( .IN1(n18673), .IN2(n18672), .IN3(n32811), .QN(n18675) );
  NOR2X0 U20434 ( .IN1(n32791), .IN2(n32801), .QN(n18674) );
  NAND2X0 U20435 ( .IN1(n18675), .IN2(n18674), .QN(n18678) );
  NAND3X0 U20436 ( .IN1(\s11/msel/gnt_p1 [0]), .IN2(n34390), .IN3(n32788), 
        .QN(n32785) );
  NOR2X0 U20437 ( .IN1(\s11/msel/gnt_p1 [0]), .IN2(n34390), .QN(n32833) );
  INVX0 U20438 ( .INP(n32833), .ZN(n18676) );
  AO22X1 U20439 ( .IN1(n18678), .IN2(n18677), .IN3(n32785), .IN4(n18676), .Q(
        n18685) );
  NAND3X0 U20440 ( .IN1(\s11/msel/gnt_p1 [1]), .IN2(n18679), .IN3(n32799), 
        .QN(n18684) );
  INVX0 U20441 ( .INP(n32811), .ZN(n32796) );
  NAND3X0 U20442 ( .IN1(n32796), .IN2(n32799), .IN3(n18680), .QN(n18681) );
  AO221X1 U20443 ( .IN1(n18682), .IN2(n32832), .IN3(n18682), .IN4(n18681), 
        .IN5(n32824), .Q(n18683) );
  NAND4X0 U20444 ( .IN1(\s11/msel/gnt_p1 [2]), .IN2(n18685), .IN3(n18684), 
        .IN4(n18683), .QN(n18686) );
  OA221X1 U20445 ( .IN1(n18688), .IN2(n32814), .IN3(n18688), .IN4(n18687), 
        .IN5(n18686), .Q(n18692) );
  NOR2X0 U20446 ( .IN1(n34655), .IN2(n32798), .QN(n18689) );
  AO222X1 U20447 ( .IN1(n18692), .IN2(\s11/msel/gnt_p1 [1]), .IN3(n18692), 
        .IN4(n32799), .IN5(n34390), .IN6(n18689), .Q(n18690) );
  NOR2X0 U20448 ( .IN1(n32800), .IN2(n18690), .QN(n18695) );
  MUX21X1 U20449 ( .IN1(n32836), .IN2(n32788), .S(\s11/msel/gnt_p1 [1]), .Q(
        n18691) );
  INVX0 U20450 ( .INP(n18691), .ZN(n32792) );
  OA21X1 U20451 ( .IN1(n34425), .IN2(n32792), .IN3(n34655), .Q(n18694) );
  INVX0 U20452 ( .INP(n18692), .ZN(n18693) );
  OA22X1 U20453 ( .IN1(\s11/msel/gnt_p1 [2]), .IN2(n18695), .IN3(n18694), 
        .IN4(n18693), .Q(n18700) );
  INVX0 U20454 ( .INP(n32789), .ZN(n32786) );
  NOR2X0 U20455 ( .IN1(n32786), .IN2(n34390), .QN(n32787) );
  NOR2X0 U20456 ( .IN1(n32787), .IN2(n34425), .QN(n18699) );
  NAND2X0 U20457 ( .IN1(\s11/msel/gnt_p1 [0]), .IN2(n32835), .QN(n18696) );
  NAND2X0 U20458 ( .IN1(n18697), .IN2(n18696), .QN(n18698) );
  NAND2X0 U20459 ( .IN1(n18699), .IN2(n18698), .QN(n32807) );
  NAND2X0 U20460 ( .IN1(n18700), .IN2(n32807), .QN(n17720) );
  NAND2X0 U20461 ( .IN1(n32008), .IN2(n32005), .QN(n31985) );
  INVX0 U20462 ( .INP(n31985), .ZN(n18715) );
  NOR2X0 U20463 ( .IN1(\s8/msel/gnt_p1 [1]), .IN2(n18715), .QN(n31997) );
  NAND2X0 U20464 ( .IN1(n18706), .IN2(n31988), .QN(n31986) );
  NOR2X0 U20465 ( .IN1(n18701), .IN2(n18709), .QN(n31994) );
  INVX0 U20466 ( .INP(n31994), .ZN(n18702) );
  NOR2X0 U20467 ( .IN1(n31986), .IN2(n18702), .QN(n34145) );
  OA21X1 U20468 ( .IN1(n18704), .IN2(n18703), .IN3(n34229), .Q(n18705) );
  NOR3X0 U20469 ( .IN1(n31997), .IN2(n34145), .IN3(n18705), .QN(n18718) );
  OR2X1 U20470 ( .IN1(n32007), .IN2(n18706), .Q(n18708) );
  NAND3X0 U20471 ( .IN1(n18708), .IN2(n18707), .IN3(n34420), .QN(n32002) );
  OAI22X1 U20472 ( .IN1(n18711), .IN2(n18710), .IN3(n18709), .IN4(n31986), 
        .QN(n18714) );
  OA21X1 U20473 ( .IN1(\s8/msel/gnt_p1 [0]), .IN2(n18713), .IN3(n18712), .Q(
        n32003) );
  OA22X1 U20474 ( .IN1(n32004), .IN2(n18714), .IN3(\s8/msel/gnt_p1 [1]), .IN4(
        n32003), .Q(n18716) );
  NOR2X0 U20475 ( .IN1(n32011), .IN2(n32009), .QN(n31984) );
  NAND2X0 U20476 ( .IN1(n18715), .IN2(n31984), .QN(n34141) );
  NAND2X0 U20477 ( .IN1(n18716), .IN2(n34141), .QN(n18717) );
  OA22X1 U20478 ( .IN1(n18718), .IN2(n34420), .IN3(n32002), .IN4(n18717), .Q(
        n18720) );
  NAND2X0 U20479 ( .IN1(n18720), .IN2(n18719), .QN(n17806) );
  NAND3X0 U20480 ( .IN1(n13684), .IN2(m4s1_cyc), .IN3(n34483), .QN(n29999) );
  NAND3X0 U20481 ( .IN1(n13580), .IN2(m6s1_cyc), .IN3(n34522), .QN(n18895) );
  MUX21X1 U20482 ( .IN1(n29999), .IN2(n18895), .S(\s1/msel/gnt_p2 [1]), .Q(
        n18910) );
  NOR2X0 U20483 ( .IN1(\s1/msel/gnt_p2 [1]), .IN2(\s1/msel/gnt_p2 [0]), .QN(
        n18729) );
  NAND3X0 U20484 ( .IN1(n13788), .IN2(m2s1_cyc), .IN3(n34558), .QN(n18897) );
  INVX0 U20485 ( .INP(n18897), .ZN(n18900) );
  NAND3X0 U20486 ( .IN1(n13528), .IN2(m7s1_cyc), .IN3(n34559), .QN(n18894) );
  NAND2X0 U20487 ( .IN1(n18895), .IN2(n29999), .QN(n18722) );
  OR3X1 U20488 ( .IN1(n18900), .IN2(n18894), .IN3(n18722), .Q(n18721) );
  INVX0 U20489 ( .INP(n29999), .ZN(n18730) );
  NAND3X0 U20490 ( .IN1(n13632), .IN2(m5s1_cyc), .IN3(n34556), .QN(n29996) );
  NAND3X0 U20491 ( .IN1(n13736), .IN2(m3s1_cyc), .IN3(n34521), .QN(n29989) );
  OA21X1 U20492 ( .IN1(n18730), .IN2(n29996), .IN3(n29989), .Q(n18733) );
  NAND3X0 U20493 ( .IN1(n13840), .IN2(m1s1_cyc), .IN3(n34555), .QN(n18905) );
  OA21X1 U20494 ( .IN1(n18900), .IN2(n18733), .IN3(n18905), .Q(n18738) );
  NAND2X0 U20495 ( .IN1(n18721), .IN2(n18738), .QN(n18728) );
  INVX0 U20496 ( .INP(n18729), .ZN(n29974) );
  NAND3X0 U20497 ( .IN1(n13898), .IN2(m0s1_cyc), .IN3(n34557), .QN(n18906) );
  INVX0 U20498 ( .INP(n18906), .ZN(n18748) );
  OA21X1 U20499 ( .IN1(n18748), .IN2(n18905), .IN3(n18894), .Q(n18731) );
  NOR2X0 U20500 ( .IN1(n18731), .IN2(n18722), .QN(n18725) );
  OR3X1 U20501 ( .IN1(n18722), .IN2(n34385), .IN3(n18748), .Q(n18723) );
  NAND2X0 U20502 ( .IN1(n18723), .IN2(n18733), .QN(n18724) );
  NOR2X0 U20503 ( .IN1(n18900), .IN2(\s1/msel/gnt_p2 [1]), .QN(n29972) );
  OA22X1 U20504 ( .IN1(n18725), .IN2(n18724), .IN3(n29972), .IN4(n34385), .Q(
        n18727) );
  INVX0 U20505 ( .INP(n18895), .ZN(n29997) );
  NAND2X0 U20506 ( .IN1(n18897), .IN2(n18906), .QN(n18732) );
  OA21X1 U20507 ( .IN1(n34385), .IN2(n18732), .IN3(n18731), .Q(n18735) );
  OA21X1 U20508 ( .IN1(n29997), .IN2(n18735), .IN3(n29996), .Q(n18737) );
  NAND2X0 U20509 ( .IN1(\s1/msel/gnt_p2 [1]), .IN2(\s1/msel/gnt_p2 [0]), .QN(
        n18749) );
  NOR3X0 U20510 ( .IN1(n18737), .IN2(n18730), .IN3(n18749), .QN(n18726) );
  AO221X1 U20511 ( .IN1(n18729), .IN2(n18728), .IN3(n29974), .IN4(n18727), 
        .IN5(n18726), .Q(n18742) );
  AND2X1 U20512 ( .IN1(n18731), .IN2(n18730), .Q(n18734) );
  OA22X1 U20513 ( .IN1(n18735), .IN2(n18734), .IN3(n18733), .IN4(n18732), .Q(
        n18736) );
  OA22X1 U20514 ( .IN1(n18737), .IN2(n29974), .IN3(n29997), .IN4(n18736), .Q(
        n18740) );
  OR3X1 U20515 ( .IN1(n34445), .IN2(n18748), .IN3(n18738), .Q(n18739) );
  NAND2X0 U20516 ( .IN1(n18740), .IN2(n18739), .QN(n18741) );
  MUX21X1 U20517 ( .IN1(n18742), .IN2(n18741), .S(\s1/msel/gnt_p2 [2]), .Q(
        n18746) );
  OA221X1 U20518 ( .IN1(\s1/msel/gnt_p2 [0]), .IN2(\s1/msel/gnt_p2 [2]), .IN3(
        \s1/msel/gnt_p2 [0]), .IN4(n18910), .IN5(n18746), .Q(n18745) );
  INVX0 U20519 ( .INP(n29996), .ZN(n18743) );
  NAND2X0 U20520 ( .IN1(\s1/msel/gnt_p2 [1]), .IN2(n18894), .QN(n29968) );
  OA21X1 U20521 ( .IN1(\s1/msel/gnt_p2 [1]), .IN2(n18743), .IN3(n29968), .Q(
        n18908) );
  AND3X1 U20522 ( .IN1(\s1/msel/gnt_p2 [2]), .IN2(\s1/msel/gnt_p2 [0]), .IN3(
        n18908), .Q(n18744) );
  NOR2X0 U20523 ( .IN1(n18745), .IN2(n18744), .QN(n18754) );
  NAND3X0 U20524 ( .IN1(\s1/msel/gnt_p2 [1]), .IN2(n18746), .IN3(n18897), .QN(
        n18751) );
  INVX0 U20525 ( .INP(n18905), .ZN(n18896) );
  NAND2X0 U20526 ( .IN1(\s1/msel/gnt_p2 [0]), .IN2(n18896), .QN(n18893) );
  INVX0 U20527 ( .INP(n18746), .ZN(n18747) );
  AO221X1 U20528 ( .IN1(n18893), .IN2(n18748), .IN3(n18893), .IN4(n18747), 
        .IN5(\s1/msel/gnt_p2 [1]), .Q(n18750) );
  OR2X1 U20529 ( .IN1(n29989), .IN2(n18749), .Q(n18901) );
  NAND3X0 U20530 ( .IN1(n18751), .IN2(n18750), .IN3(n18901), .QN(n18752) );
  NAND2X0 U20531 ( .IN1(n34437), .IN2(n18752), .QN(n18753) );
  NAND2X0 U20532 ( .IN1(n18754), .IN2(n18753), .QN(n17994) );
  NAND3X0 U20533 ( .IN1(m0s14_cyc), .IN2(n34367), .IN3(n34604), .QN(n33577) );
  INVX0 U20534 ( .INP(n33577), .ZN(n33600) );
  NAND3X0 U20535 ( .IN1(m1s14_cyc), .IN2(n34334), .IN3(n34512), .QN(n33557) );
  INVX0 U20536 ( .INP(n33557), .ZN(n33560) );
  MUX21X1 U20537 ( .IN1(n33600), .IN2(n33560), .S(\s14/msel/gnt_p3 [0]), .Q(
        n33548) );
  NOR2X0 U20538 ( .IN1(n13745), .IN2(n18755), .QN(n33566) );
  NOR2X0 U20539 ( .IN1(\s14/msel/gnt_p3 [0]), .IN2(n34447), .QN(n33579) );
  NOR2X0 U20540 ( .IN1(\s14/msel/gnt_p3 [1]), .IN2(n34468), .QN(n33554) );
  INVX0 U20541 ( .INP(n33566), .ZN(n33573) );
  NOR2X0 U20542 ( .IN1(n13797), .IN2(n18756), .QN(n33601) );
  INVX0 U20543 ( .INP(n33601), .ZN(n33595) );
  NAND2X0 U20544 ( .IN1(n33573), .IN2(n33595), .QN(n33545) );
  AO22X1 U20545 ( .IN1(n33566), .IN2(n33579), .IN3(n33554), .IN4(n33545), .Q(
        n18763) );
  NAND2X0 U20546 ( .IN1(n33577), .IN2(n33557), .QN(n21764) );
  NAND2X0 U20547 ( .IN1(\s14/msel/gnt_p3 [0]), .IN2(\s14/msel/gnt_p3 [1]), 
        .QN(n33587) );
  NOR2X0 U20548 ( .IN1(n21764), .IN2(n33587), .QN(n18759) );
  NAND3X0 U20549 ( .IN1(m7s14_cyc), .IN2(n34358), .IN3(n34513), .QN(n33556) );
  NAND3X0 U20550 ( .IN1(m6s14_cyc), .IN2(n34357), .IN3(n34544), .QN(n33584) );
  NAND2X0 U20551 ( .IN1(n33556), .IN2(n33584), .QN(n21762) );
  NOR2X0 U20552 ( .IN1(n13641), .IN2(n18757), .QN(n33564) );
  NAND2X0 U20553 ( .IN1(m4s14_cyc), .IN2(n34571), .QN(n18758) );
  NOR2X0 U20554 ( .IN1(n13693), .IN2(n18758), .QN(n33589) );
  NOR2X0 U20555 ( .IN1(n33564), .IN2(n33589), .QN(n21763) );
  OA21X1 U20556 ( .IN1(n18759), .IN2(n21762), .IN3(n21763), .Q(n18760) );
  NOR2X0 U20557 ( .IN1(\s14/msel/gnt_p3 [0]), .IN2(\s14/msel/gnt_p3 [1]), .QN(
        n33593) );
  AO21X1 U20558 ( .IN1(\s14/msel/gnt_p3 [1]), .IN2(n21763), .IN3(n33545), .Q(
        n18767) );
  INVX0 U20559 ( .INP(n33593), .ZN(n33567) );
  OA222X1 U20560 ( .IN1(n18760), .IN2(n33593), .IN3(n18760), .IN4(n18767), 
        .IN5(n33567), .IN6(n33557), .Q(n18761) );
  NOR3X0 U20561 ( .IN1(\s14/msel/gnt_p3 [2]), .IN2(n18763), .IN3(n18761), .QN(
        n18776) );
  INVX0 U20562 ( .INP(n33556), .ZN(n33582) );
  AO22X1 U20563 ( .IN1(n33582), .IN2(n33579), .IN3(n33554), .IN4(n21762), .Q(
        n18762) );
  NOR2X0 U20564 ( .IN1(n34281), .IN2(n18762), .QN(n18775) );
  INVX0 U20565 ( .INP(n21764), .ZN(n18772) );
  NOR2X0 U20566 ( .IN1(\s14/msel/gnt_p3 [0]), .IN2(n33564), .QN(n33555) );
  OA221X1 U20567 ( .IN1(n21762), .IN2(n33601), .IN3(n21762), .IN4(n18772), 
        .IN5(n33555), .Q(n18771) );
  INVX0 U20568 ( .INP(n33587), .ZN(n33572) );
  NAND2X0 U20569 ( .IN1(n33555), .IN2(n33566), .QN(n18765) );
  NAND2X0 U20570 ( .IN1(n33579), .IN2(n33601), .QN(n18777) );
  INVX0 U20571 ( .INP(n18763), .ZN(n18764) );
  NAND3X0 U20572 ( .IN1(n18765), .IN2(n18777), .IN3(n18764), .QN(n18766) );
  NOR2X0 U20573 ( .IN1(n33572), .IN2(n18766), .QN(n18769) );
  NAND2X0 U20574 ( .IN1(n18772), .IN2(n18767), .QN(n18768) );
  NOR2X0 U20575 ( .IN1(n18769), .IN2(n18768), .QN(n18770) );
  NOR2X0 U20576 ( .IN1(n18771), .IN2(n18770), .QN(n18774) );
  NAND3X0 U20577 ( .IN1(n18772), .IN2(n33579), .IN3(n21763), .QN(n18773) );
  OA221X1 U20578 ( .IN1(n18776), .IN2(n18775), .IN3(n18776), .IN4(n18774), 
        .IN5(n18773), .Q(n18781) );
  NOR2X0 U20579 ( .IN1(n33548), .IN2(n18781), .QN(n18779) );
  NAND2X0 U20580 ( .IN1(n33566), .IN2(n33572), .QN(n33602) );
  NAND2X0 U20581 ( .IN1(n33602), .IN2(n18777), .QN(n18778) );
  NOR2X0 U20582 ( .IN1(n18779), .IN2(n18778), .QN(n18780) );
  OA22X1 U20583 ( .IN1(\s14/msel/gnt_p3 [2]), .IN2(n18780), .IN3(n34447), 
        .IN4(n18781), .Q(n18785) );
  NAND2X0 U20584 ( .IN1(\s14/msel/gnt_p3 [1]), .IN2(n33582), .QN(n33538) );
  OA21X1 U20585 ( .IN1(n33564), .IN2(n18781), .IN3(n33538), .Q(n18783) );
  INVX0 U20586 ( .INP(n33584), .ZN(n33578) );
  NAND2X0 U20587 ( .IN1(\s14/msel/gnt_p3 [1]), .IN2(n33578), .QN(n33539) );
  OA21X1 U20588 ( .IN1(n33589), .IN2(n18781), .IN3(n33539), .Q(n18782) );
  AO221X1 U20589 ( .IN1(\s14/msel/gnt_p3 [0]), .IN2(n18783), .IN3(n34468), 
        .IN4(n18782), .IN5(n34281), .Q(n18784) );
  NAND2X0 U20590 ( .IN1(n18785), .IN2(n18784), .QN(n17640) );
  NAND3X0 U20591 ( .IN1(n13695), .IN2(n13669), .IN3(m4s8_cyc), .QN(n32036) );
  NAND3X0 U20592 ( .IN1(n13591), .IN2(n13565), .IN3(m6s8_cyc), .QN(n18878) );
  MUX21X1 U20593 ( .IN1(n32036), .IN2(n18878), .S(\s8/msel/gnt_p0 [1]), .Q(
        n18889) );
  NAND3X0 U20594 ( .IN1(n13916), .IN2(n13877), .IN3(m0s8_cyc), .QN(n18873) );
  INVX0 U20595 ( .INP(n18873), .ZN(n18885) );
  NAND3X0 U20596 ( .IN1(n13799), .IN2(n13773), .IN3(m2s8_cyc), .QN(n18880) );
  INVX0 U20597 ( .INP(n18880), .ZN(n18875) );
  NOR2X0 U20598 ( .IN1(n18885), .IN2(n18875), .QN(n18786) );
  NAND3X0 U20599 ( .IN1(n13747), .IN2(n13721), .IN3(m3s8_cyc), .QN(n18879) );
  INVX0 U20600 ( .INP(n18879), .ZN(n32019) );
  NAND2X0 U20601 ( .IN1(n18786), .IN2(n32019), .QN(n18791) );
  INVX0 U20602 ( .INP(n18791), .ZN(n18790) );
  NAND3X0 U20603 ( .IN1(\s8/msel/gnt_p0 [0]), .IN2(n18786), .IN3(n32036), .QN(
        n18787) );
  NAND3X0 U20604 ( .IN1(n13851), .IN2(n13825), .IN3(m1s8_cyc), .QN(n18872) );
  NAND3X0 U20605 ( .IN1(n13539), .IN2(n13489), .IN3(m7s8_cyc), .QN(n32022) );
  OA21X1 U20606 ( .IN1(n18885), .IN2(n18872), .IN3(n32022), .Q(n18797) );
  NAND2X0 U20607 ( .IN1(n18787), .IN2(n18797), .QN(n18789) );
  NOR2X0 U20608 ( .IN1(\s8/msel/gnt_p0 [0]), .IN2(n34654), .QN(n32042) );
  INVX0 U20609 ( .INP(n18878), .ZN(n32043) );
  NAND2X0 U20610 ( .IN1(\s8/msel/gnt_p0 [0]), .IN2(n34654), .QN(n18788) );
  NOR2X0 U20611 ( .IN1(n32043), .IN2(n18788), .QN(n32023) );
  OA22X1 U20612 ( .IN1(n18790), .IN2(n18789), .IN3(n32042), .IN4(n32023), .Q(
        n18811) );
  NAND3X0 U20613 ( .IN1(n13643), .IN2(n13617), .IN3(m5s8_cyc), .QN(n32038) );
  OA21X1 U20614 ( .IN1(n32043), .IN2(n18797), .IN3(n32038), .Q(n18805) );
  OR2X1 U20615 ( .IN1(\s8/msel/gnt_p0 [0]), .IN2(\s8/msel/gnt_p0 [1]), .Q(
        n32031) );
  AO221X1 U20616 ( .IN1(n18805), .IN2(n32043), .IN3(n18805), .IN4(n18791), 
        .IN5(n32031), .Q(n18796) );
  INVX0 U20617 ( .INP(n32036), .ZN(n18792) );
  NOR2X0 U20618 ( .IN1(n32043), .IN2(n18792), .QN(n18798) );
  AND2X1 U20619 ( .IN1(\s8/msel/gnt_p0 [0]), .IN2(n18798), .Q(n18794) );
  NOR2X0 U20620 ( .IN1(n32038), .IN2(n18792), .QN(n18793) );
  OR2X1 U20621 ( .IN1(n32019), .IN2(n18793), .Q(n18801) );
  INVX0 U20622 ( .INP(n18872), .ZN(n18884) );
  AO221X1 U20623 ( .IN1(n18880), .IN2(n18794), .IN3(n18880), .IN4(n18801), 
        .IN5(n18884), .Q(n18802) );
  NAND3X0 U20624 ( .IN1(\s8/msel/gnt_p0 [1]), .IN2(n18802), .IN3(n18873), .QN(
        n18795) );
  NAND3X0 U20625 ( .IN1(\s8/msel/gnt_p0 [2]), .IN2(n18796), .IN3(n18795), .QN(
        n18810) );
  INVX0 U20626 ( .INP(n18797), .ZN(n18799) );
  OA221X1 U20627 ( .IN1(n18799), .IN2(\s8/msel/gnt_p0 [0]), .IN3(n18799), 
        .IN4(n18873), .IN5(n18798), .Q(n18800) );
  NOR2X0 U20628 ( .IN1(n18801), .IN2(n18800), .QN(n18804) );
  INVX0 U20629 ( .INP(n18802), .ZN(n18803) );
  OA22X1 U20630 ( .IN1(n18875), .IN2(n18804), .IN3(n18803), .IN4(n32031), .Q(
        n18808) );
  INVX0 U20631 ( .INP(n18805), .ZN(n18806) );
  NAND4X0 U20632 ( .IN1(\s8/msel/gnt_p0 [1]), .IN2(\s8/msel/gnt_p0 [0]), .IN3(
        n18806), .IN4(n32036), .QN(n18807) );
  NAND2X0 U20633 ( .IN1(n18808), .IN2(n18807), .QN(n18809) );
  OA22X1 U20634 ( .IN1(n18811), .IN2(n18810), .IN3(\s8/msel/gnt_p0 [2]), .IN4(
        n18809), .Q(n18815) );
  OA221X1 U20635 ( .IN1(\s8/msel/gnt_p0 [0]), .IN2(\s8/msel/gnt_p0 [2]), .IN3(
        \s8/msel/gnt_p0 [0]), .IN4(n18889), .IN5(n18815), .Q(n18813) );
  NAND2X0 U20636 ( .IN1(\s8/msel/gnt_p0 [1]), .IN2(n32022), .QN(n32026) );
  NAND2X0 U20637 ( .IN1(n34654), .IN2(n32038), .QN(n18886) );
  AND4X1 U20638 ( .IN1(\s8/msel/gnt_p0 [2]), .IN2(\s8/msel/gnt_p0 [0]), .IN3(
        n32026), .IN4(n18886), .Q(n18812) );
  NOR2X0 U20639 ( .IN1(n18813), .IN2(n18812), .QN(n18818) );
  OA221X1 U20640 ( .IN1(\s8/msel/gnt_p0 [1]), .IN2(n18884), .IN3(n34654), 
        .IN4(n32019), .IN5(\s8/msel/gnt_p0 [0]), .Q(n18814) );
  AO221X1 U20641 ( .IN1(n18815), .IN2(\s8/msel/gnt_p0 [1]), .IN3(n18815), 
        .IN4(n18873), .IN5(n18814), .Q(n18816) );
  NAND2X0 U20642 ( .IN1(n34403), .IN2(n18816), .QN(n18817) );
  NAND2X0 U20643 ( .IN1(n18818), .IN2(n18817), .QN(n17801) );
  NAND2X0 U20644 ( .IN1(m6s11_cyc), .IN2(n34570), .QN(n18819) );
  NOR2X0 U20645 ( .IN1(n13594), .IN2(n18819), .QN(n32749) );
  NAND3X0 U20646 ( .IN1(m7s11_cyc), .IN2(n34324), .IN3(n34539), .QN(n32760) );
  INVX0 U20647 ( .INP(n32749), .ZN(n32730) );
  NAND2X0 U20648 ( .IN1(n32760), .IN2(n32730), .QN(n18828) );
  NAND2X0 U20649 ( .IN1(m0s11_cyc), .IN2(n34584), .QN(n18820) );
  NOR2X0 U20650 ( .IN1(n13922), .IN2(n18820), .QN(n32733) );
  NOR2X0 U20651 ( .IN1(n32733), .IN2(n34419), .QN(n32747) );
  NAND3X0 U20652 ( .IN1(m1s11_cyc), .IN2(n34326), .IN3(n34537), .QN(n32746) );
  NAND2X0 U20653 ( .IN1(m5s11_cyc), .IN2(n34585), .QN(n18821) );
  NOR2X0 U20654 ( .IN1(n13646), .IN2(n18821), .QN(n32778) );
  NAND2X0 U20655 ( .IN1(m4s11_cyc), .IN2(n34569), .QN(n18822) );
  NOR2X0 U20656 ( .IN1(n13698), .IN2(n18822), .QN(n32736) );
  NOR2X0 U20657 ( .IN1(n32778), .IN2(n32736), .QN(n32723) );
  OA221X1 U20658 ( .IN1(n18828), .IN2(n32747), .IN3(n18828), .IN4(n32746), 
        .IN5(n32723), .Q(n18832) );
  NAND3X0 U20659 ( .IN1(m3s11_cyc), .IN2(n34365), .IN3(n34601), .QN(n32739) );
  NAND3X0 U20660 ( .IN1(m2s11_cyc), .IN2(n34325), .IN3(n34538), .QN(n32771) );
  NAND2X0 U20661 ( .IN1(n32739), .IN2(n32771), .QN(n32717) );
  NAND2X0 U20662 ( .IN1(\s11/msel/gnt_p3 [0]), .IN2(\s11/msel/gnt_p3 [1]), 
        .QN(n18835) );
  AO21X1 U20663 ( .IN1(n32717), .IN2(n18835), .IN3(\s11/msel/gnt_p3 [2]), .Q(
        n32724) );
  NOR2X0 U20664 ( .IN1(\s11/msel/gnt_p3 [0]), .IN2(n34419), .QN(n18823) );
  NOR2X0 U20665 ( .IN1(\s11/msel/gnt_p3 [1]), .IN2(n34399), .QN(n32774) );
  NOR2X0 U20666 ( .IN1(n18823), .IN2(n32774), .QN(n32763) );
  INVX0 U20667 ( .INP(n32760), .ZN(n32777) );
  NOR2X0 U20668 ( .IN1(\s11/msel/gnt_p3 [1]), .IN2(n32730), .QN(n32762) );
  NOR2X0 U20669 ( .IN1(n32777), .IN2(n32762), .QN(n32721) );
  INVX0 U20670 ( .INP(n32736), .ZN(n32756) );
  NAND2X0 U20671 ( .IN1(n18823), .IN2(n32756), .QN(n18826) );
  AND2X1 U20672 ( .IN1(n32723), .IN2(\s11/msel/gnt_p3 [1]), .Q(n18824) );
  OAI22X1 U20673 ( .IN1(\s11/msel/gnt_p3 [1]), .IN2(\s11/msel/gnt_p3 [0]), 
        .IN3(n32717), .IN4(n18824), .QN(n18825) );
  OA221X1 U20674 ( .IN1(n32778), .IN2(n32739), .IN3(n32778), .IN4(n18826), 
        .IN5(n18825), .Q(n18827) );
  INVX0 U20675 ( .INP(n32733), .ZN(n32772) );
  NAND2X0 U20676 ( .IN1(n32746), .IN2(n32772), .QN(n32716) );
  OA22X1 U20677 ( .IN1(n32763), .IN2(n32721), .IN3(n18827), .IN4(n32716), .Q(
        n18830) );
  INVX0 U20678 ( .INP(n18828), .ZN(n32722) );
  INVX0 U20679 ( .INP(n32778), .ZN(n32741) );
  NAND2X0 U20680 ( .IN1(n34399), .IN2(n32741), .QN(n32755) );
  AO221X1 U20681 ( .IN1(n32722), .IN2(n32771), .IN3(n32722), .IN4(n32716), 
        .IN5(n32755), .Q(n18829) );
  NAND3X0 U20682 ( .IN1(\s11/msel/gnt_p3 [2]), .IN2(n18830), .IN3(n18829), 
        .QN(n18831) );
  OA21X1 U20683 ( .IN1(n18832), .IN2(n32724), .IN3(n18831), .Q(n18838) );
  AO22X1 U20684 ( .IN1(\s11/msel/gnt_p3 [1]), .IN2(n32749), .IN3(n18838), 
        .IN4(n32756), .Q(n18834) );
  AO22X1 U20685 ( .IN1(\s11/msel/gnt_p3 [1]), .IN2(n32777), .IN3(n18838), 
        .IN4(n32741), .Q(n18833) );
  OA221X1 U20686 ( .IN1(\s11/msel/gnt_p3 [0]), .IN2(n18834), .IN3(n34399), 
        .IN4(n18833), .IN5(\s11/msel/gnt_p3 [2]), .Q(n18837) );
  NOR2X0 U20687 ( .IN1(n32739), .IN2(n18835), .QN(n32784) );
  OA21X1 U20688 ( .IN1(\s11/msel/gnt_p3 [0]), .IN2(n32772), .IN3(n32746), .Q(
        n32725) );
  OA221X1 U20689 ( .IN1(n32784), .IN2(n18838), .IN3(n32784), .IN4(n32725), 
        .IN5(n34444), .Q(n18836) );
  NOR2X0 U20690 ( .IN1(n18837), .IN2(n18836), .QN(n18840) );
  NAND2X0 U20691 ( .IN1(n18838), .IN2(\s11/msel/gnt_p3 [1]), .QN(n18839) );
  NAND2X0 U20692 ( .IN1(n18840), .IN2(n18839), .QN(n17724) );
  INVX0 U20693 ( .INP(n18842), .ZN(n18866) );
  INVX0 U20694 ( .INP(n18843), .ZN(n18857) );
  NAND2X0 U20695 ( .IN1(n18841), .IN2(n33631), .QN(n18851) );
  INVX0 U20696 ( .INP(n33631), .ZN(n18859) );
  OA21X1 U20697 ( .IN1(n18859), .IN2(n33632), .IN3(n33625), .Q(n18850) );
  OA21X1 U20698 ( .IN1(n34394), .IN2(n18851), .IN3(n18850), .Q(n18854) );
  OA21X1 U20699 ( .IN1(n18857), .IN2(n18854), .IN3(n18864), .Q(n18855) );
  OR3X1 U20700 ( .IN1(n34242), .IN2(n18866), .IN3(n18855), .Q(n18849) );
  INVX0 U20701 ( .INP(n18841), .ZN(n33635) );
  NAND2X0 U20702 ( .IN1(n18843), .IN2(n18842), .QN(n18846) );
  OR2X1 U20703 ( .IN1(n18859), .IN2(n34394), .Q(n18845) );
  OA21X1 U20704 ( .IN1(n18866), .IN2(n18864), .IN3(n18844), .Q(n18852) );
  OA221X1 U20705 ( .IN1(n18846), .IN2(n33625), .IN3(n18846), .IN4(n18845), 
        .IN5(n18852), .Q(n18847) );
  OA21X1 U20706 ( .IN1(n33635), .IN2(n18852), .IN3(n33632), .Q(n18858) );
  NAND2X0 U20707 ( .IN1(n34394), .IN2(n34242), .QN(n33616) );
  OA22X1 U20708 ( .IN1(n33635), .IN2(n18847), .IN3(n18858), .IN4(n33616), .Q(
        n18848) );
  NAND3X0 U20709 ( .IN1(n18849), .IN2(n18848), .IN3(\s14/msel/gnt_p1 [2]), 
        .QN(n18863) );
  AND2X1 U20710 ( .IN1(n18866), .IN2(n18850), .Q(n18853) );
  OA22X1 U20711 ( .IN1(n18854), .IN2(n18853), .IN3(n18852), .IN4(n18851), .Q(
        n18856) );
  OA22X1 U20712 ( .IN1(n18857), .IN2(n18856), .IN3(n18855), .IN4(n33616), .Q(
        n18861) );
  OR4X1 U20713 ( .IN1(n34242), .IN2(n34394), .IN3(n18859), .IN4(n18858), .Q(
        n18860) );
  NAND3X0 U20714 ( .IN1(n18861), .IN2(n34386), .IN3(n18860), .QN(n18862) );
  NAND2X0 U20715 ( .IN1(n18863), .IN2(n18862), .QN(n18867) );
  AO221X1 U20716 ( .IN1(\s14/msel/gnt_p1 [1]), .IN2(n33625), .IN3(n34242), 
        .IN4(n18864), .IN5(n34394), .Q(n18865) );
  OA221X1 U20717 ( .IN1(n18867), .IN2(n18866), .IN3(n18867), .IN4(n34242), 
        .IN5(n18865), .Q(n18869) );
  OA22X1 U20718 ( .IN1(\s14/msel/gnt_p1 [2]), .IN2(n18869), .IN3(n18868), 
        .IN4(n18867), .Q(n18871) );
  NAND2X0 U20719 ( .IN1(n18871), .IN2(n18870), .QN(n17636) );
  OA21X1 U20720 ( .IN1(\s8/msel/gnt_p0 [0]), .IN2(n18873), .IN3(n18872), .Q(
        n32035) );
  NOR2X0 U20721 ( .IN1(n32035), .IN2(\s8/msel/gnt_p0 [1]), .QN(n18883) );
  NOR2X0 U20722 ( .IN1(n18879), .IN2(n34654), .QN(n18874) );
  NOR2X0 U20723 ( .IN1(\s8/msel/gnt_p0 [2]), .IN2(n18874), .QN(n18877) );
  NAND2X0 U20724 ( .IN1(n18875), .IN2(n32042), .QN(n18876) );
  NAND2X0 U20725 ( .IN1(n18877), .IN2(n18876), .QN(n32034) );
  AND2X1 U20726 ( .IN1(n32038), .IN2(n32036), .Q(n32025) );
  NAND2X0 U20727 ( .IN1(n18878), .IN2(n32022), .QN(n32030) );
  INVX0 U20728 ( .INP(n32030), .ZN(n18881) );
  NAND2X0 U20729 ( .IN1(n18880), .IN2(n18879), .QN(n32028) );
  AO22X1 U20730 ( .IN1(n32025), .IN2(n18881), .IN3(n34654), .IN4(n32028), .Q(
        n18882) );
  NOR2X0 U20731 ( .IN1(n18885), .IN2(n18884), .QN(n32027) );
  INVX0 U20732 ( .INP(n32027), .ZN(n18890) );
  INVX0 U20733 ( .INP(n32026), .ZN(n18888) );
  NOR2X0 U20734 ( .IN1(n18886), .IN2(n32030), .QN(n18887) );
  OAI222X1 U20735 ( .IN1(n18890), .IN2(n32028), .IN3(\s8/msel/gnt_p0 [0]), 
        .IN4(n18889), .IN5(n18888), .IN6(n18887), .QN(n18891) );
  NAND2X0 U20736 ( .IN1(\s8/msel/gnt_p0 [2]), .IN2(n18891), .QN(n18892) );
  NAND2X0 U20737 ( .IN1(n18197), .IN2(n18892), .QN(n17803) );
  OA21X1 U20738 ( .IN1(\s1/msel/gnt_p2 [0]), .IN2(n18906), .IN3(n18893), .Q(
        n30003) );
  NOR2X0 U20739 ( .IN1(\s1/msel/gnt_p2 [1]), .IN2(n30003), .QN(n18904) );
  NAND2X0 U20740 ( .IN1(n18895), .IN2(n18894), .QN(n29970) );
  NAND2X0 U20741 ( .IN1(n29996), .IN2(n29999), .QN(n29983) );
  NOR2X0 U20742 ( .IN1(n29970), .IN2(n29983), .QN(n34080) );
  NOR2X0 U20743 ( .IN1(\s1/msel/gnt_p2 [1]), .IN2(n34385), .QN(n29981) );
  NOR2X0 U20744 ( .IN1(n18896), .IN2(n29974), .QN(n29980) );
  NAND2X0 U20745 ( .IN1(n18897), .IN2(n29989), .QN(n18907) );
  INVX0 U20746 ( .INP(n18907), .ZN(n29979) );
  OA21X1 U20747 ( .IN1(n29981), .IN2(n29980), .IN3(n29979), .Q(n18899) );
  AND2X1 U20748 ( .IN1(\s1/msel/gnt_p2 [1]), .IN2(n29989), .Q(n18898) );
  NOR2X0 U20749 ( .IN1(n18899), .IN2(n18898), .QN(n18903) );
  NOR2X0 U20750 ( .IN1(\s1/msel/gnt_p2 [0]), .IN2(n34445), .QN(n29998) );
  NAND2X0 U20751 ( .IN1(n29998), .IN2(n18900), .QN(n18902) );
  NAND3X0 U20752 ( .IN1(n18902), .IN2(n18901), .IN3(n34437), .QN(n30004) );
  NAND2X0 U20753 ( .IN1(n18906), .IN2(n18905), .QN(n29971) );
  NOR2X0 U20754 ( .IN1(n29971), .IN2(n18907), .QN(n34081) );
  NOR2X0 U20755 ( .IN1(n18908), .IN2(n34081), .QN(n18913) );
  NAND2X0 U20756 ( .IN1(n34445), .IN2(n29970), .QN(n18909) );
  NAND2X0 U20757 ( .IN1(\s1/msel/gnt_p2 [0]), .IN2(n18909), .QN(n29969) );
  NAND2X0 U20758 ( .IN1(n18910), .IN2(n18909), .QN(n18911) );
  NAND2X0 U20759 ( .IN1(n29969), .IN2(n18911), .QN(n18912) );
  NAND2X0 U20760 ( .IN1(n18913), .IN2(n18912), .QN(n18914) );
  NAND2X0 U20761 ( .IN1(\s1/msel/gnt_p2 [2]), .IN2(n18914), .QN(n18915) );
  NAND2X0 U20762 ( .IN1(n18194), .IN2(n18915), .QN(n17996) );
  NAND3X0 U20763 ( .IN1(n13594), .IN2(m6s11_cyc), .IN3(n34570), .QN(n18935) );
  INVX0 U20764 ( .INP(n18935), .ZN(n18956) );
  NAND2X0 U20765 ( .IN1(\s11/msel/gnt_p2 [1]), .IN2(n18956), .QN(n32927) );
  AND2X1 U20766 ( .IN1(n32927), .IN2(\s11/msel/gnt_p2 [2]), .Q(n18987) );
  NAND3X0 U20767 ( .IN1(n13698), .IN2(m4s11_cyc), .IN3(n34569), .QN(n18962) );
  INVX0 U20768 ( .INP(n18962), .ZN(n18988) );
  NAND2X0 U20769 ( .IN1(n18988), .IN2(n34407), .QN(n32928) );
  NOR2X0 U20770 ( .IN1(\s11/msel/gnt_p2 [0]), .IN2(\s11/msel/gnt_p2 [1]), .QN(
        n18929) );
  NAND3X0 U20771 ( .IN1(n13802), .IN2(m2s11_cyc), .IN3(n34538), .QN(n18979) );
  NAND3X0 U20772 ( .IN1(n13542), .IN2(m7s11_cyc), .IN3(n34539), .QN(n18989) );
  INVX0 U20773 ( .INP(n18989), .ZN(n18955) );
  NOR2X0 U20774 ( .IN1(n18956), .IN2(n18988), .QN(n18920) );
  NAND3X0 U20775 ( .IN1(n18979), .IN2(n18955), .IN3(n18920), .QN(n18918) );
  INVX0 U20776 ( .INP(n18979), .ZN(n18957) );
  INVX0 U20777 ( .INP(n18920), .ZN(n18919) );
  AND3X1 U20778 ( .IN1(n13750), .IN2(m3s11_cyc), .IN3(n34601), .Q(n32937) );
  NAND3X0 U20779 ( .IN1(n13646), .IN2(m5s11_cyc), .IN3(n34585), .QN(n18969) );
  NOR2X0 U20780 ( .IN1(n18988), .IN2(n18969), .QN(n18916) );
  NOR2X0 U20781 ( .IN1(n32937), .IN2(n18916), .QN(n18921) );
  OA21X1 U20782 ( .IN1(n34470), .IN2(n18919), .IN3(n18921), .Q(n18917) );
  NAND3X0 U20783 ( .IN1(n13854), .IN2(m1s11_cyc), .IN3(n34537), .QN(n18953) );
  OA21X1 U20784 ( .IN1(n18957), .IN2(n18917), .IN3(n18953), .Q(n18938) );
  NAND2X0 U20785 ( .IN1(n18918), .IN2(n18938), .QN(n18928) );
  INVX0 U20786 ( .INP(n18929), .ZN(n18971) );
  NAND3X0 U20787 ( .IN1(n13922), .IN2(m0s11_cyc), .IN3(n34584), .QN(n18954) );
  INVX0 U20788 ( .INP(n18954), .ZN(n18985) );
  OA21X1 U20789 ( .IN1(n18985), .IN2(n18953), .IN3(n18989), .Q(n18933) );
  NOR2X0 U20790 ( .IN1(n18933), .IN2(n18919), .QN(n18924) );
  NAND3X0 U20791 ( .IN1(n18920), .IN2(\s11/msel/gnt_p2 [0]), .IN3(n18954), 
        .QN(n18922) );
  NAND2X0 U20792 ( .IN1(n18922), .IN2(n18921), .QN(n18923) );
  NOR2X0 U20793 ( .IN1(\s11/msel/gnt_p2 [1]), .IN2(n18957), .QN(n18961) );
  OA22X1 U20794 ( .IN1(n18924), .IN2(n18923), .IN3(n18961), .IN4(n34470), .Q(
        n18927) );
  NOR2X0 U20795 ( .IN1(n18957), .IN2(n18985), .QN(n18930) );
  NAND2X0 U20796 ( .IN1(\s11/msel/gnt_p2 [0]), .IN2(n18930), .QN(n18925) );
  OA221X1 U20797 ( .IN1(n18956), .IN2(n18933), .IN3(n18956), .IN4(n18925), 
        .IN5(n18969), .Q(n18937) );
  NAND2X0 U20798 ( .IN1(\s11/msel/gnt_p2 [0]), .IN2(\s11/msel/gnt_p2 [1]), 
        .QN(n18990) );
  NOR3X0 U20799 ( .IN1(n18937), .IN2(n18988), .IN3(n18990), .QN(n18926) );
  AO221X1 U20800 ( .IN1(n18929), .IN2(n18928), .IN3(n18971), .IN4(n18927), 
        .IN5(n18926), .Q(n18943) );
  NAND2X0 U20801 ( .IN1(n32937), .IN2(n18930), .QN(n18934) );
  NAND2X0 U20802 ( .IN1(n18969), .IN2(n34470), .QN(n18931) );
  NAND3X0 U20803 ( .IN1(n18931), .IN2(n18962), .IN3(n18930), .QN(n18932) );
  NAND3X0 U20804 ( .IN1(n18934), .IN2(n18933), .IN3(n18932), .QN(n18936) );
  NAND2X0 U20805 ( .IN1(\s11/msel/gnt_p2 [1]), .IN2(n34470), .QN(n18980) );
  NAND2X0 U20806 ( .IN1(n18935), .IN2(n34407), .QN(n18967) );
  NAND2X0 U20807 ( .IN1(n18980), .IN2(n18967), .QN(n18965) );
  NAND2X0 U20808 ( .IN1(n18936), .IN2(n18965), .QN(n18941) );
  OR2X1 U20809 ( .IN1(n18971), .IN2(n18937), .Q(n18940) );
  OR3X1 U20810 ( .IN1(n34407), .IN2(n18985), .IN3(n18938), .Q(n18939) );
  NAND4X0 U20811 ( .IN1(\s11/msel/gnt_p2 [2]), .IN2(n18941), .IN3(n18940), 
        .IN4(n18939), .QN(n18942) );
  OA21X1 U20812 ( .IN1(\s11/msel/gnt_p2 [2]), .IN2(n18943), .IN3(n18942), .Q(
        n18945) );
  OA221X1 U20813 ( .IN1(\s11/msel/gnt_p2 [0]), .IN2(n18987), .IN3(
        \s11/msel/gnt_p2 [0]), .IN4(n32928), .IN5(n18945), .Q(n18944) );
  MUX21X1 U20814 ( .IN1(n18969), .IN2(n18989), .S(\s11/msel/gnt_p2 [1]), .Q(
        n32929) );
  NAND2X0 U20815 ( .IN1(\s11/msel/gnt_p2 [2]), .IN2(\s11/msel/gnt_p2 [0]), 
        .QN(n18986) );
  NOR2X0 U20816 ( .IN1(n32929), .IN2(n18986), .QN(n32926) );
  NOR2X0 U20817 ( .IN1(n18944), .IN2(n32926), .QN(n18952) );
  INVX0 U20818 ( .INP(n18990), .ZN(n18963) );
  NAND2X0 U20819 ( .IN1(n32937), .IN2(n18963), .QN(n18981) );
  NAND3X0 U20820 ( .IN1(\s11/msel/gnt_p2 [1]), .IN2(n18945), .IN3(n18979), 
        .QN(n18949) );
  INVX0 U20821 ( .INP(n18953), .ZN(n18984) );
  NAND2X0 U20822 ( .IN1(\s11/msel/gnt_p2 [0]), .IN2(n18984), .QN(n18947) );
  INVX0 U20823 ( .INP(n18945), .ZN(n18946) );
  AO221X1 U20824 ( .IN1(n18947), .IN2(n18985), .IN3(n18947), .IN4(n18946), 
        .IN5(\s11/msel/gnt_p2 [1]), .Q(n18948) );
  NAND3X0 U20825 ( .IN1(n18981), .IN2(n18949), .IN3(n18948), .QN(n18950) );
  NAND2X0 U20826 ( .IN1(n34401), .IN2(n18950), .QN(n18951) );
  NAND2X0 U20827 ( .IN1(n18952), .IN2(n18951), .QN(n17714) );
  INVX0 U20828 ( .INP(n18969), .ZN(n18978) );
  NAND2X0 U20829 ( .IN1(n18954), .IN2(n18953), .QN(n34172) );
  NAND2X0 U20830 ( .IN1(n18969), .IN2(n18962), .QN(n32933) );
  NOR2X0 U20831 ( .IN1(n34172), .IN2(n32933), .QN(n18968) );
  NOR2X0 U20832 ( .IN1(n18956), .IN2(n18955), .QN(n32935) );
  NOR2X0 U20833 ( .IN1(n32935), .IN2(n32933), .QN(n18958) );
  NOR3X0 U20834 ( .IN1(n32937), .IN2(n18968), .IN3(n18958), .QN(n18960) );
  OR2X1 U20835 ( .IN1(\s11/msel/gnt_p2 [1]), .IN2(n18984), .Q(n32936) );
  NOR2X0 U20836 ( .IN1(n32937), .IN2(n18957), .QN(n18964) );
  INVX0 U20837 ( .INP(n18964), .ZN(n34171) );
  NOR2X0 U20838 ( .IN1(n18958), .IN2(n34171), .QN(n18959) );
  OA22X1 U20839 ( .IN1(n18960), .IN2(n18980), .IN3(n32936), .IN4(n18959), .Q(
        n18977) );
  OAI21X1 U20840 ( .IN1(n18961), .IN2(n34172), .IN3(n32935), .QN(n18970) );
  NAND4X0 U20841 ( .IN1(n18963), .IN2(n18962), .IN3(n18969), .IN4(n18970), 
        .QN(n18976) );
  NOR2X0 U20842 ( .IN1(n18964), .IN2(n34172), .QN(n18974) );
  NAND2X0 U20843 ( .IN1(n18989), .IN2(n18965), .QN(n18966) );
  AO22X1 U20844 ( .IN1(n18968), .IN2(n18967), .IN3(n18990), .IN4(n18966), .Q(
        n18973) );
  OA21X1 U20845 ( .IN1(n18974), .IN2(n18970), .IN3(n18969), .Q(n18972) );
  OAI22X1 U20846 ( .IN1(n18974), .IN2(n18973), .IN3(n18972), .IN4(n18971), 
        .QN(n18975) );
  OA222X1 U20847 ( .IN1(\s11/msel/gnt_p2 [2]), .IN2(n18977), .IN3(
        \s11/msel/gnt_p2 [2]), .IN4(n18976), .IN5(n18975), .IN6(n34401), .Q(
        n18994) );
  AO221X1 U20848 ( .IN1(n34407), .IN2(n18978), .IN3(n34407), .IN4(n18986), 
        .IN5(n18994), .Q(n18996) );
  NOR2X0 U20849 ( .IN1(n18980), .IN2(n18979), .QN(n18983) );
  NAND2X0 U20850 ( .IN1(n18981), .IN2(n34401), .QN(n18982) );
  NOR2X0 U20851 ( .IN1(n18983), .IN2(n18982), .QN(n32940) );
  MUX21X1 U20852 ( .IN1(n18985), .IN2(n18984), .S(\s11/msel/gnt_p2 [0]), .Q(
        n32932) );
  INVX0 U20853 ( .INP(n18986), .ZN(n18992) );
  OA21X1 U20854 ( .IN1(n18988), .IN2(n18994), .IN3(n18987), .Q(n18991) );
  OA22X1 U20855 ( .IN1(n18992), .IN2(n18991), .IN3(n18990), .IN4(n18989), .Q(
        n18993) );
  AO221X1 U20856 ( .IN1(n32940), .IN2(n18994), .IN3(n32940), .IN4(n32932), 
        .IN5(n18993), .Q(n18995) );
  NAND2X0 U20857 ( .IN1(n18996), .IN2(n18995), .QN(n17715) );
  NAND3X0 U20858 ( .IN1(n13525), .IN2(n13469), .IN3(m7s6_cyc), .QN(n31504) );
  NAND2X0 U20859 ( .IN1(\s6/msel/gnt_p0 [1]), .IN2(n31504), .QN(n18998) );
  NAND3X0 U20860 ( .IN1(n13629), .IN2(n13603), .IN3(m5s6_cyc), .QN(n31530) );
  NAND2X0 U20861 ( .IN1(n34675), .IN2(n31530), .QN(n18997) );
  AND4X1 U20862 ( .IN1(\s6/msel/gnt_p0 [2]), .IN2(\s6/msel/gnt_p0 [0]), .IN3(
        n18998), .IN4(n18997), .Q(n19146) );
  NAND3X0 U20863 ( .IN1(n13577), .IN2(n13551), .IN3(m6s6_cyc), .QN(n31505) );
  INVX0 U20864 ( .INP(n31505), .ZN(n31535) );
  INVX0 U20865 ( .INP(n31504), .ZN(n19117) );
  NOR2X0 U20866 ( .IN1(n31535), .IN2(n19117), .QN(n31511) );
  INVX0 U20867 ( .INP(n31511), .ZN(n18999) );
  NAND3X0 U20868 ( .IN1(n13681), .IN2(n13655), .IN3(m4s6_cyc), .QN(n31512) );
  NAND2X0 U20869 ( .IN1(n31530), .IN2(n31512), .QN(n31506) );
  NOR2X0 U20870 ( .IN1(n18999), .IN2(n31506), .QN(n19006) );
  NAND3X0 U20871 ( .IN1(n13733), .IN2(n13707), .IN3(m3s6_cyc), .QN(n19148) );
  INVX0 U20872 ( .INP(n19148), .ZN(n31509) );
  AND3X1 U20873 ( .IN1(n13785), .IN2(n13759), .IN3(m2s6_cyc), .Q(n19137) );
  NOR2X0 U20874 ( .IN1(n31509), .IN2(n19137), .QN(n31507) );
  NAND3X0 U20875 ( .IN1(n13837), .IN2(n13811), .IN3(m1s6_cyc), .QN(n19149) );
  AND2X1 U20876 ( .IN1(n34675), .IN2(n19149), .Q(n31508) );
  NAND2X0 U20877 ( .IN1(n31507), .IN2(n31508), .QN(n19000) );
  AND2X1 U20878 ( .IN1(n19000), .IN2(n34675), .Q(n19005) );
  NAND3X0 U20879 ( .IN1(n13892), .IN2(n13863), .IN3(m0s6_cyc), .QN(n19151) );
  MUX21X1 U20880 ( .IN1(n19151), .IN2(n19149), .S(\s6/msel/gnt_p0 [0]), .Q(
        n31528) );
  NOR2X0 U20881 ( .IN1(\s6/msel/gnt_p0 [1]), .IN2(n31528), .QN(n19004) );
  NOR2X0 U20882 ( .IN1(n19148), .IN2(n34675), .QN(n19001) );
  NOR2X0 U20883 ( .IN1(\s6/msel/gnt_p0 [2]), .IN2(n19001), .QN(n19003) );
  NOR2X0 U20884 ( .IN1(\s6/msel/gnt_p0 [0]), .IN2(n34675), .QN(n31534) );
  NAND2X0 U20885 ( .IN1(n19137), .IN2(n31534), .QN(n19002) );
  NAND2X0 U20886 ( .IN1(n19003), .IN2(n19002), .QN(n31527) );
  NOR4X0 U20887 ( .IN1(n19006), .IN2(n19005), .IN3(n19004), .IN4(n31527), .QN(
        n19007) );
  NOR2X0 U20888 ( .IN1(n19146), .IN2(n19007), .QN(n19012) );
  NAND2X0 U20889 ( .IN1(n31530), .IN2(n31511), .QN(n19009) );
  NOR2X0 U20890 ( .IN1(n31535), .IN2(n34671), .QN(n19120) );
  OAI21X1 U20891 ( .IN1(\s6/msel/gnt_p0 [1]), .IN2(n19120), .IN3(n31504), .QN(
        n31520) );
  MUX21X1 U20892 ( .IN1(n31512), .IN2(n31505), .S(\s6/msel/gnt_p0 [1]), .Q(
        n19145) );
  INVX0 U20893 ( .INP(n19145), .ZN(n19008) );
  NAND2X0 U20894 ( .IN1(n19151), .IN2(n19149), .QN(n31510) );
  INVX0 U20895 ( .INP(n31510), .ZN(n31519) );
  AO222X1 U20896 ( .IN1(n19009), .IN2(n31520), .IN3(n34671), .IN4(n19008), 
        .IN5(n31507), .IN6(n31519), .Q(n19010) );
  NAND2X0 U20897 ( .IN1(\s6/msel/gnt_p0 [2]), .IN2(n19010), .QN(n19011) );
  NAND2X0 U20898 ( .IN1(n19012), .IN2(n19011), .QN(n17859) );
  NAND3X0 U20899 ( .IN1(m0s15_cyc), .IN2(n13876), .IN3(n34298), .QN(n33871) );
  NOR2X0 U20900 ( .IN1(\s15/msel/gnt_p1 [1]), .IN2(n33871), .QN(n19029) );
  NAND3X0 U20901 ( .IN1(m6s15_cyc), .IN2(n13564), .IN3(n34360), .QN(n21757) );
  INVX0 U20902 ( .INP(n21757), .ZN(n33897) );
  INVX0 U20903 ( .INP(n33871), .ZN(n19016) );
  NAND3X0 U20904 ( .IN1(m1s15_cyc), .IN2(n13824), .IN3(n34302), .QN(n33870) );
  NAND3X0 U20905 ( .IN1(m7s15_cyc), .IN2(n13485), .IN3(n34301), .QN(n21756) );
  OA21X1 U20906 ( .IN1(n19016), .IN2(n33870), .IN3(n21756), .Q(n19017) );
  NAND3X0 U20907 ( .IN1(m5s15_cyc), .IN2(n13616), .IN3(n34300), .QN(n33895) );
  OA21X1 U20908 ( .IN1(n33897), .IN2(n19017), .IN3(n33895), .Q(n19020) );
  NAND3X0 U20909 ( .IN1(m4s15_cyc), .IN2(n13668), .IN3(n34299), .QN(n33880) );
  INVX0 U20910 ( .INP(n33880), .ZN(n33894) );
  NAND3X0 U20911 ( .IN1(m3s15_cyc), .IN2(n13720), .IN3(n34303), .QN(n33888) );
  OA21X1 U20912 ( .IN1(n33894), .IN2(n33895), .IN3(n33888), .Q(n19019) );
  NAND3X0 U20913 ( .IN1(m2s15_cyc), .IN2(n13772), .IN3(n34359), .QN(n33889) );
  INVX0 U20914 ( .INP(n33889), .ZN(n33868) );
  AO221X1 U20915 ( .IN1(n19019), .IN2(n33894), .IN3(n19019), .IN4(n34272), 
        .IN5(n33868), .Q(n19013) );
  OA21X1 U20916 ( .IN1(n19016), .IN2(n19013), .IN3(n19017), .Q(n19014) );
  OA22X1 U20917 ( .IN1(\s15/msel/gnt_p1 [1]), .IN2(n19020), .IN3(n33897), 
        .IN4(n19014), .Q(n19027) );
  OA21X1 U20918 ( .IN1(n33868), .IN2(n19019), .IN3(n33870), .Q(n19015) );
  OR3X1 U20919 ( .IN1(n34412), .IN2(n19016), .IN3(n19015), .Q(n19026) );
  NOR2X0 U20920 ( .IN1(n19015), .IN2(\s15/msel/gnt_p1 [1]), .QN(n19024) );
  AO221X1 U20921 ( .IN1(n19017), .IN2(n19016), .IN3(n19017), .IN4(n34272), 
        .IN5(n33894), .Q(n19018) );
  AO221X1 U20922 ( .IN1(n19019), .IN2(n33897), .IN3(n19019), .IN4(n19018), 
        .IN5(n33868), .Q(n19022) );
  OR4X1 U20923 ( .IN1(n34412), .IN2(n34272), .IN3(n33894), .IN4(n19020), .Q(
        n19021) );
  NAND2X0 U20924 ( .IN1(n19022), .IN2(n19021), .QN(n19023) );
  NOR2X0 U20925 ( .IN1(n19024), .IN2(n19023), .QN(n19025) );
  OA222X1 U20926 ( .IN1(n34448), .IN2(n19027), .IN3(n34448), .IN4(n19026), 
        .IN5(n19025), .IN6(\s15/msel/gnt_p1 [2]), .Q(n19030) );
  NAND2X0 U20927 ( .IN1(\s15/msel/gnt_p1 [0]), .IN2(\s15/msel/gnt_p1 [1]), 
        .QN(n19028) );
  OA22X1 U20928 ( .IN1(n19029), .IN2(n19030), .IN3(n19028), .IN4(n33888), .Q(
        n19032) );
  MUX21X1 U20929 ( .IN1(n33894), .IN2(n33897), .S(\s15/msel/gnt_p1 [1]), .Q(
        n33863) );
  OA21X1 U20930 ( .IN1(n34448), .IN2(n33863), .IN3(n34272), .Q(n19031) );
  OA22X1 U20931 ( .IN1(\s15/msel/gnt_p1 [2]), .IN2(n19032), .IN3(n19031), 
        .IN4(n19030), .Q(n19034) );
  INVX0 U20932 ( .INP(n33895), .ZN(n19033) );
  NAND2X0 U20933 ( .IN1(\s15/msel/gnt_p1 [1]), .IN2(n21756), .QN(n33886) );
  OA21X1 U20934 ( .IN1(\s15/msel/gnt_p1 [1]), .IN2(n19033), .IN3(n33886), .Q(
        n33864) );
  NAND3X0 U20935 ( .IN1(\s15/msel/gnt_p1 [0]), .IN2(\s15/msel/gnt_p1 [2]), 
        .IN3(n33864), .QN(n33877) );
  NAND2X0 U20936 ( .IN1(n19034), .IN2(n33877), .QN(n17608) );
  NAND3X0 U20937 ( .IN1(m5s8_cyc), .IN2(n34588), .IN3(n34239), .QN(n31961) );
  NAND2X0 U20938 ( .IN1(m7s8_cyc), .IN2(n34592), .QN(n19035) );
  NOR2X0 U20939 ( .IN1(n13539), .IN2(n19035), .QN(n31958) );
  NAND2X0 U20940 ( .IN1(\s8/msel/gnt_p3 [1]), .IN2(n31958), .QN(n31976) );
  OA21X1 U20941 ( .IN1(\s8/msel/gnt_p3 [1]), .IN2(n31961), .IN3(n31976), .Q(
        n31943) );
  NAND2X0 U20942 ( .IN1(\s8/msel/gnt_p3 [0]), .IN2(n34223), .QN(n19037) );
  NAND2X0 U20943 ( .IN1(m1s8_cyc), .IN2(n34593), .QN(n19036) );
  NOR2X0 U20944 ( .IN1(n13851), .IN2(n19036), .QN(n31945) );
  INVX0 U20945 ( .INP(n31945), .ZN(n19042) );
  NOR2X0 U20946 ( .IN1(n19037), .IN2(n19042), .QN(n19070) );
  NAND2X0 U20947 ( .IN1(m2s8_cyc), .IN2(n34591), .QN(n19038) );
  NOR2X0 U20948 ( .IN1(n13799), .IN2(n19038), .QN(n31955) );
  NAND2X0 U20949 ( .IN1(m0s8_cyc), .IN2(n34589), .QN(n19039) );
  NOR2X0 U20950 ( .IN1(n13916), .IN2(n19039), .QN(n31946) );
  INVX0 U20951 ( .INP(n31961), .ZN(n31977) );
  NAND2X0 U20952 ( .IN1(n34223), .IN2(n31977), .QN(n19049) );
  NOR2X0 U20953 ( .IN1(n34228), .IN2(n34223), .QN(n31944) );
  INVX0 U20954 ( .INP(n31944), .ZN(n19067) );
  NAND3X0 U20955 ( .IN1(m4s8_cyc), .IN2(n34238), .IN3(n34369), .QN(n31948) );
  INVX0 U20956 ( .INP(n31948), .ZN(n31975) );
  AO21X1 U20957 ( .IN1(n34228), .IN2(n31961), .IN3(n31975), .Q(n19043) );
  NAND2X0 U20958 ( .IN1(m6s8_cyc), .IN2(n34580), .QN(n19040) );
  NOR2X0 U20959 ( .IN1(n13591), .IN2(n19040), .QN(n31973) );
  NAND2X0 U20960 ( .IN1(m3s8_cyc), .IN2(n34590), .QN(n19041) );
  NOR2X0 U20961 ( .IN1(n13747), .IN2(n19041), .QN(n31962) );
  INVX0 U20962 ( .INP(n31962), .ZN(n31949) );
  OA221X1 U20963 ( .IN1(n19043), .IN2(n31973), .IN3(n19043), .IN4(n31961), 
        .IN5(n31949), .Q(n19052) );
  OA21X1 U20964 ( .IN1(n31955), .IN2(n19052), .IN3(n19042), .Q(n19054) );
  OR3X1 U20965 ( .IN1(n19067), .IN2(n31946), .IN3(n19054), .Q(n19048) );
  INVX0 U20966 ( .INP(n31958), .ZN(n19050) );
  OA21X1 U20967 ( .IN1(n31946), .IN2(n19042), .IN3(n19050), .Q(n19056) );
  NOR2X0 U20968 ( .IN1(n31955), .IN2(n31946), .QN(n19045) );
  NAND2X0 U20969 ( .IN1(n31949), .IN2(n19043), .QN(n19044) );
  NAND2X0 U20970 ( .IN1(n19045), .IN2(n19044), .QN(n19046) );
  AO21X1 U20971 ( .IN1(n19056), .IN2(n19046), .IN3(n31973), .Q(n19047) );
  NAND4X0 U20972 ( .IN1(\s8/msel/gnt_p3 [2]), .IN2(n19049), .IN3(n19048), 
        .IN4(n19047), .QN(n19066) );
  AND3X1 U20973 ( .IN1(n31946), .IN2(n31949), .IN3(n31961), .Q(n19051) );
  OR2X1 U20974 ( .IN1(n31975), .IN2(n31973), .Q(n19057) );
  OA22X1 U20975 ( .IN1(n19052), .IN2(n19051), .IN3(n19050), .IN4(n19057), .Q(
        n19055) );
  NAND2X0 U20976 ( .IN1(n34228), .IN2(n34223), .QN(n19053) );
  OA22X1 U20977 ( .IN1(n31955), .IN2(n19055), .IN3(n19054), .IN4(n19053), .Q(
        n19064) );
  NOR2X0 U20978 ( .IN1(n31975), .IN2(n19067), .QN(n19060) );
  NOR2X0 U20979 ( .IN1(n19057), .IN2(n19056), .QN(n19061) );
  INVX0 U20980 ( .INP(n19061), .ZN(n19058) );
  NAND2X0 U20981 ( .IN1(n31961), .IN2(n19058), .QN(n19059) );
  NAND2X0 U20982 ( .IN1(n19060), .IN2(n19059), .QN(n19063) );
  NAND2X0 U20983 ( .IN1(\s8/msel/gnt_p3 [1]), .IN2(n19061), .QN(n19062) );
  NAND4X0 U20984 ( .IN1(n19064), .IN2(n34456), .IN3(n19063), .IN4(n19062), 
        .QN(n19065) );
  NAND2X0 U20985 ( .IN1(n19066), .IN2(n19065), .QN(n19072) );
  AO221X1 U20986 ( .IN1(\s8/msel/gnt_p3 [1]), .IN2(n31955), .IN3(n34223), 
        .IN4(n31946), .IN5(n19072), .Q(n19068) );
  OA21X1 U20987 ( .IN1(n31949), .IN2(n19067), .IN3(n34456), .Q(n31971) );
  NAND2X0 U20988 ( .IN1(n19068), .IN2(n31971), .QN(n19069) );
  NOR2X0 U20989 ( .IN1(n19070), .IN2(n19069), .QN(n19071) );
  AO221X1 U20990 ( .IN1(\s8/msel/gnt_p3 [2]), .IN2(n31943), .IN3(
        \s8/msel/gnt_p3 [2]), .IN4(n34228), .IN5(n19071), .Q(n19074) );
  MUX21X1 U20991 ( .IN1(n31975), .IN2(n31973), .S(\s8/msel/gnt_p3 [1]), .Q(
        n31940) );
  AO221X1 U20992 ( .IN1(n34228), .IN2(n34456), .IN3(n34228), .IN4(n31940), 
        .IN5(n19072), .Q(n19073) );
  NAND2X0 U20993 ( .IN1(n19074), .IN2(n19073), .QN(n17807) );
  INVX0 U20994 ( .INP(n19075), .ZN(n30423) );
  NOR2X0 U20995 ( .IN1(n19078), .IN2(n30423), .QN(n19110) );
  INVX0 U20996 ( .INP(n19091), .ZN(n19105) );
  OA21X1 U20997 ( .IN1(n30446), .IN2(n19079), .IN3(n19076), .Q(n19095) );
  OA21X1 U20998 ( .IN1(n19106), .IN2(n19095), .IN3(n19078), .Q(n19099) );
  OR3X1 U20999 ( .IN1(n34388), .IN2(n19105), .IN3(n19099), .Q(n19086) );
  NAND2X0 U21000 ( .IN1(n19077), .IN2(n19091), .QN(n19081) );
  NOR2X0 U21001 ( .IN1(n19105), .IN2(n19078), .QN(n19089) );
  NOR2X0 U21002 ( .IN1(n30440), .IN2(n19089), .QN(n19080) );
  OA21X1 U21003 ( .IN1(n34658), .IN2(n19081), .IN3(n19080), .Q(n19083) );
  OA21X1 U21004 ( .IN1(n30442), .IN2(n19083), .IN3(n19079), .Q(n19087) );
  AND2X1 U21005 ( .IN1(n19080), .IN2(n30446), .Q(n19082) );
  OA22X1 U21006 ( .IN1(n19083), .IN2(n19082), .IN3(n19095), .IN4(n19081), .Q(
        n19084) );
  OA22X1 U21007 ( .IN1(n19087), .IN2(n30430), .IN3(n30442), .IN4(n19084), .Q(
        n19085) );
  NAND3X0 U21008 ( .IN1(n19086), .IN2(n19085), .IN3(\s3/msel/gnt_p1 [2]), .QN(
        n19104) );
  OR3X1 U21009 ( .IN1(n34388), .IN2(n19087), .IN3(n30446), .Q(n19102) );
  NOR2X0 U21010 ( .IN1(n30442), .IN2(n30446), .QN(n19088) );
  NAND2X0 U21011 ( .IN1(n30440), .IN2(n19088), .QN(n19098) );
  NAND3X0 U21012 ( .IN1(n19089), .IN2(n19092), .IN3(n19090), .QN(n19094) );
  NAND4X0 U21013 ( .IN1(\s3/msel/gnt_p1 [0]), .IN2(n19092), .IN3(n19091), 
        .IN4(n19090), .QN(n19093) );
  NAND4X0 U21014 ( .IN1(n19095), .IN2(n19098), .IN3(n19094), .IN4(n19093), 
        .QN(n19096) );
  NAND2X0 U21015 ( .IN1(n19097), .IN2(n19096), .QN(n19101) );
  AO221X1 U21016 ( .IN1(n19099), .IN2(n19106), .IN3(n19099), .IN4(n19098), 
        .IN5(n30430), .Q(n19100) );
  NAND4X0 U21017 ( .IN1(n34418), .IN2(n19102), .IN3(n19101), .IN4(n19100), 
        .QN(n19103) );
  NAND2X0 U21018 ( .IN1(n19104), .IN2(n19103), .QN(n19112) );
  AO221X1 U21019 ( .IN1(\s3/msel/gnt_p1 [1]), .IN2(n19106), .IN3(n34388), 
        .IN4(n19105), .IN5(n19112), .Q(n19107) );
  NAND2X0 U21020 ( .IN1(n19108), .IN2(n19107), .QN(n19109) );
  NOR2X0 U21021 ( .IN1(n19110), .IN2(n19109), .QN(n19114) );
  OA21X1 U21022 ( .IN1(n19111), .IN2(n34418), .IN3(n34658), .Q(n19113) );
  OA22X1 U21023 ( .IN1(\s3/msel/gnt_p1 [2]), .IN2(n19114), .IN3(n19113), .IN4(
        n19112), .Q(n19116) );
  NAND2X0 U21024 ( .IN1(n19116), .IN2(n19115), .QN(n17944) );
  INVX0 U21025 ( .INP(n19151), .ZN(n19130) );
  NOR2X0 U21026 ( .IN1(n19149), .IN2(n19130), .QN(n19131) );
  NOR2X0 U21027 ( .IN1(n19117), .IN2(n19131), .QN(n19122) );
  INVX0 U21028 ( .INP(n19122), .ZN(n19119) );
  NOR2X0 U21029 ( .IN1(n19130), .IN2(n19137), .QN(n19125) );
  OA221X1 U21030 ( .IN1(n31509), .IN2(\s6/msel/gnt_p0 [0]), .IN3(n31509), 
        .IN4(n31512), .IN5(n19125), .Q(n19118) );
  OA22X1 U21031 ( .IN1(n31534), .IN2(n19120), .IN3(n19119), .IN4(n19118), .Q(
        n19144) );
  NAND2X0 U21032 ( .IN1(n31505), .IN2(n31512), .QN(n19129) );
  OR2X1 U21033 ( .IN1(n34671), .IN2(n19129), .Q(n19121) );
  INVX0 U21034 ( .INP(n31512), .ZN(n19138) );
  NOR2X0 U21035 ( .IN1(n31530), .IN2(n19138), .QN(n19124) );
  NOR2X0 U21036 ( .IN1(n31509), .IN2(n19124), .QN(n19134) );
  OA221X1 U21037 ( .IN1(n19137), .IN2(n19121), .IN3(n19137), .IN4(n19134), 
        .IN5(n19149), .Q(n19135) );
  OR3X1 U21038 ( .IN1(n34675), .IN2(n19130), .IN3(n19135), .Q(n19128) );
  OA21X1 U21039 ( .IN1(n31535), .IN2(n19122), .IN3(n31530), .Q(n19139) );
  NAND2X0 U21040 ( .IN1(n31509), .IN2(n19125), .QN(n19123) );
  NAND2X0 U21041 ( .IN1(n34671), .IN2(n34675), .QN(n31516) );
  AO221X1 U21042 ( .IN1(n19139), .IN2(n31535), .IN3(n19139), .IN4(n19123), 
        .IN5(n31516), .Q(n19127) );
  NAND2X0 U21043 ( .IN1(n19125), .IN2(n19124), .QN(n19126) );
  NAND4X0 U21044 ( .IN1(\s6/msel/gnt_p0 [2]), .IN2(n19128), .IN3(n19127), 
        .IN4(n19126), .QN(n19143) );
  AO221X1 U21045 ( .IN1(n31504), .IN2(n19130), .IN3(n31504), .IN4(n34671), 
        .IN5(n19129), .Q(n19133) );
  NOR2X0 U21046 ( .IN1(\s6/msel/gnt_p0 [0]), .IN2(n19138), .QN(n31529) );
  NAND3X0 U21047 ( .IN1(n19131), .IN2(n31505), .IN3(n31529), .QN(n19132) );
  AND3X1 U21048 ( .IN1(n19134), .IN2(n19133), .IN3(n19132), .Q(n19136) );
  OA22X1 U21049 ( .IN1(n19137), .IN2(n19136), .IN3(n19135), .IN4(n31516), .Q(
        n19141) );
  OR4X1 U21050 ( .IN1(n34675), .IN2(n34671), .IN3(n19139), .IN4(n19138), .Q(
        n19140) );
  NAND2X0 U21051 ( .IN1(n19141), .IN2(n19140), .QN(n19142) );
  OA22X1 U21052 ( .IN1(n19144), .IN2(n19143), .IN3(\s6/msel/gnt_p0 [2]), .IN4(
        n19142), .Q(n19152) );
  OA221X1 U21053 ( .IN1(\s6/msel/gnt_p0 [0]), .IN2(\s6/msel/gnt_p0 [2]), .IN3(
        \s6/msel/gnt_p0 [0]), .IN4(n19145), .IN5(n19152), .Q(n19147) );
  NOR2X0 U21054 ( .IN1(n19147), .IN2(n19146), .QN(n19155) );
  AOI221X1 U21055 ( .IN1(n34675), .IN2(n19149), .IN3(\s6/msel/gnt_p0 [1]), 
        .IN4(n19148), .IN5(n34671), .QN(n19150) );
  AO221X1 U21056 ( .IN1(n19152), .IN2(\s6/msel/gnt_p0 [1]), .IN3(n19152), 
        .IN4(n19151), .IN5(n19150), .Q(n19153) );
  NAND2X0 U21057 ( .IN1(n34402), .IN2(n19153), .QN(n19154) );
  NAND2X0 U21058 ( .IN1(n19155), .IN2(n19154), .QN(n17857) );
  NAND3X0 U21059 ( .IN1(n13743), .IN2(m3s12_cyc), .IN3(n34507), .QN(n33209) );
  NAND2X0 U21060 ( .IN1(\s12/msel/gnt_p2 [0]), .IN2(\s12/msel/gnt_p2 [1]), 
        .QN(n33190) );
  NOR2X0 U21061 ( .IN1(n33209), .IN2(n33190), .QN(n33195) );
  NAND3X0 U21062 ( .IN1(n13908), .IN2(m0s12_cyc), .IN3(n34509), .QN(n33184) );
  NAND3X0 U21063 ( .IN1(n13587), .IN2(m6s12_cyc), .IN3(n34540), .QN(n33220) );
  INVX0 U21064 ( .INP(n33220), .ZN(n19168) );
  INVX0 U21065 ( .INP(n33184), .ZN(n33192) );
  NAND3X0 U21066 ( .IN1(n13847), .IN2(m1s12_cyc), .IN3(n34508), .QN(n33191) );
  OR2X1 U21067 ( .IN1(n34474), .IN2(n19156), .Q(n33219) );
  OA21X1 U21068 ( .IN1(n33192), .IN2(n33191), .IN3(n33219), .Q(n19160) );
  NAND3X0 U21069 ( .IN1(n13639), .IN2(m5s12_cyc), .IN3(n34506), .QN(n33227) );
  OA21X1 U21070 ( .IN1(n19168), .IN2(n19160), .IN3(n33227), .Q(n19166) );
  NAND2X0 U21071 ( .IN1(n34244), .IN2(n34422), .QN(n33222) );
  NOR2X0 U21072 ( .IN1(n19166), .IN2(n33222), .QN(n19164) );
  NAND3X0 U21073 ( .IN1(n13795), .IN2(m2s12_cyc), .IN3(n34541), .QN(n33183) );
  INVX0 U21074 ( .INP(n33183), .ZN(n33197) );
  NOR2X0 U21075 ( .IN1(n34475), .IN2(n19157), .QN(n19169) );
  OA21X1 U21076 ( .IN1(n19169), .IN2(n33227), .IN3(n33209), .Q(n19167) );
  INVX0 U21077 ( .INP(n19169), .ZN(n33230) );
  NAND3X0 U21078 ( .IN1(\s12/msel/gnt_p2 [0]), .IN2(n33230), .IN3(n33220), 
        .QN(n19158) );
  OA221X1 U21079 ( .IN1(n33197), .IN2(n19167), .IN3(n33197), .IN4(n19158), 
        .IN5(n33191), .Q(n19165) );
  NOR3X0 U21080 ( .IN1(n33192), .IN2(n19165), .IN3(n33190), .QN(n19163) );
  NOR2X0 U21081 ( .IN1(\s12/msel/gnt_p2 [0]), .IN2(n34422), .QN(n33196) );
  OA21X1 U21082 ( .IN1(n19169), .IN2(n34244), .IN3(n19167), .Q(n19159) );
  NOR3X0 U21083 ( .IN1(n33197), .IN2(n33192), .IN3(n19159), .QN(n19161) );
  INVX0 U21084 ( .INP(n19160), .ZN(n19171) );
  OA22X1 U21085 ( .IN1(n33220), .IN2(n33196), .IN3(n19161), .IN4(n19171), .Q(
        n19162) );
  NOR4X0 U21086 ( .IN1(n19164), .IN2(n19163), .IN3(n19162), .IN4(n34553), .QN(
        n19178) );
  NOR2X0 U21087 ( .IN1(n19165), .IN2(n33222), .QN(n19176) );
  NOR3X0 U21088 ( .IN1(n19169), .IN2(n19166), .IN3(n33190), .QN(n19175) );
  INVX0 U21089 ( .INP(n19167), .ZN(n19173) );
  NOR2X0 U21090 ( .IN1(n19169), .IN2(n19168), .QN(n19170) );
  OA221X1 U21091 ( .IN1(n19171), .IN2(\s12/msel/gnt_p2 [0]), .IN3(n19171), 
        .IN4(n33184), .IN5(n19170), .Q(n19172) );
  OA21X1 U21092 ( .IN1(n19173), .IN2(n19172), .IN3(n33183), .Q(n19174) );
  NOR4X0 U21093 ( .IN1(\s12/msel/gnt_p2 [2]), .IN2(n19176), .IN3(n19175), 
        .IN4(n19174), .QN(n19177) );
  NOR2X0 U21094 ( .IN1(n19178), .IN2(n19177), .QN(n19181) );
  OA21X1 U21095 ( .IN1(\s12/msel/gnt_p2 [1]), .IN2(n33184), .IN3(n19181), .Q(
        n19180) );
  NOR3X0 U21096 ( .IN1(n34244), .IN2(n33191), .IN3(\s12/msel/gnt_p2 [1]), .QN(
        n19179) );
  NOR3X0 U21097 ( .IN1(n33195), .IN2(n19180), .IN3(n19179), .QN(n19184) );
  NOR2X0 U21098 ( .IN1(\s12/msel/gnt_p2 [1]), .IN2(n33230), .QN(n33185) );
  NOR2X0 U21099 ( .IN1(n34422), .IN2(n33220), .QN(n33186) );
  OR2X1 U21100 ( .IN1(n34553), .IN2(n33186), .Q(n33231) );
  OA21X1 U21101 ( .IN1(n33185), .IN2(n33231), .IN3(n34244), .Q(n19183) );
  INVX0 U21102 ( .INP(n19181), .ZN(n19182) );
  OA22X1 U21103 ( .IN1(\s12/msel/gnt_p2 [2]), .IN2(n19184), .IN3(n19183), 
        .IN4(n19182), .Q(n19186) );
  NAND2X0 U21104 ( .IN1(\s12/msel/gnt_p2 [1]), .IN2(n33219), .QN(n33189) );
  NAND2X0 U21105 ( .IN1(n34422), .IN2(n33227), .QN(n33188) );
  NAND4X0 U21106 ( .IN1(\s12/msel/gnt_p2 [2]), .IN2(\s12/msel/gnt_p2 [0]), 
        .IN3(n33189), .IN4(n33188), .QN(n19185) );
  NAND2X0 U21107 ( .IN1(n19186), .IN2(n19185), .QN(n17686) );
  INVX0 U21108 ( .INP(m3s0_addr[2]), .ZN(n28592) );
  INVX0 U21109 ( .INP(m7s0_addr[2]), .ZN(n28596) );
  OA22X1 U21110 ( .IN1(n23812), .IN2(n28592), .IN3(n23824), .IN4(n28596), .Q(
        n19190) );
  INVX0 U21111 ( .INP(m0s0_addr[2]), .ZN(n28591) );
  INVX0 U21112 ( .INP(m2s0_addr[2]), .ZN(n28594) );
  OA22X1 U21113 ( .IN1(n23838), .IN2(n28591), .IN3(n23837), .IN4(n28594), .Q(
        n19189) );
  INVX0 U21114 ( .INP(m4s0_addr[2]), .ZN(n28590) );
  INVX0 U21115 ( .INP(m1s0_addr[2]), .ZN(n28589) );
  OA22X1 U21116 ( .IN1(n23825), .IN2(n28590), .IN3(n23818), .IN4(n28589), .Q(
        n19188) );
  INVX0 U21117 ( .INP(m5s0_addr[2]), .ZN(n28593) );
  INVX0 U21118 ( .INP(m6s0_addr[2]), .ZN(n28595) );
  OA22X1 U21119 ( .IN1(n23826), .IN2(n28593), .IN3(n23833), .IN4(n28595), .Q(
        n19187) );
  NAND4X0 U21120 ( .IN1(n19190), .IN2(n19189), .IN3(n19188), .IN4(n19187), 
        .QN(s15_addr_o[2]) );
  INVX0 U21121 ( .INP(m5s0_addr[28]), .ZN(n28910) );
  NOR2X0 U21122 ( .IN1(m5s0_addr[29]), .IN2(n28910), .QN(n19198) );
  NOR2X0 U21123 ( .IN1(m5s0_addr[31]), .IN2(m5s0_addr[30]), .QN(n19197) );
  AND2X1 U21124 ( .IN1(n19198), .IN2(n19197), .Q(n29345) );
  INVX0 U21125 ( .INP(n29345), .ZN(n21727) );
  INVX0 U21126 ( .INP(m0s1_data_i[30]), .ZN(n22601) );
  INVX0 U21127 ( .INP(m5s0_addr[29]), .ZN(n28920) );
  NOR2X0 U21128 ( .IN1(m5s0_addr[28]), .IN2(n28920), .QN(n19201) );
  AND2X1 U21129 ( .IN1(n19197), .IN2(n19201), .Q(n29344) );
  INVX0 U21130 ( .INP(n29344), .ZN(n21742) );
  INVX0 U21131 ( .INP(m0s2_data_i[30]), .ZN(n22603) );
  OA22X1 U21132 ( .IN1(n21727), .IN2(n22601), .IN3(n21742), .IN4(n22603), .Q(
        n19194) );
  INVX0 U21133 ( .INP(m5s0_addr[31]), .ZN(n28954) );
  NOR2X0 U21134 ( .IN1(m5s0_addr[30]), .IN2(n28954), .QN(n19195) );
  NOR2X0 U21135 ( .IN1(m5s0_addr[29]), .IN2(m5s0_addr[28]), .QN(n19199) );
  AND2X1 U21136 ( .IN1(n19195), .IN2(n19199), .Q(n29338) );
  INVX0 U21137 ( .INP(n29338), .ZN(n21740) );
  INVX0 U21138 ( .INP(m0s8_data_i[30]), .ZN(n21061) );
  INVX0 U21139 ( .INP(m5s0_addr[30]), .ZN(n28936) );
  NOR2X0 U21140 ( .IN1(n28954), .IN2(n28936), .QN(n19202) );
  AND2X1 U21141 ( .IN1(n19202), .IN2(n19199), .Q(n29334) );
  INVX0 U21142 ( .INP(n29334), .ZN(n21735) );
  INVX0 U21143 ( .INP(m0s12_data_i[30]), .ZN(n22600) );
  OA22X1 U21144 ( .IN1(n21740), .IN2(n21061), .IN3(n21735), .IN4(n22600), .Q(
        n19193) );
  NOR2X0 U21145 ( .IN1(n28920), .IN2(n28910), .QN(n19196) );
  AND2X1 U21146 ( .IN1(n19196), .IN2(n19195), .Q(n29335) );
  INVX0 U21147 ( .INP(m0s11_data_i[30]), .ZN(n21062) );
  NOR2X0 U21148 ( .IN1(m5s0_addr[31]), .IN2(n28936), .QN(n19200) );
  NAND2X0 U21149 ( .IN1(n19196), .IN2(n19200), .QN(n21738) );
  INVX0 U21150 ( .INP(m0s7_data_i[30]), .ZN(n21060) );
  OA22X1 U21151 ( .IN1(n21728), .IN2(n21062), .IN3(n21738), .IN4(n21060), .Q(
        n19192) );
  NAND2X0 U21152 ( .IN1(n19198), .IN2(n19195), .QN(n21746) );
  INVX0 U21153 ( .INP(n21746), .ZN(n29337) );
  NAND2X0 U21154 ( .IN1(n29337), .IN2(m0s9_data_i[30]), .QN(n19191) );
  NAND4X0 U21155 ( .IN1(n19194), .IN2(n19193), .IN3(n19192), .IN4(n19191), 
        .QN(n19208) );
  AND2X1 U21156 ( .IN1(n19201), .IN2(n19195), .Q(n29336) );
  INVX0 U21157 ( .INP(n29336), .ZN(n21730) );
  INVX0 U21158 ( .INP(m0s10_data_i[30]), .ZN(n22598) );
  AND2X1 U21159 ( .IN1(n19196), .IN2(n19197), .Q(n29343) );
  INVX0 U21160 ( .INP(n29343), .ZN(n21744) );
  INVX0 U21161 ( .INP(m0s3_data_i[30]), .ZN(n21070) );
  OA22X1 U21162 ( .IN1(n21730), .IN2(n22598), .IN3(n21744), .IN4(n21070), .Q(
        n19206) );
  AND2X1 U21163 ( .IN1(n19202), .IN2(n19198), .Q(n29333) );
  INVX0 U21164 ( .INP(m0s13_data_i[30]), .ZN(n22602) );
  AND2X1 U21165 ( .IN1(n19197), .IN2(n19199), .Q(n29347) );
  INVX0 U21166 ( .INP(n29347), .ZN(n21724) );
  INVX0 U21167 ( .INP(m0s0_data_i[30]), .ZN(n22177) );
  OA22X1 U21168 ( .IN1(n21704), .IN2(n22602), .IN3(n21724), .IN4(n22177), .Q(
        n19205) );
  AND2X1 U21169 ( .IN1(n19198), .IN2(n19200), .Q(n29341) );
  INVX0 U21170 ( .INP(n29341), .ZN(n21736) );
  INVX0 U21171 ( .INP(m0s5_data_i[30]), .ZN(n21072) );
  AND2X1 U21172 ( .IN1(n19200), .IN2(n19201), .Q(n29340) );
  INVX0 U21173 ( .INP(n29340), .ZN(n21745) );
  INVX0 U21174 ( .INP(m0s6_data_i[30]), .ZN(n21071) );
  OA22X1 U21175 ( .IN1(n21736), .IN2(n21072), .IN3(n21745), .IN4(n21071), .Q(
        n19204) );
  AND2X1 U21176 ( .IN1(n19200), .IN2(n19199), .Q(n29342) );
  INVX0 U21177 ( .INP(n29342), .ZN(n21712) );
  INVX0 U21178 ( .INP(m0s4_data_i[30]), .ZN(n21069) );
  NAND2X0 U21179 ( .IN1(n19202), .IN2(n19201), .QN(n21726) );
  INVX0 U21180 ( .INP(m0s14_data_i[30]), .ZN(n22597) );
  OA22X1 U21181 ( .IN1(n21712), .IN2(n21069), .IN3(n21726), .IN4(n22597), .Q(
        n19203) );
  NAND4X0 U21182 ( .IN1(n19206), .IN2(n19205), .IN3(n19204), .IN4(n19203), 
        .QN(n19207) );
  NOR2X0 U21183 ( .IN1(n19208), .IN2(n19207), .QN(n19223) );
  NAND4X0 U21184 ( .IN1(m2s0_addr[29]), .IN2(m2s0_addr[28]), .IN3(
        m2s0_addr[31]), .IN4(m2s0_addr[30]), .QN(n20112) );
  NOR2X0 U21185 ( .IN1(n23837), .IN2(n20112), .QN(n20051) );
  NAND2X0 U21186 ( .IN1(m2_stb_i), .IN2(n20051), .QN(n23632) );
  NAND4X0 U21187 ( .IN1(m2s0_addr[25]), .IN2(m2s0_addr[24]), .IN3(
        m2s0_addr[27]), .IN4(m2s0_addr[26]), .QN(n19210) );
  NAND4X0 U21188 ( .IN1(m6s0_addr[29]), .IN2(m6s0_addr[28]), .IN3(
        m6s0_addr[31]), .IN4(m6s0_addr[30]), .QN(n20886) );
  NOR2X0 U21189 ( .IN1(n23799), .IN2(n20886), .QN(n23389) );
  NAND2X0 U21190 ( .IN1(m6_stb_i), .IN2(n23389), .QN(n23631) );
  NAND4X0 U21191 ( .IN1(m6s0_addr[25]), .IN2(m6s0_addr[24]), .IN3(
        m6s0_addr[27]), .IN4(m6s0_addr[26]), .QN(n19209) );
  OA22X1 U21192 ( .IN1(n23632), .IN2(n19210), .IN3(n23631), .IN4(n19209), .Q(
        n19220) );
  NAND4X0 U21193 ( .IN1(m1s0_addr[29]), .IN2(m1s0_addr[28]), .IN3(
        m1s0_addr[31]), .IN4(m1s0_addr[30]), .QN(n22217) );
  NOR2X0 U21194 ( .IN1(n23818), .IN2(n22217), .QN(n23289) );
  NAND2X0 U21195 ( .IN1(m1_stb_i), .IN2(n23289), .QN(n23628) );
  NAND4X0 U21196 ( .IN1(m1s0_addr[25]), .IN2(m1s0_addr[24]), .IN3(
        m1s0_addr[27]), .IN4(m1s0_addr[26]), .QN(n19212) );
  NAND4X0 U21197 ( .IN1(m7s0_addr[28]), .IN2(m7s0_addr[29]), .IN3(
        m7s0_addr[31]), .IN4(m7s0_addr[30]), .QN(n20454) );
  NOR2X0 U21198 ( .IN1(n23824), .IN2(n20454), .QN(n23446) );
  NAND2X0 U21199 ( .IN1(m7_stb_i), .IN2(n23446), .QN(n23627) );
  NAND4X0 U21200 ( .IN1(m7s0_addr[25]), .IN2(m7s0_addr[24]), .IN3(
        m7s0_addr[27]), .IN4(m7s0_addr[26]), .QN(n19211) );
  OA22X1 U21201 ( .IN1(n23628), .IN2(n19212), .IN3(n23627), .IN4(n19211), .Q(
        n19219) );
  NAND4X0 U21202 ( .IN1(m5s0_addr[29]), .IN2(m5s0_addr[28]), .IN3(
        m5s0_addr[31]), .IN4(m5s0_addr[30]), .QN(n21170) );
  NOR2X0 U21203 ( .IN1(n23832), .IN2(n21170), .QN(n23364) );
  NAND2X0 U21204 ( .IN1(m5_stb_i), .IN2(n23364), .QN(n23626) );
  NAND4X0 U21205 ( .IN1(m5s0_addr[25]), .IN2(m5s0_addr[24]), .IN3(
        m5s0_addr[27]), .IN4(m5s0_addr[26]), .QN(n19214) );
  NAND4X0 U21206 ( .IN1(m0s0_addr[28]), .IN2(m0s0_addr[29]), .IN3(
        m0s0_addr[31]), .IN4(m0s0_addr[30]), .QN(n22021) );
  NOR2X0 U21207 ( .IN1(n23838), .IN2(n22021), .QN(n23203) );
  NAND2X0 U21208 ( .IN1(m0_stb_i), .IN2(n23203), .QN(n23625) );
  NAND4X0 U21209 ( .IN1(m0s0_addr[25]), .IN2(m0s0_addr[24]), .IN3(
        m0s0_addr[27]), .IN4(m0s0_addr[26]), .QN(n19213) );
  OA22X1 U21210 ( .IN1(n23626), .IN2(n19214), .IN3(n23625), .IN4(n19213), .Q(
        n19218) );
  NAND4X0 U21211 ( .IN1(m3s0_addr[28]), .IN2(m3s0_addr[29]), .IN3(
        m3s0_addr[31]), .IN4(m3s0_addr[30]), .QN(n19808) );
  NOR2X0 U21212 ( .IN1(n23835), .IN2(n19808), .QN(n23314) );
  NAND2X0 U21213 ( .IN1(m3_stb_i), .IN2(n23314), .QN(n23630) );
  NAND4X0 U21214 ( .IN1(m3s0_addr[25]), .IN2(m3s0_addr[24]), .IN3(
        m3s0_addr[27]), .IN4(m3s0_addr[26]), .QN(n19216) );
  NAND4X0 U21215 ( .IN1(m4s0_addr[28]), .IN2(m4s0_addr[29]), .IN3(
        m4s0_addr[31]), .IN4(m4s0_addr[30]), .QN(n19458) );
  NOR2X0 U21216 ( .IN1(n23825), .IN2(n19458), .QN(n23339) );
  NAND2X0 U21217 ( .IN1(m4_stb_i), .IN2(n23339), .QN(n23629) );
  NAND4X0 U21218 ( .IN1(m4s0_addr[25]), .IN2(m4s0_addr[24]), .IN3(
        m4s0_addr[27]), .IN4(m4s0_addr[26]), .QN(n19215) );
  OA22X1 U21219 ( .IN1(n23630), .IN2(n19216), .IN3(n23629), .IN4(n19215), .Q(
        n19217) );
  NAND4X0 U21220 ( .IN1(n19220), .IN2(n19219), .IN3(n19218), .IN4(n19217), 
        .QN(n23451) );
  INVX0 U21221 ( .INP(n23451), .ZN(n19221) );
  OR2X1 U21222 ( .IN1(n18178), .IN2(n19221), .Q(n23445) );
  INVX0 U21223 ( .INP(n23445), .ZN(n23501) );
  NOR2X0 U21224 ( .IN1(n23501), .IN2(n21170), .QN(n21753) );
  NAND2X0 U21225 ( .IN1(s15_data_i[30]), .IN2(n21753), .QN(n19222) );
  NAND2X0 U21226 ( .IN1(n19223), .IN2(n19222), .QN(m5_data_o[30]) );
  INVX0 U21227 ( .INP(m0s7_data_i[31]), .ZN(n21090) );
  INVX0 U21228 ( .INP(n29333), .ZN(n21704) );
  INVX0 U21229 ( .INP(m0s13_data_i[31]), .ZN(n22618) );
  OA22X1 U21230 ( .IN1(n21738), .IN2(n21090), .IN3(n21704), .IN4(n22618), .Q(
        n19227) );
  INVX0 U21231 ( .INP(m0s8_data_i[31]), .ZN(n21083) );
  INVX0 U21232 ( .INP(m0s14_data_i[31]), .ZN(n21096) );
  OA22X1 U21233 ( .IN1(n21740), .IN2(n21083), .IN3(n21726), .IN4(n21096), .Q(
        n19226) );
  INVX0 U21234 ( .INP(m0s5_data_i[31]), .ZN(n22616) );
  INVX0 U21235 ( .INP(m0s0_data_i[31]), .ZN(n21107) );
  OA22X1 U21236 ( .IN1(n21736), .IN2(n22616), .IN3(n21724), .IN4(n21107), .Q(
        n19225) );
  NAND2X0 U21237 ( .IN1(n29334), .IN2(m0s12_data_i[31]), .QN(n19224) );
  NAND4X0 U21238 ( .IN1(n19227), .IN2(n19226), .IN3(n19225), .IN4(n19224), 
        .QN(n19233) );
  INVX0 U21239 ( .INP(m0s2_data_i[31]), .ZN(n22619) );
  INVX0 U21240 ( .INP(m0s6_data_i[31]), .ZN(n21081) );
  OA22X1 U21241 ( .IN1(n21742), .IN2(n22619), .IN3(n21745), .IN4(n21081), .Q(
        n19231) );
  INVX0 U21242 ( .INP(m0s10_data_i[31]), .ZN(n21088) );
  INVX0 U21243 ( .INP(m0s3_data_i[31]), .ZN(n22617) );
  OA22X1 U21244 ( .IN1(n21730), .IN2(n21088), .IN3(n21744), .IN4(n22617), .Q(
        n19230) );
  INVX0 U21245 ( .INP(m0s1_data_i[31]), .ZN(n21099) );
  INVX0 U21246 ( .INP(m0s9_data_i[31]), .ZN(n21102) );
  OA22X1 U21247 ( .IN1(n21727), .IN2(n21099), .IN3(n21746), .IN4(n21102), .Q(
        n19229) );
  INVX0 U21248 ( .INP(n29335), .ZN(n21728) );
  INVX0 U21249 ( .INP(m0s11_data_i[31]), .ZN(n21086) );
  INVX0 U21250 ( .INP(m0s4_data_i[31]), .ZN(n21105) );
  OA22X1 U21251 ( .IN1(n21728), .IN2(n21086), .IN3(n21712), .IN4(n21105), .Q(
        n19228) );
  NAND4X0 U21252 ( .IN1(n19231), .IN2(n19230), .IN3(n19229), .IN4(n19228), 
        .QN(n19232) );
  NOR2X0 U21253 ( .IN1(n19233), .IN2(n19232), .QN(n19235) );
  NAND2X0 U21254 ( .IN1(s15_data_i[31]), .IN2(n21753), .QN(n19234) );
  NAND2X0 U21255 ( .IN1(n19235), .IN2(n19234), .QN(m5_data_o[31]) );
  INVX0 U21256 ( .INP(s5_ack_i), .ZN(n21144) );
  INVX0 U21257 ( .INP(m4s0_addr[30]), .ZN(n28939) );
  NOR2X0 U21258 ( .IN1(m4s0_addr[31]), .IN2(n28939), .QN(n19242) );
  INVX0 U21259 ( .INP(m4s0_addr[28]), .ZN(n28906) );
  NOR2X0 U21260 ( .IN1(m4s0_addr[29]), .IN2(n28906), .QN(n19240) );
  AND2X1 U21261 ( .IN1(n19242), .IN2(n19240), .Q(n29322) );
  MUX41X1 U21262 ( .IN1(\s5/msel/gnt_p0 [0]), .IN3(\s5/msel/gnt_p1 [0]), .IN2(
        \s5/msel/gnt_p2 [0]), .IN4(\s5/msel/gnt_p3 [0]), .S0(
        \s5/msel/pri_out [0]), .S1(\s5/msel/pri_out [1]), .Q(n23227) );
  MUX41X1 U21263 ( .IN1(\s5/msel/gnt_p0 [2]), .IN3(\s5/msel/gnt_p1 [2]), .IN2(
        \s5/msel/gnt_p2 [2]), .IN4(\s5/msel/gnt_p3 [2]), .S0(
        \s5/msel/pri_out [0]), .S1(\s5/msel/pri_out [1]), .Q(n23133) );
  INVX0 U21264 ( .INP(n23133), .ZN(n21143) );
  MUX41X1 U21265 ( .IN1(\s5/msel/gnt_p0 [1]), .IN3(\s5/msel/gnt_p1 [1]), .IN2(
        \s5/msel/gnt_p2 [1]), .IN4(\s5/msel/gnt_p3 [1]), .S0(
        \s5/msel/pri_out [0]), .S1(\s5/msel/pri_out [1]), .Q(n23132) );
  NOR3X0 U21266 ( .IN1(n23227), .IN2(n21143), .IN3(n23132), .QN(n29063) );
  NAND2X0 U21267 ( .IN1(n29322), .IN2(n29063), .QN(n26584) );
  INVX0 U21268 ( .INP(s1_ack_i), .ZN(n21138) );
  NOR2X0 U21269 ( .IN1(m4s0_addr[31]), .IN2(m4s0_addr[30]), .QN(n19245) );
  AND2X1 U21270 ( .IN1(n19245), .IN2(n19240), .Q(n29326) );
  MUX41X1 U21271 ( .IN1(\s1/msel/gnt_p0 [0]), .IN3(\s1/msel/gnt_p2 [0]), .IN2(
        \s1/msel/gnt_p1 [0]), .IN4(\s1/msel/gnt_p3 [0]), .S0(
        \s1/msel/pri_out [1]), .S1(\s1/msel/pri_out [0]), .Q(n23236) );
  MUX41X1 U21272 ( .IN1(\s1/msel/gnt_p0 [1]), .IN3(\s1/msel/gnt_p2 [1]), .IN2(
        \s1/msel/gnt_p1 [1]), .IN4(\s1/msel/gnt_p3 [1]), .S0(
        \s1/msel/pri_out [1]), .S1(\s1/msel/pri_out [0]), .Q(n23140) );
  MUX41X1 U21273 ( .IN1(\s1/msel/gnt_p0 [2]), .IN3(\s1/msel/gnt_p2 [2]), .IN2(
        \s1/msel/gnt_p1 [2]), .IN4(\s1/msel/gnt_p3 [2]), .S0(
        \s1/msel/pri_out [1]), .S1(\s1/msel/pri_out [0]), .Q(n23141) );
  INVX0 U21274 ( .INP(n23141), .ZN(n21135) );
  NOR3X0 U21275 ( .IN1(n23236), .IN2(n23140), .IN3(n21135), .QN(n28992) );
  NAND2X0 U21276 ( .IN1(n29326), .IN2(n28992), .QN(n27805) );
  OA22X1 U21277 ( .IN1(n21144), .IN2(n26584), .IN3(n21138), .IN4(n27805), .Q(
        n19239) );
  INVX0 U21278 ( .INP(s6_ack_i), .ZN(n21126) );
  INVX0 U21279 ( .INP(m4s0_addr[29]), .ZN(n28923) );
  NOR2X0 U21280 ( .IN1(m4s0_addr[28]), .IN2(n28923), .QN(n19246) );
  NAND2X0 U21281 ( .IN1(n19242), .IN2(n19246), .QN(n19643) );
  INVX0 U21282 ( .INP(n19643), .ZN(n29321) );
  MUX41X1 U21283 ( .IN1(\s6/msel/gnt_p0 [2]), .IN3(\s6/msel/gnt_p2 [2]), .IN2(
        \s6/msel/gnt_p1 [2]), .IN4(\s6/msel/gnt_p3 [2]), .S0(
        \s6/msel/pri_out [1]), .S1(\s6/msel/pri_out [0]), .Q(n23137) );
  INVX0 U21284 ( .INP(n23137), .ZN(n21125) );
  MUX41X1 U21285 ( .IN1(\s6/msel/gnt_p0 [0]), .IN3(\s6/msel/gnt_p2 [0]), .IN2(
        \s6/msel/gnt_p1 [0]), .IN4(\s6/msel/gnt_p3 [0]), .S0(
        \s6/msel/pri_out [1]), .S1(\s6/msel/pri_out [0]), .Q(n23230) );
  MUX41X1 U21286 ( .IN1(\s6/msel/gnt_p0 [1]), .IN3(\s6/msel/gnt_p2 [1]), .IN2(
        \s6/msel/gnt_p1 [1]), .IN4(\s6/msel/gnt_p3 [1]), .S0(
        \s6/msel/pri_out [1]), .S1(\s6/msel/pri_out [0]), .Q(n23136) );
  NOR3X0 U21287 ( .IN1(n21125), .IN2(n23230), .IN3(n23136), .QN(n29083) );
  NAND2X0 U21288 ( .IN1(n29321), .IN2(n29083), .QN(n26283) );
  INVX0 U21289 ( .INP(s3_ack_i), .ZN(n21120) );
  NOR2X0 U21290 ( .IN1(n28906), .IN2(n28923), .QN(n19241) );
  NAND2X0 U21291 ( .IN1(n19241), .IN2(n19245), .QN(n19633) );
  INVX0 U21292 ( .INP(n19633), .ZN(n29324) );
  MUX41X1 U21293 ( .IN1(\s3/msel/gnt_p0 [2]), .IN3(\s3/msel/gnt_p2 [2]), .IN2(
        \s3/msel/gnt_p1 [2]), .IN4(\s3/msel/gnt_p3 [2]), .S0(
        \s3/msel/pri_out [1]), .S1(\s3/msel/pri_out [0]), .Q(n23165) );
  INVX0 U21294 ( .INP(n23165), .ZN(n21118) );
  MUX41X1 U21295 ( .IN1(\s3/msel/gnt_p0 [0]), .IN3(\s3/msel/gnt_p2 [0]), .IN2(
        \s3/msel/gnt_p1 [0]), .IN4(\s3/msel/gnt_p3 [0]), .S0(
        \s3/msel/pri_out [1]), .S1(\s3/msel/pri_out [0]), .Q(n23233) );
  MUX41X1 U21296 ( .IN1(\s3/msel/gnt_p0 [1]), .IN3(\s3/msel/gnt_p2 [1]), .IN2(
        \s3/msel/gnt_p1 [1]), .IN4(\s3/msel/gnt_p3 [1]), .S0(
        \s3/msel/pri_out [1]), .S1(\s3/msel/pri_out [0]), .Q(n23164) );
  NOR3X0 U21297 ( .IN1(n21118), .IN2(n23233), .IN3(n23164), .QN(n29022) );
  NAND2X0 U21298 ( .IN1(n29324), .IN2(n29022), .QN(n27195) );
  OA22X1 U21299 ( .IN1(n21126), .IN2(n26283), .IN3(n21120), .IN4(n27195), .Q(
        n19238) );
  INVX0 U21300 ( .INP(s2_ack_i), .ZN(n23214) );
  AND2X1 U21301 ( .IN1(n19245), .IN2(n19246), .Q(n29325) );
  MUX41X1 U21302 ( .IN1(\s2/msel/gnt_p0 [2]), .IN3(\s2/msel/gnt_p1 [2]), .IN2(
        \s2/msel/gnt_p2 [2]), .IN4(\s2/msel/gnt_p3 [2]), .S0(
        \s2/msel/pri_out [0]), .S1(\s2/msel/pri_out [1]), .Q(n23112) );
  INVX0 U21303 ( .INP(n23112), .ZN(n21133) );
  MUX41X1 U21304 ( .IN1(\s2/msel/gnt_p0 [1]), .IN3(\s2/msel/gnt_p1 [1]), .IN2(
        \s2/msel/gnt_p2 [1]), .IN4(\s2/msel/gnt_p3 [1]), .S0(
        \s2/msel/pri_out [0]), .S1(\s2/msel/pri_out [1]), .Q(n23113) );
  MUX41X1 U21305 ( .IN1(\s2/msel/gnt_p0 [0]), .IN3(\s2/msel/gnt_p1 [0]), .IN2(
        \s2/msel/gnt_p2 [0]), .IN4(\s2/msel/gnt_p3 [0]), .S0(
        \s2/msel/pri_out [0]), .S1(\s2/msel/pri_out [1]), .Q(n23114) );
  NOR3X0 U21306 ( .IN1(n21133), .IN2(n23113), .IN3(n23114), .QN(n29012) );
  NAND2X0 U21307 ( .IN1(n29325), .IN2(n29012), .QN(n27504) );
  INVX0 U21308 ( .INP(s12_ack_i), .ZN(n21141) );
  INVX0 U21309 ( .INP(m4s0_addr[31]), .ZN(n28946) );
  NOR2X0 U21310 ( .IN1(n28946), .IN2(n28939), .QN(n19243) );
  NOR2X0 U21311 ( .IN1(m4s0_addr[28]), .IN2(m4s0_addr[29]), .QN(n19244) );
  AND2X1 U21312 ( .IN1(n19243), .IN2(n19244), .Q(n29315) );
  MUX41X1 U21313 ( .IN1(\s12/msel/gnt_p0 [1]), .IN3(\s12/msel/gnt_p1 [1]), 
        .IN2(\s12/msel/gnt_p2 [1]), .IN4(\s12/msel/gnt_p3 [1]), .S0(
        \s12/msel/pri_out [0]), .S1(\s12/msel/pri_out [1]), .Q(n23151) );
  MUX41X1 U21314 ( .IN1(\s12/msel/gnt_p0 [2]), .IN3(\s12/msel/gnt_p1 [2]), 
        .IN2(\s12/msel/gnt_p2 [2]), .IN4(\s12/msel/gnt_p3 [2]), .S0(
        \s12/msel/pri_out [0]), .S1(\s12/msel/pri_out [1]), .Q(n23150) );
  INVX0 U21315 ( .INP(n23150), .ZN(n21139) );
  MUX41X1 U21316 ( .IN1(\s12/msel/gnt_p0 [0]), .IN3(\s12/msel/gnt_p1 [0]), 
        .IN2(\s12/msel/gnt_p2 [0]), .IN4(\s12/msel/gnt_p3 [0]), .S0(
        \s12/msel/pri_out [0]), .S1(\s12/msel/pri_out [1]), .Q(n23224) );
  NOR3X0 U21317 ( .IN1(n23151), .IN2(n21139), .IN3(n23224), .QN(n29182) );
  NAND2X0 U21318 ( .IN1(n29315), .IN2(n29182), .QN(n24452) );
  OA22X1 U21319 ( .IN1(n23214), .IN2(n27504), .IN3(n21141), .IN4(n24452), .Q(
        n19237) );
  INVX0 U21320 ( .INP(s8_ack_i), .ZN(n23246) );
  NOR2X0 U21321 ( .IN1(m4s0_addr[30]), .IN2(n28946), .QN(n19247) );
  AND2X1 U21322 ( .IN1(n19247), .IN2(n19244), .Q(n29319) );
  MUX41X1 U21323 ( .IN1(\s8/msel/gnt_p0 [2]), .IN3(\s8/msel/gnt_p2 [2]), .IN2(
        \s8/msel/gnt_p1 [2]), .IN4(\s8/msel/gnt_p3 [2]), .S0(
        \s8/msel/pri_out [1]), .S1(\s8/msel/pri_out [0]), .Q(n23121) );
  INVX0 U21324 ( .INP(n23121), .ZN(n19665) );
  MUX41X1 U21325 ( .IN1(\s8/msel/gnt_p0 [1]), .IN3(\s8/msel/gnt_p2 [1]), .IN2(
        \s8/msel/gnt_p1 [1]), .IN4(\s8/msel/gnt_p3 [1]), .S0(
        \s8/msel/pri_out [1]), .S1(\s8/msel/pri_out [0]), .Q(n23122) );
  NOR2X0 U21326 ( .IN1(n19665), .IN2(n23122), .QN(n21121) );
  MUX41X1 U21327 ( .IN1(\s8/msel/gnt_p0 [0]), .IN3(\s8/msel/gnt_p2 [0]), .IN2(
        \s8/msel/gnt_p1 [0]), .IN4(\s8/msel/gnt_p3 [0]), .S0(
        \s8/msel/pri_out [1]), .S1(\s8/msel/pri_out [0]), .Q(n23123) );
  INVX0 U21328 ( .INP(n23123), .ZN(n23245) );
  NAND2X0 U21329 ( .IN1(n21121), .IN2(n23245), .QN(n25969) );
  NAND2X0 U21330 ( .IN1(n29319), .IN2(n29110), .QN(n25673) );
  OR2X1 U21331 ( .IN1(n23246), .IN2(n25673), .Q(n19236) );
  NAND4X0 U21332 ( .IN1(n19239), .IN2(n19238), .IN3(n19237), .IN4(n19236), 
        .QN(n19253) );
  INVX0 U21333 ( .INP(s13_ack_i), .ZN(n23213) );
  AND2X1 U21334 ( .IN1(n19243), .IN2(n19240), .Q(n29314) );
  MUX41X1 U21335 ( .IN1(\s13/msel/gnt_p0 [0]), .IN3(\s13/msel/gnt_p1 [0]), 
        .IN2(\s13/msel/gnt_p2 [0]), .IN4(\s13/msel/gnt_p3 [0]), .S0(
        \s13/msel/pri_out [0]), .S1(\s13/msel/pri_out [1]), .Q(n23212) );
  MUX41X1 U21336 ( .IN1(\s13/msel/gnt_p0 [2]), .IN3(\s13/msel/gnt_p1 [2]), 
        .IN2(\s13/msel/gnt_p2 [2]), .IN4(\s13/msel/gnt_p3 [2]), .S0(
        \s13/msel/pri_out [0]), .S1(\s13/msel/pri_out [1]), .Q(n23128) );
  INVX0 U21337 ( .INP(n23128), .ZN(n21127) );
  MUX41X1 U21338 ( .IN1(\s13/msel/gnt_p0 [1]), .IN3(\s13/msel/gnt_p1 [1]), 
        .IN2(\s13/msel/gnt_p2 [1]), .IN4(\s13/msel/gnt_p3 [1]), .S0(
        \s13/msel/pri_out [0]), .S1(\s13/msel/pri_out [1]), .Q(n23129) );
  NOR3X0 U21339 ( .IN1(n23212), .IN2(n21127), .IN3(n23129), .QN(n29209) );
  NAND2X0 U21340 ( .IN1(n29314), .IN2(n29209), .QN(n24154) );
  INVX0 U21341 ( .INP(s11_ack_i), .ZN(n21137) );
  AND2X1 U21342 ( .IN1(n19241), .IN2(n19247), .Q(n29316) );
  MUX41X1 U21343 ( .IN1(\s11/msel/gnt_p0 [1]), .IN3(\s11/msel/gnt_p2 [1]), 
        .IN2(\s11/msel/gnt_p1 [1]), .IN4(\s11/msel/gnt_p3 [1]), .S0(
        \s11/msel/pri_out [1]), .S1(\s11/msel/pri_out [0]), .Q(n23147) );
  MUX41X1 U21344 ( .IN1(\s11/msel/gnt_p0 [0]), .IN3(\s11/msel/gnt_p2 [0]), 
        .IN2(\s11/msel/gnt_p1 [0]), .IN4(\s11/msel/gnt_p3 [0]), .S0(
        \s11/msel/pri_out [1]), .S1(\s11/msel/pri_out [0]), .Q(n23221) );
  MUX41X1 U21345 ( .IN1(\s11/msel/gnt_p0 [2]), .IN3(\s11/msel/gnt_p2 [2]), 
        .IN2(\s11/msel/gnt_p1 [2]), .IN4(\s11/msel/gnt_p3 [2]), .S0(
        \s11/msel/pri_out [1]), .S1(\s11/msel/pri_out [0]), .Q(n23146) );
  INVX0 U21346 ( .INP(n23146), .ZN(n21136) );
  NOR3X0 U21347 ( .IN1(n23147), .IN2(n23221), .IN3(n21136), .QN(n29172) );
  NAND2X0 U21348 ( .IN1(n29316), .IN2(n29172), .QN(n24760) );
  OA22X1 U21349 ( .IN1(n23213), .IN2(n24154), .IN3(n21137), .IN4(n24760), .Q(
        n19251) );
  INVX0 U21350 ( .INP(s9_ack_i), .ZN(n23253) );
  AND2X1 U21351 ( .IN1(n19247), .IN2(n19240), .Q(n29318) );
  MUX41X1 U21352 ( .IN1(\s9/msel/gnt_p0 [2]), .IN3(\s9/msel/gnt_p1 [2]), .IN2(
        \s9/msel/gnt_p2 [2]), .IN4(\s9/msel/gnt_p3 [2]), .S0(
        \s9/msel/pri_out [0]), .S1(\s9/msel/pri_out [1]), .Q(n23115) );
  INVX0 U21353 ( .INP(n23115), .ZN(n21142) );
  MUX41X1 U21354 ( .IN1(\s9/msel/gnt_p0 [1]), .IN3(\s9/msel/gnt_p1 [1]), .IN2(
        \s9/msel/gnt_p2 [1]), .IN4(\s9/msel/gnt_p3 [1]), .S0(
        \s9/msel/pri_out [0]), .S1(\s9/msel/pri_out [1]), .Q(n23116) );
  MUX41X1 U21355 ( .IN1(\s9/msel/gnt_p0 [0]), .IN3(\s9/msel/gnt_p1 [0]), .IN2(
        \s9/msel/gnt_p2 [0]), .IN4(\s9/msel/gnt_p3 [0]), .S0(
        \s9/msel/pri_out [0]), .S1(\s9/msel/pri_out [1]), .Q(n23117) );
  NOR3X0 U21356 ( .IN1(n21142), .IN2(n23116), .IN3(n23117), .QN(n29128) );
  NAND2X0 U21357 ( .IN1(n29318), .IN2(n29128), .QN(n25367) );
  INVX0 U21358 ( .INP(s7_ack_i), .ZN(n23220) );
  NAND2X0 U21359 ( .IN1(n19241), .IN2(n19242), .QN(n19645) );
  INVX0 U21360 ( .INP(n19645), .ZN(n29320) );
  MUX41X1 U21361 ( .IN1(\s7/msel/gnt_p0 [0]), .IN3(\s7/msel/gnt_p1 [0]), .IN2(
        \s7/msel/gnt_p2 [0]), .IN4(\s7/msel/gnt_p3 [0]), .S0(
        \s7/msel/pri_out [0]), .S1(\s7/msel/pri_out [1]), .Q(n23215) );
  MUX41X1 U21362 ( .IN1(\s7/msel/gnt_p0 [2]), .IN3(\s7/msel/gnt_p1 [2]), .IN2(
        \s7/msel/gnt_p2 [2]), .IN4(\s7/msel/gnt_p3 [2]), .S0(
        \s7/msel/pri_out [0]), .S1(\s7/msel/pri_out [1]), .Q(n23144) );
  INVX0 U21363 ( .INP(n23144), .ZN(n21119) );
  MUX41X1 U21364 ( .IN1(\s7/msel/gnt_p0 [1]), .IN3(\s7/msel/gnt_p1 [1]), .IN2(
        \s7/msel/gnt_p2 [1]), .IN4(\s7/msel/gnt_p3 [1]), .S0(
        \s7/msel/pri_out [0]), .S1(\s7/msel/pri_out [1]), .Q(n23143) );
  NOR3X0 U21365 ( .IN1(n23215), .IN2(n21119), .IN3(n23143), .QN(n29101) );
  NAND2X0 U21366 ( .IN1(n29320), .IN2(n29101), .QN(n25975) );
  OA22X1 U21367 ( .IN1(n23253), .IN2(n25367), .IN3(n23220), .IN4(n25975), .Q(
        n19250) );
  INVX0 U21368 ( .INP(s4_ack_i), .ZN(n23247) );
  AND2X1 U21369 ( .IN1(n19244), .IN2(n19242), .Q(n29323) );
  MUX41X1 U21370 ( .IN1(\s4/msel/gnt_p0 [2]), .IN3(\s4/msel/gnt_p2 [2]), .IN2(
        \s4/msel/gnt_p1 [2]), .IN4(\s4/msel/gnt_p3 [2]), .S0(
        \s4/msel/pri_out [1]), .S1(\s4/msel/pri_out [0]), .Q(n23119) );
  INVX0 U21371 ( .INP(n23119), .ZN(n21124) );
  MUX41X1 U21372 ( .IN1(\s4/msel/gnt_p0 [0]), .IN3(\s4/msel/gnt_p2 [0]), .IN2(
        \s4/msel/gnt_p1 [0]), .IN4(\s4/msel/gnt_p3 [0]), .S0(
        \s4/msel/pri_out [1]), .S1(\s4/msel/pri_out [0]), .Q(n23120) );
  MUX41X1 U21373 ( .IN1(\s4/msel/gnt_p0 [1]), .IN3(\s4/msel/gnt_p2 [1]), .IN2(
        \s4/msel/gnt_p1 [1]), .IN4(\s4/msel/gnt_p3 [1]), .S0(
        \s4/msel/pri_out [1]), .S1(\s4/msel/pri_out [0]), .Q(n23118) );
  NOR3X0 U21374 ( .IN1(n21124), .IN2(n23120), .IN3(n23118), .QN(n29048) );
  NAND2X0 U21375 ( .IN1(n29323), .IN2(n29048), .QN(n26891) );
  INVX0 U21376 ( .INP(s14_ack_i), .ZN(n21123) );
  AND2X1 U21377 ( .IN1(n19243), .IN2(n19246), .Q(n29313) );
  MUX41X1 U21378 ( .IN1(\s14/msel/gnt_p0 [0]), .IN3(\s14/msel/gnt_p1 [0]), 
        .IN2(\s14/msel/gnt_p2 [0]), .IN4(\s14/msel/gnt_p3 [0]), .S0(
        \s14/msel/pri_out [0]), .S1(\s14/msel/pri_out [1]), .Q(n23240) );
  MUX41X1 U21379 ( .IN1(\s14/msel/gnt_p0 [1]), .IN3(\s14/msel/gnt_p1 [1]), 
        .IN2(\s14/msel/gnt_p2 [1]), .IN4(\s14/msel/gnt_p3 [1]), .S0(
        \s14/msel/pri_out [0]), .S1(\s14/msel/pri_out [1]), .Q(n23124) );
  MUX41X1 U21380 ( .IN1(\s14/msel/gnt_p0 [2]), .IN3(\s14/msel/gnt_p1 [2]), 
        .IN2(\s14/msel/gnt_p2 [2]), .IN4(\s14/msel/gnt_p3 [2]), .S0(
        \s14/msel/pri_out [0]), .S1(\s14/msel/pri_out [1]), .Q(n23125) );
  INVX0 U21381 ( .INP(n23125), .ZN(n21122) );
  NOR3X0 U21382 ( .IN1(n23240), .IN2(n23124), .IN3(n21122), .QN(n29219) );
  NAND2X0 U21383 ( .IN1(n29313), .IN2(n29219), .QN(n23848) );
  OA22X1 U21384 ( .IN1(n23247), .IN2(n26891), .IN3(n21123), .IN4(n23848), .Q(
        n19249) );
  INVX0 U21385 ( .INP(s0_ack_i), .ZN(n23252) );
  AND2X1 U21386 ( .IN1(n19245), .IN2(n19244), .Q(n29328) );
  MUX41X1 U21387 ( .IN1(\s0/msel/gnt_p0 [0]), .IN3(\s0/msel/gnt_p2 [0]), .IN2(
        \s0/msel/gnt_p1 [0]), .IN4(\s0/msel/gnt_p3 [0]), .S0(
        \s0/msel/pri_out [1]), .S1(\s0/msel/pri_out [0]), .Q(n23251) );
  MUX41X1 U21388 ( .IN1(\s0/msel/gnt_p0 [1]), .IN3(\s0/msel/gnt_p2 [1]), .IN2(
        \s0/msel/gnt_p1 [1]), .IN4(\s0/msel/gnt_p3 [1]), .S0(
        \s0/msel/pri_out [1]), .S1(\s0/msel/pri_out [0]), .Q(n23154) );
  MUX41X1 U21389 ( .IN1(\s0/msel/gnt_p0 [2]), .IN3(\s0/msel/gnt_p2 [2]), .IN2(
        \s0/msel/gnt_p1 [2]), .IN4(\s0/msel/gnt_p3 [2]), .S0(
        \s0/msel/pri_out [1]), .S1(\s0/msel/pri_out [0]), .Q(n23155) );
  INVX0 U21390 ( .INP(n23155), .ZN(n21140) );
  NOR3X0 U21391 ( .IN1(n23251), .IN2(n23154), .IN3(n21140), .QN(n28973) );
  NAND2X0 U21392 ( .IN1(n29328), .IN2(n28973), .QN(n28115) );
  INVX0 U21393 ( .INP(s10_ack_i), .ZN(n23219) );
  AND2X1 U21394 ( .IN1(n19247), .IN2(n19246), .Q(n29317) );
  MUX41X1 U21395 ( .IN1(\s10/msel/gnt_p0 [0]), .IN3(\s10/msel/gnt_p1 [0]), 
        .IN2(\s10/msel/gnt_p2 [0]), .IN4(\s10/msel/gnt_p3 [0]), .S0(
        \s10/msel/pri_out [0]), .S1(\s10/msel/pri_out [1]), .Q(n23217) );
  MUX41X1 U21396 ( .IN1(\s10/msel/gnt_p0 [2]), .IN3(\s10/msel/gnt_p1 [2]), 
        .IN2(\s10/msel/gnt_p2 [2]), .IN4(\s10/msel/gnt_p3 [2]), .S0(
        \s10/msel/pri_out [0]), .S1(\s10/msel/pri_out [1]), .Q(n23159) );
  INVX0 U21397 ( .INP(n23159), .ZN(n21134) );
  MUX41X1 U21398 ( .IN1(\s10/msel/gnt_p0 [1]), .IN3(\s10/msel/gnt_p1 [1]), 
        .IN2(\s10/msel/gnt_p2 [1]), .IN4(\s10/msel/gnt_p3 [1]), .S0(
        \s10/msel/pri_out [0]), .S1(\s10/msel/pri_out [1]), .Q(n23158) );
  NOR3X0 U21399 ( .IN1(n23217), .IN2(n21134), .IN3(n23158), .QN(n29154) );
  NAND2X0 U21400 ( .IN1(n29317), .IN2(n29154), .QN(n25067) );
  OA22X1 U21401 ( .IN1(n23252), .IN2(n28115), .IN3(n23219), .IN4(n25067), .Q(
        n19248) );
  NAND4X0 U21402 ( .IN1(n19251), .IN2(n19250), .IN3(n19249), .IN4(n19248), 
        .QN(n19252) );
  NOR2X0 U21403 ( .IN1(n19253), .IN2(n19252), .QN(n19255) );
  MUX21X1 U21404 ( .IN1(s15_ack_i), .IN2(\rf/rf_ack ), .S(n23501), .Q(n23261)
         );
  NAND2X0 U21405 ( .IN1(n23339), .IN2(n23261), .QN(n19254) );
  NAND2X0 U21406 ( .IN1(n19255), .IN2(n19254), .QN(m4_ack_o) );
  INVX0 U21407 ( .INP(m0s14_data_i[0]), .ZN(n21154) );
  INVX0 U21408 ( .INP(n29313), .ZN(n19617) );
  INVX0 U21409 ( .INP(m0s0_data_i[0]), .ZN(n22204) );
  INVX0 U21410 ( .INP(n29328), .ZN(n19630) );
  OA22X1 U21411 ( .IN1(n21154), .IN2(n19617), .IN3(n22204), .IN4(n19630), .Q(
        n19259) );
  INVX0 U21412 ( .INP(m0s10_data_i[0]), .ZN(n22207) );
  INVX0 U21413 ( .INP(n29317), .ZN(n19642) );
  INVX0 U21414 ( .INP(m0s7_data_i[0]), .ZN(n21162) );
  OA22X1 U21415 ( .IN1(n22207), .IN2(n19642), .IN3(n21162), .IN4(n19645), .Q(
        n19258) );
  INVX0 U21416 ( .INP(m0s8_data_i[0]), .ZN(n21163) );
  INVX0 U21417 ( .INP(n29319), .ZN(n19644) );
  INVX0 U21418 ( .INP(m0s1_data_i[0]), .ZN(n21161) );
  INVX0 U21419 ( .INP(n29326), .ZN(n19646) );
  OA22X1 U21420 ( .IN1(n21163), .IN2(n19644), .IN3(n21161), .IN4(n19646), .Q(
        n19257) );
  NAND2X0 U21421 ( .IN1(m0s5_data_i[0]), .IN2(n29322), .QN(n19256) );
  NAND4X0 U21422 ( .IN1(n19259), .IN2(n19258), .IN3(n19257), .IN4(n19256), 
        .QN(n19265) );
  INVX0 U21423 ( .INP(m0s13_data_i[0]), .ZN(n21823) );
  INVX0 U21424 ( .INP(n29314), .ZN(n19641) );
  INVX0 U21425 ( .INP(m0s4_data_i[0]), .ZN(n22203) );
  INVX0 U21426 ( .INP(n29323), .ZN(n19632) );
  OA22X1 U21427 ( .IN1(n21823), .IN2(n19641), .IN3(n22203), .IN4(n19632), .Q(
        n19263) );
  INVX0 U21428 ( .INP(m0s11_data_i[0]), .ZN(n22208) );
  INVX0 U21429 ( .INP(n29316), .ZN(n19631) );
  INVX0 U21430 ( .INP(m0s3_data_i[0]), .ZN(n22206) );
  OA22X1 U21431 ( .IN1(n22208), .IN2(n19631), .IN3(n22206), .IN4(n19633), .Q(
        n19262) );
  INVX0 U21432 ( .INP(m0s6_data_i[0]), .ZN(n21153) );
  INVX0 U21433 ( .INP(m0s2_data_i[0]), .ZN(n22205) );
  INVX0 U21434 ( .INP(n29325), .ZN(n19634) );
  OA22X1 U21435 ( .IN1(n21153), .IN2(n19643), .IN3(n22205), .IN4(n19634), .Q(
        n19261) );
  INVX0 U21436 ( .INP(m0s12_data_i[0]), .ZN(n20251) );
  INVX0 U21437 ( .INP(n29315), .ZN(n19635) );
  INVX0 U21438 ( .INP(m0s9_data_i[0]), .ZN(n21159) );
  INVX0 U21439 ( .INP(n29318), .ZN(n19640) );
  OA22X1 U21440 ( .IN1(n20251), .IN2(n19635), .IN3(n21159), .IN4(n19640), .Q(
        n19260) );
  NAND4X0 U21441 ( .IN1(n19263), .IN2(n19262), .IN3(n19261), .IN4(n19260), 
        .QN(n19264) );
  NOR2X0 U21442 ( .IN1(n19265), .IN2(n19264), .QN(n19267) );
  INVX0 U21443 ( .INP(n19458), .ZN(n29312) );
  MUX21X1 U21444 ( .IN1(s15_data_i[0]), .IN2(\rf/rf_dout [0]), .S(n23501), .Q(
        n22218) );
  NAND2X0 U21445 ( .IN1(n29312), .IN2(n22218), .QN(n19266) );
  NAND2X0 U21446 ( .IN1(n19267), .IN2(n19266), .QN(m4_data_o[0]) );
  INVX0 U21447 ( .INP(m0s5_data_i[1]), .ZN(n21177) );
  INVX0 U21448 ( .INP(n29322), .ZN(n19647) );
  INVX0 U21449 ( .INP(m0s0_data_i[1]), .ZN(n22223) );
  OA22X1 U21450 ( .IN1(n21177), .IN2(n19647), .IN3(n22223), .IN4(n19630), .Q(
        n19271) );
  INVX0 U21451 ( .INP(m0s12_data_i[1]), .ZN(n21185) );
  INVX0 U21452 ( .INP(m0s10_data_i[1]), .ZN(n21186) );
  OA22X1 U21453 ( .IN1(n21185), .IN2(n19635), .IN3(n21186), .IN4(n19642), .Q(
        n19270) );
  INVX0 U21454 ( .INP(m0s3_data_i[1]), .ZN(n21176) );
  INVX0 U21455 ( .INP(m0s2_data_i[1]), .ZN(n22225) );
  OA22X1 U21456 ( .IN1(n21176), .IN2(n19633), .IN3(n22225), .IN4(n19634), .Q(
        n19269) );
  NAND2X0 U21457 ( .IN1(m0s11_data_i[1]), .IN2(n29316), .QN(n19268) );
  NAND4X0 U21458 ( .IN1(n19271), .IN2(n19270), .IN3(n19269), .IN4(n19268), 
        .QN(n19277) );
  INVX0 U21459 ( .INP(m0s6_data_i[1]), .ZN(n21175) );
  INVX0 U21460 ( .INP(m0s9_data_i[1]), .ZN(n21183) );
  OA22X1 U21461 ( .IN1(n21175), .IN2(n19643), .IN3(n21183), .IN4(n19640), .Q(
        n19275) );
  INVX0 U21462 ( .INP(m0s1_data_i[1]), .ZN(n21182) );
  INVX0 U21463 ( .INP(m0s8_data_i[1]), .ZN(n21174) );
  OA22X1 U21464 ( .IN1(n21182), .IN2(n19646), .IN3(n21174), .IN4(n19644), .Q(
        n19274) );
  INVX0 U21465 ( .INP(m0s7_data_i[1]), .ZN(n22226) );
  INVX0 U21466 ( .INP(m0s13_data_i[1]), .ZN(n21184) );
  OA22X1 U21467 ( .IN1(n22226), .IN2(n19645), .IN3(n21184), .IN4(n19641), .Q(
        n19273) );
  INVX0 U21468 ( .INP(m0s14_data_i[1]), .ZN(n22224) );
  INVX0 U21469 ( .INP(m0s4_data_i[1]), .ZN(n21173) );
  OA22X1 U21470 ( .IN1(n22224), .IN2(n19617), .IN3(n21173), .IN4(n19632), .Q(
        n19272) );
  NAND4X0 U21471 ( .IN1(n19275), .IN2(n19274), .IN3(n19273), .IN4(n19272), 
        .QN(n19276) );
  NOR2X0 U21472 ( .IN1(n19277), .IN2(n19276), .QN(n19279) );
  INVX0 U21473 ( .INP(n23445), .ZN(n23622) );
  MUX21X1 U21474 ( .IN1(s15_data_i[1]), .IN2(\rf/rf_dout [1]), .S(n23622), .Q(
        n22235) );
  NAND2X0 U21475 ( .IN1(n29312), .IN2(n22235), .QN(n19278) );
  NAND2X0 U21476 ( .IN1(n19279), .IN2(n19278), .QN(m4_data_o[1]) );
  INVX0 U21477 ( .INP(m0s5_data_i[2]), .ZN(n21211) );
  INVX0 U21478 ( .INP(m0s1_data_i[2]), .ZN(n21199) );
  OA22X1 U21479 ( .IN1(n21211), .IN2(n19647), .IN3(n21199), .IN4(n19646), .Q(
        n19283) );
  INVX0 U21480 ( .INP(m0s9_data_i[2]), .ZN(n21210) );
  INVX0 U21481 ( .INP(m0s11_data_i[2]), .ZN(n20702) );
  OA22X1 U21482 ( .IN1(n21210), .IN2(n19640), .IN3(n20702), .IN4(n19631), .Q(
        n19282) );
  INVX0 U21483 ( .INP(m0s4_data_i[2]), .ZN(n21197) );
  INVX0 U21484 ( .INP(m0s0_data_i[2]), .ZN(n21205) );
  OA22X1 U21485 ( .IN1(n21197), .IN2(n19632), .IN3(n21205), .IN4(n19630), .Q(
        n19281) );
  NAND2X0 U21486 ( .IN1(m0s3_data_i[2]), .IN2(n29324), .QN(n19280) );
  NAND4X0 U21487 ( .IN1(n19283), .IN2(n19282), .IN3(n19281), .IN4(n19280), 
        .QN(n19289) );
  INVX0 U21488 ( .INP(m0s12_data_i[2]), .ZN(n21198) );
  INVX0 U21489 ( .INP(m0s10_data_i[2]), .ZN(n21206) );
  OA22X1 U21490 ( .IN1(n21198), .IN2(n19635), .IN3(n21206), .IN4(n19642), .Q(
        n19287) );
  INVX0 U21491 ( .INP(m0s14_data_i[2]), .ZN(n21195) );
  INVX0 U21492 ( .INP(m0s2_data_i[2]), .ZN(n21207) );
  OA22X1 U21493 ( .IN1(n21195), .IN2(n19617), .IN3(n21207), .IN4(n19634), .Q(
        n19286) );
  INVX0 U21494 ( .INP(m0s13_data_i[2]), .ZN(n21212) );
  INVX0 U21495 ( .INP(m0s6_data_i[2]), .ZN(n21208) );
  OA22X1 U21496 ( .IN1(n21212), .IN2(n19641), .IN3(n21208), .IN4(n19643), .Q(
        n19285) );
  INVX0 U21497 ( .INP(m0s7_data_i[2]), .ZN(n21209) );
  INVX0 U21498 ( .INP(m0s8_data_i[2]), .ZN(n21196) );
  OA22X1 U21499 ( .IN1(n21209), .IN2(n19645), .IN3(n21196), .IN4(n19644), .Q(
        n19284) );
  NAND4X0 U21500 ( .IN1(n19287), .IN2(n19286), .IN3(n19285), .IN4(n19284), 
        .QN(n19288) );
  NOR2X0 U21501 ( .IN1(n19289), .IN2(n19288), .QN(n19291) );
  MUX21X1 U21502 ( .IN1(s15_data_i[2]), .IN2(\rf/rf_dout [2]), .S(n23501), .Q(
        n22247) );
  NAND2X0 U21503 ( .IN1(n29312), .IN2(n22247), .QN(n19290) );
  NAND2X0 U21504 ( .IN1(n19291), .IN2(n19290), .QN(m4_data_o[2]) );
  INVX0 U21505 ( .INP(m0s3_data_i[3]), .ZN(n21221) );
  INVX0 U21506 ( .INP(m0s13_data_i[3]), .ZN(n22636) );
  OA22X1 U21507 ( .IN1(n21221), .IN2(n19633), .IN3(n22636), .IN4(n19641), .Q(
        n19295) );
  INVX0 U21508 ( .INP(m0s11_data_i[3]), .ZN(n21234) );
  INVX0 U21509 ( .INP(m0s6_data_i[3]), .ZN(n21224) );
  OA22X1 U21510 ( .IN1(n21234), .IN2(n19631), .IN3(n21224), .IN4(n19643), .Q(
        n19294) );
  INVX0 U21511 ( .INP(m0s12_data_i[3]), .ZN(n22635) );
  INVX0 U21512 ( .INP(m0s9_data_i[3]), .ZN(n21223) );
  OA22X1 U21513 ( .IN1(n22635), .IN2(n19635), .IN3(n21223), .IN4(n19640), .Q(
        n19293) );
  NAND2X0 U21514 ( .IN1(m0s5_data_i[3]), .IN2(n29322), .QN(n19292) );
  NAND4X0 U21515 ( .IN1(n19295), .IN2(n19294), .IN3(n19293), .IN4(n19292), 
        .QN(n19301) );
  INVX0 U21516 ( .INP(m0s0_data_i[3]), .ZN(n21235) );
  INVX0 U21517 ( .INP(m0s14_data_i[3]), .ZN(n21231) );
  OA22X1 U21518 ( .IN1(n21235), .IN2(n19630), .IN3(n21231), .IN4(n19617), .Q(
        n19299) );
  INVX0 U21519 ( .INP(m0s4_data_i[3]), .ZN(n22634) );
  INVX0 U21520 ( .INP(m0s10_data_i[3]), .ZN(n21232) );
  OA22X1 U21521 ( .IN1(n22634), .IN2(n19632), .IN3(n21232), .IN4(n19642), .Q(
        n19298) );
  INVX0 U21522 ( .INP(m0s2_data_i[3]), .ZN(n21225) );
  INVX0 U21523 ( .INP(m0s8_data_i[3]), .ZN(n21233) );
  OA22X1 U21524 ( .IN1(n21225), .IN2(n19634), .IN3(n21233), .IN4(n19644), .Q(
        n19297) );
  INVX0 U21525 ( .INP(m0s7_data_i[3]), .ZN(n21222) );
  INVX0 U21526 ( .INP(m0s1_data_i[3]), .ZN(n21226) );
  OA22X1 U21527 ( .IN1(n21222), .IN2(n19645), .IN3(n21226), .IN4(n19646), .Q(
        n19296) );
  NAND4X0 U21528 ( .IN1(n19299), .IN2(n19298), .IN3(n19297), .IN4(n19296), 
        .QN(n19300) );
  NOR2X0 U21529 ( .IN1(n19301), .IN2(n19300), .QN(n19303) );
  MUX21X1 U21530 ( .IN1(s15_data_i[3]), .IN2(\rf/rf_dout [3]), .S(n23622), .Q(
        n22646) );
  NAND2X0 U21531 ( .IN1(n29312), .IN2(n22646), .QN(n19302) );
  NAND2X0 U21532 ( .IN1(n19303), .IN2(n19302), .QN(m4_data_o[3]) );
  INVX0 U21533 ( .INP(m0s7_data_i[4]), .ZN(n21257) );
  INVX0 U21534 ( .INP(m0s11_data_i[4]), .ZN(n21255) );
  OA22X1 U21535 ( .IN1(n21257), .IN2(n19645), .IN3(n21255), .IN4(n19631), .Q(
        n19307) );
  INVX0 U21536 ( .INP(m0s3_data_i[4]), .ZN(n20727) );
  INVX0 U21537 ( .INP(m0s1_data_i[4]), .ZN(n21246) );
  OA22X1 U21538 ( .IN1(n20727), .IN2(n19633), .IN3(n21246), .IN4(n19646), .Q(
        n19306) );
  INVX0 U21539 ( .INP(m0s6_data_i[4]), .ZN(n21248) );
  INVX0 U21540 ( .INP(m0s4_data_i[4]), .ZN(n22651) );
  OA22X1 U21541 ( .IN1(n21248), .IN2(n19643), .IN3(n22651), .IN4(n19632), .Q(
        n19305) );
  NAND2X0 U21542 ( .IN1(m0s8_data_i[4]), .IN2(n29319), .QN(n19304) );
  NAND4X0 U21543 ( .IN1(n19307), .IN2(n19306), .IN3(n19305), .IN4(n19304), 
        .QN(n19313) );
  INVX0 U21544 ( .INP(m0s12_data_i[4]), .ZN(n22654) );
  INVX0 U21545 ( .INP(m0s10_data_i[4]), .ZN(n21245) );
  OA22X1 U21546 ( .IN1(n22654), .IN2(n19635), .IN3(n21245), .IN4(n19642), .Q(
        n19311) );
  INVX0 U21547 ( .INP(m0s2_data_i[4]), .ZN(n22652) );
  INVX0 U21548 ( .INP(m0s13_data_i[4]), .ZN(n22653) );
  OA22X1 U21549 ( .IN1(n22652), .IN2(n19634), .IN3(n22653), .IN4(n19641), .Q(
        n19310) );
  INVX0 U21550 ( .INP(m0s5_data_i[4]), .ZN(n21253) );
  INVX0 U21551 ( .INP(m0s0_data_i[4]), .ZN(n21254) );
  OA22X1 U21552 ( .IN1(n21253), .IN2(n19647), .IN3(n21254), .IN4(n19630), .Q(
        n19309) );
  INVX0 U21553 ( .INP(m0s9_data_i[4]), .ZN(n21247) );
  INVX0 U21554 ( .INP(m0s14_data_i[4]), .ZN(n21244) );
  OA22X1 U21555 ( .IN1(n21247), .IN2(n19640), .IN3(n21244), .IN4(n19617), .Q(
        n19308) );
  NAND4X0 U21556 ( .IN1(n19311), .IN2(n19310), .IN3(n19309), .IN4(n19308), 
        .QN(n19312) );
  NOR2X0 U21557 ( .IN1(n19313), .IN2(n19312), .QN(n19315) );
  MUX21X1 U21558 ( .IN1(s15_data_i[4]), .IN2(\rf/rf_dout [4]), .S(n23622), .Q(
        n22663) );
  NAND2X0 U21559 ( .IN1(n29312), .IN2(n22663), .QN(n19314) );
  NAND2X0 U21560 ( .IN1(n19315), .IN2(n19314), .QN(m4_data_o[4]) );
  INVX0 U21561 ( .INP(m0s3_data_i[5]), .ZN(n22668) );
  INVX0 U21562 ( .INP(m0s11_data_i[5]), .ZN(n21268) );
  OA22X1 U21563 ( .IN1(n22668), .IN2(n19633), .IN3(n21268), .IN4(n19631), .Q(
        n19319) );
  INVX0 U21564 ( .INP(m0s0_data_i[5]), .ZN(n21277) );
  INVX0 U21565 ( .INP(m0s7_data_i[5]), .ZN(n22670) );
  OA22X1 U21566 ( .IN1(n21277), .IN2(n19630), .IN3(n22670), .IN4(n19645), .Q(
        n19318) );
  INVX0 U21567 ( .INP(m0s4_data_i[5]), .ZN(n21269) );
  INVX0 U21568 ( .INP(m0s13_data_i[5]), .ZN(n22671) );
  OA22X1 U21569 ( .IN1(n21269), .IN2(n19632), .IN3(n22671), .IN4(n19641), .Q(
        n19317) );
  NAND2X0 U21570 ( .IN1(m0s10_data_i[5]), .IN2(n29317), .QN(n19316) );
  NAND4X0 U21571 ( .IN1(n19319), .IN2(n19318), .IN3(n19317), .IN4(n19316), 
        .QN(n19325) );
  INVX0 U21572 ( .INP(m0s2_data_i[5]), .ZN(n22669) );
  INVX0 U21573 ( .INP(m0s1_data_i[5]), .ZN(n21274) );
  OA22X1 U21574 ( .IN1(n22669), .IN2(n19634), .IN3(n21274), .IN4(n19646), .Q(
        n19323) );
  INVX0 U21575 ( .INP(m0s12_data_i[5]), .ZN(n21266) );
  INVX0 U21576 ( .INP(m0s9_data_i[5]), .ZN(n21267) );
  OA22X1 U21577 ( .IN1(n21266), .IN2(n19635), .IN3(n21267), .IN4(n19640), .Q(
        n19322) );
  INVX0 U21578 ( .INP(m0s6_data_i[5]), .ZN(n21279) );
  INVX0 U21579 ( .INP(m0s14_data_i[5]), .ZN(n21275) );
  OA22X1 U21580 ( .IN1(n21279), .IN2(n19643), .IN3(n21275), .IN4(n19617), .Q(
        n19321) );
  INVX0 U21581 ( .INP(m0s5_data_i[5]), .ZN(n20736) );
  INVX0 U21582 ( .INP(m0s8_data_i[5]), .ZN(n21276) );
  OA22X1 U21583 ( .IN1(n20736), .IN2(n19647), .IN3(n21276), .IN4(n19644), .Q(
        n19320) );
  NAND4X0 U21584 ( .IN1(n19323), .IN2(n19322), .IN3(n19321), .IN4(n19320), 
        .QN(n19324) );
  NOR2X0 U21585 ( .IN1(n19325), .IN2(n19324), .QN(n19327) );
  MUX21X1 U21586 ( .IN1(s15_data_i[5]), .IN2(\rf/rf_dout [5]), .S(n23622), .Q(
        n22680) );
  NAND2X0 U21587 ( .IN1(n29312), .IN2(n22680), .QN(n19326) );
  NAND2X0 U21588 ( .IN1(n19327), .IN2(n19326), .QN(m4_data_o[5]) );
  INVX0 U21589 ( .INP(m0s6_data_i[6]), .ZN(n21298) );
  INVX0 U21590 ( .INP(m0s3_data_i[6]), .ZN(n22685) );
  OA22X1 U21591 ( .IN1(n21298), .IN2(n19643), .IN3(n22685), .IN4(n19633), .Q(
        n19331) );
  INVX0 U21592 ( .INP(m0s10_data_i[6]), .ZN(n22686) );
  INVX0 U21593 ( .INP(m0s4_data_i[6]), .ZN(n21290) );
  OA22X1 U21594 ( .IN1(n22686), .IN2(n19642), .IN3(n21290), .IN4(n19632), .Q(
        n19330) );
  INVX0 U21595 ( .INP(m0s2_data_i[6]), .ZN(n21297) );
  INVX0 U21596 ( .INP(m0s11_data_i[6]), .ZN(n20753) );
  OA22X1 U21597 ( .IN1(n21297), .IN2(n19634), .IN3(n20753), .IN4(n19631), .Q(
        n19329) );
  NAND2X0 U21598 ( .IN1(m0s7_data_i[6]), .IN2(n29320), .QN(n19328) );
  NAND4X0 U21599 ( .IN1(n19331), .IN2(n19330), .IN3(n19329), .IN4(n19328), 
        .QN(n19337) );
  INVX0 U21600 ( .INP(m0s8_data_i[6]), .ZN(n22688) );
  INVX0 U21601 ( .INP(m0s14_data_i[6]), .ZN(n21288) );
  OA22X1 U21602 ( .IN1(n22688), .IN2(n19644), .IN3(n21288), .IN4(n19617), .Q(
        n19335) );
  INVX0 U21603 ( .INP(m0s13_data_i[6]), .ZN(n22687) );
  INVX0 U21604 ( .INP(m0s0_data_i[6]), .ZN(n21299) );
  OA22X1 U21605 ( .IN1(n22687), .IN2(n19641), .IN3(n21299), .IN4(n19630), .Q(
        n19334) );
  INVX0 U21606 ( .INP(m0s5_data_i[6]), .ZN(n21292) );
  INVX0 U21607 ( .INP(m0s1_data_i[6]), .ZN(n21301) );
  OA22X1 U21608 ( .IN1(n21292), .IN2(n19647), .IN3(n21301), .IN4(n19646), .Q(
        n19333) );
  INVX0 U21609 ( .INP(m0s12_data_i[6]), .ZN(n21291) );
  INVX0 U21610 ( .INP(m0s9_data_i[6]), .ZN(n21300) );
  OA22X1 U21611 ( .IN1(n21291), .IN2(n19635), .IN3(n21300), .IN4(n19640), .Q(
        n19332) );
  NAND4X0 U21612 ( .IN1(n19335), .IN2(n19334), .IN3(n19333), .IN4(n19332), 
        .QN(n19336) );
  NOR2X0 U21613 ( .IN1(n19337), .IN2(n19336), .QN(n19339) );
  MUX21X1 U21614 ( .IN1(s15_data_i[6]), .IN2(\rf/rf_dout [6]), .S(n23622), .Q(
        n22697) );
  NAND2X0 U21615 ( .IN1(n29312), .IN2(n22697), .QN(n19338) );
  NAND2X0 U21616 ( .IN1(n19339), .IN2(n19338), .QN(m4_data_o[6]) );
  INVX0 U21617 ( .INP(m0s12_data_i[7]), .ZN(n22704) );
  INVX0 U21618 ( .INP(m0s7_data_i[7]), .ZN(n20766) );
  OA22X1 U21619 ( .IN1(n22704), .IN2(n19635), .IN3(n20766), .IN4(n19645), .Q(
        n19343) );
  INVX0 U21620 ( .INP(m0s6_data_i[7]), .ZN(n21321) );
  INVX0 U21621 ( .INP(m0s13_data_i[7]), .ZN(n21313) );
  OA22X1 U21622 ( .IN1(n21321), .IN2(n19643), .IN3(n21313), .IN4(n19641), .Q(
        n19342) );
  INVX0 U21623 ( .INP(m0s9_data_i[7]), .ZN(n21322) );
  INVX0 U21624 ( .INP(m0s11_data_i[7]), .ZN(n21310) );
  OA22X1 U21625 ( .IN1(n21322), .IN2(n19640), .IN3(n21310), .IN4(n19631), .Q(
        n19341) );
  NAND2X0 U21626 ( .IN1(m0s0_data_i[7]), .IN2(n29328), .QN(n19340) );
  NAND4X0 U21627 ( .IN1(n19343), .IN2(n19342), .IN3(n19341), .IN4(n19340), 
        .QN(n19349) );
  INVX0 U21628 ( .INP(m0s8_data_i[7]), .ZN(n21319) );
  INVX0 U21629 ( .INP(m0s3_data_i[7]), .ZN(n21320) );
  OA22X1 U21630 ( .IN1(n21319), .IN2(n19644), .IN3(n21320), .IN4(n19633), .Q(
        n19347) );
  INVX0 U21631 ( .INP(m0s5_data_i[7]), .ZN(n21312) );
  INVX0 U21632 ( .INP(m0s10_data_i[7]), .ZN(n21314) );
  OA22X1 U21633 ( .IN1(n21312), .IN2(n19647), .IN3(n21314), .IN4(n19642), .Q(
        n19346) );
  INVX0 U21634 ( .INP(m0s4_data_i[7]), .ZN(n22705) );
  INVX0 U21635 ( .INP(m0s2_data_i[7]), .ZN(n22702) );
  OA22X1 U21636 ( .IN1(n22705), .IN2(n19632), .IN3(n22702), .IN4(n19634), .Q(
        n19345) );
  INVX0 U21637 ( .INP(m0s1_data_i[7]), .ZN(n21311) );
  INVX0 U21638 ( .INP(m0s14_data_i[7]), .ZN(n21323) );
  OA22X1 U21639 ( .IN1(n21311), .IN2(n19646), .IN3(n21323), .IN4(n19617), .Q(
        n19344) );
  NAND4X0 U21640 ( .IN1(n19347), .IN2(n19346), .IN3(n19345), .IN4(n19344), 
        .QN(n19348) );
  NOR2X0 U21641 ( .IN1(n19349), .IN2(n19348), .QN(n19351) );
  MUX21X1 U21642 ( .IN1(s15_data_i[7]), .IN2(\rf/rf_dout [7]), .S(n23622), .Q(
        n22714) );
  NAND2X0 U21643 ( .IN1(n29312), .IN2(n22714), .QN(n19350) );
  NAND2X0 U21644 ( .IN1(n19351), .IN2(n19350), .QN(m4_data_o[7]) );
  INVX0 U21645 ( .INP(m0s6_data_i[8]), .ZN(n21345) );
  INVX0 U21646 ( .INP(m0s2_data_i[8]), .ZN(n21336) );
  OA22X1 U21647 ( .IN1(n21345), .IN2(n19643), .IN3(n21336), .IN4(n19634), .Q(
        n19355) );
  INVX0 U21648 ( .INP(m0s7_data_i[8]), .ZN(n22720) );
  INVX0 U21649 ( .INP(m0s14_data_i[8]), .ZN(n21343) );
  OA22X1 U21650 ( .IN1(n22720), .IN2(n19645), .IN3(n21343), .IN4(n19617), .Q(
        n19354) );
  INVX0 U21651 ( .INP(m0s5_data_i[8]), .ZN(n21342) );
  INVX0 U21652 ( .INP(m0s1_data_i[8]), .ZN(n22722) );
  OA22X1 U21653 ( .IN1(n21342), .IN2(n19647), .IN3(n22722), .IN4(n19646), .Q(
        n19353) );
  NAND2X0 U21654 ( .IN1(m0s11_data_i[8]), .IN2(n29316), .QN(n19352) );
  NAND4X0 U21655 ( .IN1(n19355), .IN2(n19354), .IN3(n19353), .IN4(n19352), 
        .QN(n19361) );
  INVX0 U21656 ( .INP(m0s4_data_i[8]), .ZN(n21335) );
  INVX0 U21657 ( .INP(m0s0_data_i[8]), .ZN(n22721) );
  OA22X1 U21658 ( .IN1(n21335), .IN2(n19632), .IN3(n22721), .IN4(n19630), .Q(
        n19359) );
  INVX0 U21659 ( .INP(m0s10_data_i[8]), .ZN(n21337) );
  INVX0 U21660 ( .INP(m0s9_data_i[8]), .ZN(n21332) );
  OA22X1 U21661 ( .IN1(n21337), .IN2(n19642), .IN3(n21332), .IN4(n19640), .Q(
        n19358) );
  INVX0 U21662 ( .INP(m0s13_data_i[8]), .ZN(n21346) );
  INVX0 U21663 ( .INP(m0s3_data_i[8]), .ZN(n21334) );
  OA22X1 U21664 ( .IN1(n21346), .IN2(n19641), .IN3(n21334), .IN4(n19633), .Q(
        n19357) );
  INVX0 U21665 ( .INP(m0s12_data_i[8]), .ZN(n21344) );
  INVX0 U21666 ( .INP(m0s8_data_i[8]), .ZN(n22719) );
  OA22X1 U21667 ( .IN1(n21344), .IN2(n19635), .IN3(n22719), .IN4(n19644), .Q(
        n19356) );
  NAND4X0 U21668 ( .IN1(n19359), .IN2(n19358), .IN3(n19357), .IN4(n19356), 
        .QN(n19360) );
  NOR2X0 U21669 ( .IN1(n19361), .IN2(n19360), .QN(n19363) );
  MUX21X1 U21670 ( .IN1(s15_data_i[8]), .IN2(\rf/rf_dout [8]), .S(n23622), .Q(
        n22731) );
  NAND2X0 U21671 ( .IN1(n29312), .IN2(n22731), .QN(n19362) );
  NAND2X0 U21672 ( .IN1(n19363), .IN2(n19362), .QN(m4_data_o[8]) );
  INVX0 U21673 ( .INP(m0s4_data_i[9]), .ZN(n22980) );
  INVX0 U21674 ( .INP(m0s14_data_i[9]), .ZN(n21365) );
  OA22X1 U21675 ( .IN1(n22980), .IN2(n19632), .IN3(n21365), .IN4(n19617), .Q(
        n19367) );
  INVX0 U21676 ( .INP(m0s3_data_i[9]), .ZN(n22981) );
  INVX0 U21677 ( .INP(m0s0_data_i[9]), .ZN(n21362) );
  OA22X1 U21678 ( .IN1(n22981), .IN2(n19633), .IN3(n21362), .IN4(n19630), .Q(
        n19366) );
  INVX0 U21679 ( .INP(m0s2_data_i[9]), .ZN(n21357) );
  INVX0 U21680 ( .INP(m0s8_data_i[9]), .ZN(n22978) );
  OA22X1 U21681 ( .IN1(n21357), .IN2(n19634), .IN3(n22978), .IN4(n19644), .Q(
        n19365) );
  NAND2X0 U21682 ( .IN1(m0s13_data_i[9]), .IN2(n29314), .QN(n19364) );
  NAND4X0 U21683 ( .IN1(n19367), .IN2(n19366), .IN3(n19365), .IN4(n19364), 
        .QN(n19373) );
  INVX0 U21684 ( .INP(m0s6_data_i[9]), .ZN(n21356) );
  INVX0 U21685 ( .INP(m0s7_data_i[9]), .ZN(n22736) );
  OA22X1 U21686 ( .IN1(n21356), .IN2(n19643), .IN3(n22736), .IN4(n19645), .Q(
        n19371) );
  INVX0 U21687 ( .INP(m0s10_data_i[9]), .ZN(n21364) );
  INVX0 U21688 ( .INP(m0s1_data_i[9]), .ZN(n20787) );
  OA22X1 U21689 ( .IN1(n21364), .IN2(n19642), .IN3(n20787), .IN4(n19646), .Q(
        n19370) );
  INVX0 U21690 ( .INP(m0s12_data_i[9]), .ZN(n22979) );
  INVX0 U21691 ( .INP(m0s11_data_i[9]), .ZN(n21355) );
  OA22X1 U21692 ( .IN1(n22979), .IN2(n19635), .IN3(n21355), .IN4(n19631), .Q(
        n19369) );
  INVX0 U21693 ( .INP(m0s9_data_i[9]), .ZN(n22984) );
  INVX0 U21694 ( .INP(m0s5_data_i[9]), .ZN(n22983) );
  OA22X1 U21695 ( .IN1(n22984), .IN2(n19640), .IN3(n22983), .IN4(n19647), .Q(
        n19368) );
  NAND4X0 U21696 ( .IN1(n19371), .IN2(n19370), .IN3(n19369), .IN4(n19368), 
        .QN(n19372) );
  NOR2X0 U21697 ( .IN1(n19373), .IN2(n19372), .QN(n19375) );
  MUX21X1 U21698 ( .IN1(s15_data_i[9]), .IN2(\rf/rf_dout [9]), .S(n23622), .Q(
        n22993) );
  NAND2X0 U21699 ( .IN1(n29312), .IN2(n22993), .QN(n19374) );
  NAND2X0 U21700 ( .IN1(n19375), .IN2(n19374), .QN(m4_data_o[9]) );
  INVX0 U21701 ( .INP(m0s7_data_i[10]), .ZN(n22750) );
  INVX0 U21702 ( .INP(m0s0_data_i[10]), .ZN(n21375) );
  OA22X1 U21703 ( .IN1(n22750), .IN2(n19645), .IN3(n21375), .IN4(n19630), .Q(
        n19379) );
  INVX0 U21704 ( .INP(m0s13_data_i[10]), .ZN(n21383) );
  INVX0 U21705 ( .INP(m0s1_data_i[10]), .ZN(n21384) );
  OA22X1 U21706 ( .IN1(n21383), .IN2(n19641), .IN3(n21384), .IN4(n19646), .Q(
        n19378) );
  INVX0 U21707 ( .INP(m0s3_data_i[10]), .ZN(n22752) );
  INVX0 U21708 ( .INP(m0s14_data_i[10]), .ZN(n22329) );
  OA22X1 U21709 ( .IN1(n22752), .IN2(n19633), .IN3(n22329), .IN4(n19617), .Q(
        n19377) );
  NAND2X0 U21710 ( .IN1(m0s2_data_i[10]), .IN2(n29325), .QN(n19376) );
  NAND4X0 U21711 ( .IN1(n19379), .IN2(n19378), .IN3(n19377), .IN4(n19376), 
        .QN(n19385) );
  INVX0 U21712 ( .INP(m0s4_data_i[10]), .ZN(n22753) );
  INVX0 U21713 ( .INP(m0s5_data_i[10]), .ZN(n21376) );
  OA22X1 U21714 ( .IN1(n22753), .IN2(n19632), .IN3(n21376), .IN4(n19647), .Q(
        n19383) );
  INVX0 U21715 ( .INP(m0s11_data_i[10]), .ZN(n21382) );
  INVX0 U21716 ( .INP(m0s6_data_i[10]), .ZN(n21374) );
  OA22X1 U21717 ( .IN1(n21382), .IN2(n19631), .IN3(n21374), .IN4(n19643), .Q(
        n19382) );
  INVX0 U21718 ( .INP(m0s8_data_i[10]), .ZN(n21377) );
  INVX0 U21719 ( .INP(m0s10_data_i[10]), .ZN(n22751) );
  OA22X1 U21720 ( .IN1(n21377), .IN2(n19644), .IN3(n22751), .IN4(n19642), .Q(
        n19381) );
  INVX0 U21721 ( .INP(m0s9_data_i[10]), .ZN(n21385) );
  INVX0 U21722 ( .INP(m0s12_data_i[10]), .ZN(n22754) );
  OA22X1 U21723 ( .IN1(n21385), .IN2(n19640), .IN3(n22754), .IN4(n19635), .Q(
        n19380) );
  NAND4X0 U21724 ( .IN1(n19383), .IN2(n19382), .IN3(n19381), .IN4(n19380), 
        .QN(n19384) );
  NOR2X0 U21725 ( .IN1(n19385), .IN2(n19384), .QN(n19387) );
  MUX21X1 U21726 ( .IN1(s15_data_i[10]), .IN2(\rf/rf_dout [10]), .S(n23622), 
        .Q(n22763) );
  NAND2X0 U21727 ( .IN1(n29312), .IN2(n22763), .QN(n19386) );
  NAND2X0 U21728 ( .IN1(n19387), .IN2(n19386), .QN(m4_data_o[10]) );
  INVX0 U21729 ( .INP(m0s12_data_i[11]), .ZN(n21397) );
  INVX0 U21730 ( .INP(m0s3_data_i[11]), .ZN(n23002) );
  OA22X1 U21731 ( .IN1(n21397), .IN2(n19635), .IN3(n23002), .IN4(n19633), .Q(
        n19391) );
  INVX0 U21732 ( .INP(m0s0_data_i[11]), .ZN(n21398) );
  INVX0 U21733 ( .INP(m0s8_data_i[11]), .ZN(n23000) );
  OA22X1 U21734 ( .IN1(n21398), .IN2(n19630), .IN3(n23000), .IN4(n19644), .Q(
        n19390) );
  INVX0 U21735 ( .INP(m0s14_data_i[11]), .ZN(n22999) );
  INVX0 U21736 ( .INP(m0s9_data_i[11]), .ZN(n21396) );
  OA22X1 U21737 ( .IN1(n22999), .IN2(n19617), .IN3(n21396), .IN4(n19640), .Q(
        n19389) );
  NAND2X0 U21738 ( .IN1(m0s5_data_i[11]), .IN2(n29322), .QN(n19388) );
  NAND4X0 U21739 ( .IN1(n19391), .IN2(n19390), .IN3(n19389), .IN4(n19388), 
        .QN(n19397) );
  INVX0 U21740 ( .INP(m0s6_data_i[11]), .ZN(n23004) );
  INVX0 U21741 ( .INP(m0s11_data_i[11]), .ZN(n23001) );
  OA22X1 U21742 ( .IN1(n23004), .IN2(n19643), .IN3(n23001), .IN4(n19631), .Q(
        n19395) );
  INVX0 U21743 ( .INP(m0s2_data_i[11]), .ZN(n21399) );
  INVX0 U21744 ( .INP(m0s4_data_i[11]), .ZN(n22998) );
  OA22X1 U21745 ( .IN1(n21399), .IN2(n19634), .IN3(n22998), .IN4(n19632), .Q(
        n19394) );
  INVX0 U21746 ( .INP(m0s7_data_i[11]), .ZN(n21405) );
  INVX0 U21747 ( .INP(m0s10_data_i[11]), .ZN(n21395) );
  OA22X1 U21748 ( .IN1(n21405), .IN2(n19645), .IN3(n21395), .IN4(n19642), .Q(
        n19393) );
  INVX0 U21749 ( .INP(m0s13_data_i[11]), .ZN(n21406) );
  INVX0 U21750 ( .INP(m0s1_data_i[11]), .ZN(n21404) );
  OA22X1 U21751 ( .IN1(n21406), .IN2(n19641), .IN3(n21404), .IN4(n19646), .Q(
        n19392) );
  NAND4X0 U21752 ( .IN1(n19395), .IN2(n19394), .IN3(n19393), .IN4(n19392), 
        .QN(n19396) );
  NOR2X0 U21753 ( .IN1(n19397), .IN2(n19396), .QN(n19399) );
  MUX21X1 U21754 ( .IN1(s15_data_i[11]), .IN2(\rf/rf_dout [11]), .S(n23622), 
        .Q(n23013) );
  NAND2X0 U21755 ( .IN1(n29312), .IN2(n23013), .QN(n19398) );
  NAND2X0 U21756 ( .IN1(n19399), .IN2(n19398), .QN(m4_data_o[11]) );
  INVX0 U21757 ( .INP(m0s14_data_i[12]), .ZN(n23024) );
  INVX0 U21758 ( .INP(m0s2_data_i[12]), .ZN(n23026) );
  OA22X1 U21759 ( .IN1(n23024), .IN2(n19617), .IN3(n23026), .IN4(n19634), .Q(
        n19403) );
  INVX0 U21760 ( .INP(m0s8_data_i[12]), .ZN(n21416) );
  INVX0 U21761 ( .INP(m0s1_data_i[12]), .ZN(n23020) );
  OA22X1 U21762 ( .IN1(n21416), .IN2(n19644), .IN3(n23020), .IN4(n19646), .Q(
        n19402) );
  INVX0 U21763 ( .INP(m0s12_data_i[12]), .ZN(n23025) );
  INVX0 U21764 ( .INP(m0s13_data_i[12]), .ZN(n22780) );
  OA22X1 U21765 ( .IN1(n23025), .IN2(n19635), .IN3(n22780), .IN4(n19641), .Q(
        n19401) );
  NAND2X0 U21766 ( .IN1(m0s5_data_i[12]), .IN2(n29322), .QN(n19400) );
  NAND4X0 U21767 ( .IN1(n19403), .IN2(n19402), .IN3(n19401), .IN4(n19400), 
        .QN(n19409) );
  INVX0 U21768 ( .INP(m0s7_data_i[12]), .ZN(n21422) );
  INVX0 U21769 ( .INP(m0s11_data_i[12]), .ZN(n23018) );
  OA22X1 U21770 ( .IN1(n21422), .IN2(n19645), .IN3(n23018), .IN4(n19631), .Q(
        n19407) );
  INVX0 U21771 ( .INP(m0s9_data_i[12]), .ZN(n23022) );
  INVX0 U21772 ( .INP(m0s6_data_i[12]), .ZN(n20824) );
  OA22X1 U21773 ( .IN1(n23022), .IN2(n19640), .IN3(n20824), .IN4(n19643), .Q(
        n19406) );
  INVX0 U21774 ( .INP(m0s4_data_i[12]), .ZN(n21421) );
  INVX0 U21775 ( .INP(m0s3_data_i[12]), .ZN(n23023) );
  OA22X1 U21776 ( .IN1(n21421), .IN2(n19632), .IN3(n23023), .IN4(n19633), .Q(
        n19405) );
  INVX0 U21777 ( .INP(m0s10_data_i[12]), .ZN(n21423) );
  INVX0 U21778 ( .INP(m0s0_data_i[12]), .ZN(n23019) );
  OA22X1 U21779 ( .IN1(n21423), .IN2(n19642), .IN3(n23019), .IN4(n19630), .Q(
        n19404) );
  NAND4X0 U21780 ( .IN1(n19407), .IN2(n19406), .IN3(n19405), .IN4(n19404), 
        .QN(n19408) );
  NOR2X0 U21781 ( .IN1(n19409), .IN2(n19408), .QN(n19411) );
  MUX21X1 U21782 ( .IN1(s15_data_i[12]), .IN2(\rf/rf_dout [12]), .S(n23501), 
        .Q(n23034) );
  NAND2X0 U21783 ( .IN1(n29312), .IN2(n23034), .QN(n19410) );
  NAND2X0 U21784 ( .IN1(n19411), .IN2(n19410), .QN(m4_data_o[12]) );
  INVX0 U21785 ( .INP(m0s1_data_i[13]), .ZN(n21433) );
  INVX0 U21786 ( .INP(m0s14_data_i[13]), .ZN(n23039) );
  OA22X1 U21787 ( .IN1(n21433), .IN2(n19646), .IN3(n23039), .IN4(n19617), .Q(
        n19415) );
  INVX0 U21788 ( .INP(m0s11_data_i[13]), .ZN(n23041) );
  INVX0 U21789 ( .INP(m0s12_data_i[13]), .ZN(n21435) );
  OA22X1 U21790 ( .IN1(n23041), .IN2(n19631), .IN3(n21435), .IN4(n19635), .Q(
        n19414) );
  INVX0 U21791 ( .INP(m0s2_data_i[13]), .ZN(n23040) );
  INVX0 U21792 ( .INP(m0s3_data_i[13]), .ZN(n22793) );
  OA22X1 U21793 ( .IN1(n23040), .IN2(n19634), .IN3(n22793), .IN4(n19633), .Q(
        n19413) );
  NAND2X0 U21794 ( .IN1(m0s8_data_i[13]), .IN2(n29319), .QN(n19412) );
  NAND4X0 U21795 ( .IN1(n19415), .IN2(n19414), .IN3(n19413), .IN4(n19412), 
        .QN(n19421) );
  INVX0 U21796 ( .INP(m0s6_data_i[13]), .ZN(n21436) );
  INVX0 U21797 ( .INP(m0s0_data_i[13]), .ZN(n23042) );
  OA22X1 U21798 ( .IN1(n21436), .IN2(n19643), .IN3(n23042), .IN4(n19630), .Q(
        n19419) );
  INVX0 U21799 ( .INP(m0s4_data_i[13]), .ZN(n21441) );
  INVX0 U21800 ( .INP(m0s5_data_i[13]), .ZN(n21432) );
  OA22X1 U21801 ( .IN1(n21441), .IN2(n19632), .IN3(n21432), .IN4(n19647), .Q(
        n19418) );
  INVX0 U21802 ( .INP(m0s7_data_i[13]), .ZN(n21443) );
  INVX0 U21803 ( .INP(m0s10_data_i[13]), .ZN(n23044) );
  OA22X1 U21804 ( .IN1(n21443), .IN2(n19645), .IN3(n23044), .IN4(n19642), .Q(
        n19417) );
  INVX0 U21805 ( .INP(m0s13_data_i[13]), .ZN(n21434) );
  INVX0 U21806 ( .INP(m0s9_data_i[13]), .ZN(n23043) );
  OA22X1 U21807 ( .IN1(n21434), .IN2(n19641), .IN3(n23043), .IN4(n19640), .Q(
        n19416) );
  NAND4X0 U21808 ( .IN1(n19419), .IN2(n19418), .IN3(n19417), .IN4(n19416), 
        .QN(n19420) );
  NOR2X0 U21809 ( .IN1(n19421), .IN2(n19420), .QN(n19423) );
  MUX21X1 U21810 ( .IN1(s15_data_i[13]), .IN2(\rf/rf_dout [13]), .S(n23501), 
        .Q(n23053) );
  NAND2X0 U21811 ( .IN1(n29312), .IN2(n23053), .QN(n19422) );
  NAND2X0 U21812 ( .IN1(n19423), .IN2(n19422), .QN(m4_data_o[13]) );
  INVX0 U21813 ( .INP(m0s4_data_i[14]), .ZN(n23064) );
  INVX0 U21814 ( .INP(m0s5_data_i[14]), .ZN(n21452) );
  OA22X1 U21815 ( .IN1(n23064), .IN2(n19632), .IN3(n21452), .IN4(n19647), .Q(
        n19427) );
  INVX0 U21816 ( .INP(m0s7_data_i[14]), .ZN(n21457) );
  INVX0 U21817 ( .INP(m0s12_data_i[14]), .ZN(n21458) );
  OA22X1 U21818 ( .IN1(n21457), .IN2(n19645), .IN3(n21458), .IN4(n19635), .Q(
        n19426) );
  INVX0 U21819 ( .INP(m0s2_data_i[14]), .ZN(n23060) );
  INVX0 U21820 ( .INP(m0s11_data_i[14]), .ZN(n23068) );
  OA22X1 U21821 ( .IN1(n23060), .IN2(n19634), .IN3(n23068), .IN4(n19631), .Q(
        n19425) );
  NAND2X0 U21822 ( .IN1(m0s3_data_i[14]), .IN2(n29324), .QN(n19424) );
  NAND4X0 U21823 ( .IN1(n19427), .IN2(n19426), .IN3(n19425), .IN4(n19424), 
        .QN(n19433) );
  INVX0 U21824 ( .INP(m0s6_data_i[14]), .ZN(n21460) );
  INVX0 U21825 ( .INP(m0s13_data_i[14]), .ZN(n20849) );
  OA22X1 U21826 ( .IN1(n21460), .IN2(n19643), .IN3(n20849), .IN4(n19641), .Q(
        n19431) );
  INVX0 U21827 ( .INP(m0s1_data_i[14]), .ZN(n23061) );
  INVX0 U21828 ( .INP(m0s10_data_i[14]), .ZN(n21461) );
  OA22X1 U21829 ( .IN1(n23061), .IN2(n19646), .IN3(n21461), .IN4(n19642), .Q(
        n19430) );
  INVX0 U21830 ( .INP(m0s0_data_i[14]), .ZN(n23066) );
  INVX0 U21831 ( .INP(m0s8_data_i[14]), .ZN(n23062) );
  OA22X1 U21832 ( .IN1(n23066), .IN2(n19630), .IN3(n23062), .IN4(n19644), .Q(
        n19429) );
  INVX0 U21833 ( .INP(m0s9_data_i[14]), .ZN(n23058) );
  INVX0 U21834 ( .INP(m0s14_data_i[14]), .ZN(n23070) );
  OA22X1 U21835 ( .IN1(n23058), .IN2(n19640), .IN3(n23070), .IN4(n19617), .Q(
        n19428) );
  NAND4X0 U21836 ( .IN1(n19431), .IN2(n19430), .IN3(n19429), .IN4(n19428), 
        .QN(n19432) );
  NOR2X0 U21837 ( .IN1(n19433), .IN2(n19432), .QN(n19435) );
  MUX21X1 U21838 ( .IN1(s15_data_i[14]), .IN2(\rf/rf_dout [14]), .S(n23501), 
        .Q(n23078) );
  NAND2X0 U21839 ( .IN1(n29312), .IN2(n23078), .QN(n19434) );
  NAND2X0 U21840 ( .IN1(n19435), .IN2(n19434), .QN(m4_data_o[14]) );
  INVX0 U21841 ( .INP(m0s14_data_i[15]), .ZN(n21481) );
  INVX0 U21842 ( .INP(m0s11_data_i[15]), .ZN(n21478) );
  OA22X1 U21843 ( .IN1(n21481), .IN2(n19617), .IN3(n21478), .IN4(n19631), .Q(
        n19439) );
  INVX0 U21844 ( .INP(m0s3_data_i[15]), .ZN(n23090) );
  INVX0 U21845 ( .INP(m0s13_data_i[15]), .ZN(n20862) );
  OA22X1 U21846 ( .IN1(n23090), .IN2(n19633), .IN3(n20862), .IN4(n19641), .Q(
        n19438) );
  INVX0 U21847 ( .INP(m0s10_data_i[15]), .ZN(n23084) );
  INVX0 U21848 ( .INP(m0s12_data_i[15]), .ZN(n23088) );
  OA22X1 U21849 ( .IN1(n23084), .IN2(n19642), .IN3(n23088), .IN4(n19635), .Q(
        n19437) );
  NAND2X0 U21850 ( .IN1(m0s2_data_i[15]), .IN2(n29325), .QN(n19436) );
  NAND4X0 U21851 ( .IN1(n19439), .IN2(n19438), .IN3(n19437), .IN4(n19436), 
        .QN(n19445) );
  INVX0 U21852 ( .INP(m0s8_data_i[15]), .ZN(n23092) );
  INVX0 U21853 ( .INP(m0s4_data_i[15]), .ZN(n21480) );
  OA22X1 U21854 ( .IN1(n23092), .IN2(n19644), .IN3(n21480), .IN4(n19632), .Q(
        n19443) );
  INVX0 U21855 ( .INP(m0s1_data_i[15]), .ZN(n23086) );
  INVX0 U21856 ( .INP(m0s0_data_i[15]), .ZN(n21477) );
  OA22X1 U21857 ( .IN1(n23086), .IN2(n19646), .IN3(n21477), .IN4(n19630), .Q(
        n19442) );
  INVX0 U21858 ( .INP(m0s9_data_i[15]), .ZN(n21471) );
  INVX0 U21859 ( .INP(m0s5_data_i[15]), .ZN(n21472) );
  OA22X1 U21860 ( .IN1(n21471), .IN2(n19640), .IN3(n21472), .IN4(n19647), .Q(
        n19441) );
  INVX0 U21861 ( .INP(m0s7_data_i[15]), .ZN(n23094) );
  INVX0 U21862 ( .INP(m0s6_data_i[15]), .ZN(n21479) );
  OA22X1 U21863 ( .IN1(n23094), .IN2(n19645), .IN3(n21479), .IN4(n19643), .Q(
        n19440) );
  NAND4X0 U21864 ( .IN1(n19443), .IN2(n19442), .IN3(n19441), .IN4(n19440), 
        .QN(n19444) );
  NOR2X0 U21865 ( .IN1(n19445), .IN2(n19444), .QN(n19447) );
  MUX21X1 U21866 ( .IN1(s15_data_i[15]), .IN2(\rf/rf_dout [15]), .S(n23501), 
        .Q(n23103) );
  NAND2X0 U21867 ( .IN1(n29312), .IN2(n23103), .QN(n19446) );
  NAND2X0 U21868 ( .IN1(n19447), .IN2(n19446), .QN(m4_data_o[15]) );
  INVX0 U21869 ( .INP(m0s12_data_i[16]), .ZN(n22012) );
  INVX0 U21870 ( .INP(m0s14_data_i[16]), .ZN(n21492) );
  OA22X1 U21871 ( .IN1(n19635), .IN2(n22012), .IN3(n19617), .IN4(n21492), .Q(
        n19451) );
  INVX0 U21872 ( .INP(m0s11_data_i[16]), .ZN(n22011) );
  INVX0 U21873 ( .INP(m0s3_data_i[16]), .ZN(n21491) );
  OA22X1 U21874 ( .IN1(n19631), .IN2(n22011), .IN3(n19633), .IN4(n21491), .Q(
        n19450) );
  INVX0 U21875 ( .INP(m0s6_data_i[16]), .ZN(n21502) );
  INVX0 U21876 ( .INP(m0s1_data_i[16]), .ZN(n21503) );
  OA22X1 U21877 ( .IN1(n19643), .IN2(n21502), .IN3(n19646), .IN4(n21503), .Q(
        n19449) );
  NAND2X0 U21878 ( .IN1(n29314), .IN2(m0s13_data_i[16]), .QN(n19448) );
  NAND4X0 U21879 ( .IN1(n19451), .IN2(n19450), .IN3(n19449), .IN4(n19448), 
        .QN(n19457) );
  INVX0 U21880 ( .INP(m0s0_data_i[16]), .ZN(n20879) );
  INVX0 U21881 ( .INP(m0s8_data_i[16]), .ZN(n21499) );
  OA22X1 U21882 ( .IN1(n19630), .IN2(n20879), .IN3(n19644), .IN4(n21499), .Q(
        n19455) );
  INVX0 U21883 ( .INP(m0s9_data_i[16]), .ZN(n21493) );
  INVX0 U21884 ( .INP(m0s10_data_i[16]), .ZN(n21501) );
  OA22X1 U21885 ( .IN1(n19640), .IN2(n21493), .IN3(n19642), .IN4(n21501), .Q(
        n19454) );
  INVX0 U21886 ( .INP(m0s2_data_i[16]), .ZN(n21490) );
  INVX0 U21887 ( .INP(m0s5_data_i[16]), .ZN(n22009) );
  OA22X1 U21888 ( .IN1(n19634), .IN2(n21490), .IN3(n19647), .IN4(n22009), .Q(
        n19453) );
  INVX0 U21889 ( .INP(m0s4_data_i[16]), .ZN(n21494) );
  INVX0 U21890 ( .INP(m0s7_data_i[16]), .ZN(n21500) );
  OA22X1 U21891 ( .IN1(n19632), .IN2(n21494), .IN3(n19645), .IN4(n21500), .Q(
        n19452) );
  NAND4X0 U21892 ( .IN1(n19455), .IN2(n19454), .IN3(n19453), .IN4(n19452), 
        .QN(n19456) );
  NOR2X0 U21893 ( .IN1(n19457), .IN2(n19456), .QN(n19460) );
  NOR2X0 U21894 ( .IN1(n23501), .IN2(n19458), .QN(n19654) );
  NAND2X0 U21895 ( .IN1(s15_data_i[16]), .IN2(n19654), .QN(n19459) );
  NAND2X0 U21896 ( .IN1(n19460), .IN2(n19459), .QN(m4_data_o[16]) );
  INVX0 U21897 ( .INP(m0s10_data_i[17]), .ZN(n22834) );
  INVX0 U21898 ( .INP(m0s7_data_i[17]), .ZN(n22831) );
  OA22X1 U21899 ( .IN1(n19642), .IN2(n22834), .IN3(n19645), .IN4(n22831), .Q(
        n19464) );
  INVX0 U21900 ( .INP(m0s2_data_i[17]), .ZN(n21512) );
  INVX0 U21901 ( .INP(m0s5_data_i[17]), .ZN(n21513) );
  OA22X1 U21902 ( .IN1(n19634), .IN2(n21512), .IN3(n19647), .IN4(n21513), .Q(
        n19463) );
  INVX0 U21903 ( .INP(m0s6_data_i[17]), .ZN(n21521) );
  INVX0 U21904 ( .INP(m0s8_data_i[17]), .ZN(n22397) );
  OA22X1 U21905 ( .IN1(n19643), .IN2(n21521), .IN3(n19644), .IN4(n22397), .Q(
        n19462) );
  NAND2X0 U21906 ( .IN1(n29315), .IN2(m0s12_data_i[17]), .QN(n19461) );
  NAND4X0 U21907 ( .IN1(n19464), .IN2(n19463), .IN3(n19462), .IN4(n19461), 
        .QN(n19470) );
  INVX0 U21908 ( .INP(m0s11_data_i[17]), .ZN(n22832) );
  INVX0 U21909 ( .INP(m0s9_data_i[17]), .ZN(n22835) );
  OA22X1 U21910 ( .IN1(n19631), .IN2(n22832), .IN3(n19640), .IN4(n22835), .Q(
        n19468) );
  INVX0 U21911 ( .INP(m0s4_data_i[17]), .ZN(n22833) );
  INVX0 U21912 ( .INP(m0s1_data_i[17]), .ZN(n21518) );
  OA22X1 U21913 ( .IN1(n19632), .IN2(n22833), .IN3(n19646), .IN4(n21518), .Q(
        n19467) );
  INVX0 U21914 ( .INP(m0s13_data_i[17]), .ZN(n22836) );
  INVX0 U21915 ( .INP(m0s0_data_i[17]), .ZN(n21520) );
  OA22X1 U21916 ( .IN1(n19641), .IN2(n22836), .IN3(n19630), .IN4(n21520), .Q(
        n19466) );
  INVX0 U21917 ( .INP(m0s3_data_i[17]), .ZN(n22830) );
  INVX0 U21918 ( .INP(m0s14_data_i[17]), .ZN(n21519) );
  OA22X1 U21919 ( .IN1(n19633), .IN2(n22830), .IN3(n19617), .IN4(n21519), .Q(
        n19465) );
  NAND4X0 U21920 ( .IN1(n19468), .IN2(n19467), .IN3(n19466), .IN4(n19465), 
        .QN(n19469) );
  NOR2X0 U21921 ( .IN1(n19470), .IN2(n19469), .QN(n19472) );
  NAND2X0 U21922 ( .IN1(s15_data_i[17]), .IN2(n19654), .QN(n19471) );
  NAND2X0 U21923 ( .IN1(n19472), .IN2(n19471), .QN(m4_data_o[17]) );
  INVX0 U21924 ( .INP(m0s9_data_i[18]), .ZN(n21530) );
  INVX0 U21925 ( .INP(m0s2_data_i[18]), .ZN(n21538) );
  OA22X1 U21926 ( .IN1(n19640), .IN2(n21530), .IN3(n19634), .IN4(n21538), .Q(
        n19476) );
  INVX0 U21927 ( .INP(m0s4_data_i[18]), .ZN(n21536) );
  INVX0 U21928 ( .INP(m0s14_data_i[18]), .ZN(n20901) );
  OA22X1 U21929 ( .IN1(n19632), .IN2(n21536), .IN3(n19617), .IN4(n20901), .Q(
        n19475) );
  INVX0 U21930 ( .INP(m0s0_data_i[18]), .ZN(n22415) );
  INVX0 U21931 ( .INP(m0s1_data_i[18]), .ZN(n22037) );
  OA22X1 U21932 ( .IN1(n19630), .IN2(n22415), .IN3(n19646), .IN4(n22037), .Q(
        n19474) );
  NAND2X0 U21933 ( .IN1(n29321), .IN2(m0s6_data_i[18]), .QN(n19473) );
  NAND4X0 U21934 ( .IN1(n19476), .IN2(n19475), .IN3(n19474), .IN4(n19473), 
        .QN(n19482) );
  INVX0 U21935 ( .INP(m0s3_data_i[18]), .ZN(n22413) );
  INVX0 U21936 ( .INP(m0s10_data_i[18]), .ZN(n21540) );
  OA22X1 U21937 ( .IN1(n19633), .IN2(n22413), .IN3(n19642), .IN4(n21540), .Q(
        n19480) );
  INVX0 U21938 ( .INP(m0s12_data_i[18]), .ZN(n22410) );
  INVX0 U21939 ( .INP(m0s7_data_i[18]), .ZN(n22411) );
  OA22X1 U21940 ( .IN1(n19635), .IN2(n22410), .IN3(n19645), .IN4(n22411), .Q(
        n19479) );
  INVX0 U21941 ( .INP(m0s11_data_i[18]), .ZN(n21537) );
  INVX0 U21942 ( .INP(m0s5_data_i[18]), .ZN(n22414) );
  OA22X1 U21943 ( .IN1(n19631), .IN2(n21537), .IN3(n19647), .IN4(n22414), .Q(
        n19478) );
  INVX0 U21944 ( .INP(m0s13_data_i[18]), .ZN(n21539) );
  INVX0 U21945 ( .INP(m0s8_data_i[18]), .ZN(n21531) );
  OA22X1 U21946 ( .IN1(n19641), .IN2(n21539), .IN3(n19644), .IN4(n21531), .Q(
        n19477) );
  NAND4X0 U21947 ( .IN1(n19480), .IN2(n19479), .IN3(n19478), .IN4(n19477), 
        .QN(n19481) );
  NOR2X0 U21948 ( .IN1(n19482), .IN2(n19481), .QN(n19484) );
  NAND2X0 U21949 ( .IN1(s15_data_i[18]), .IN2(n19654), .QN(n19483) );
  NAND2X0 U21950 ( .IN1(n19484), .IN2(n19483), .QN(m4_data_o[18]) );
  INVX0 U21951 ( .INP(m0s5_data_i[19]), .ZN(n22050) );
  INVX0 U21952 ( .INP(m0s1_data_i[19]), .ZN(n21557) );
  OA22X1 U21953 ( .IN1(n19647), .IN2(n22050), .IN3(n19646), .IN4(n21557), .Q(
        n19488) );
  INVX0 U21954 ( .INP(m0s4_data_i[19]), .ZN(n21556) );
  INVX0 U21955 ( .INP(m0s8_data_i[19]), .ZN(n21550) );
  OA22X1 U21956 ( .IN1(n19632), .IN2(n21556), .IN3(n19644), .IN4(n21550), .Q(
        n19487) );
  INVX0 U21957 ( .INP(m0s6_data_i[19]), .ZN(n21551) );
  INVX0 U21958 ( .INP(m0s7_data_i[19]), .ZN(n22435) );
  OA22X1 U21959 ( .IN1(n19643), .IN2(n21551), .IN3(n19645), .IN4(n22435), .Q(
        n19486) );
  NAND2X0 U21960 ( .IN1(n29314), .IN2(m0s13_data_i[19]), .QN(n19485) );
  NAND4X0 U21961 ( .IN1(n19488), .IN2(n19487), .IN3(n19486), .IN4(n19485), 
        .QN(n19494) );
  INVX0 U21962 ( .INP(m0s9_data_i[19]), .ZN(n22429) );
  INVX0 U21963 ( .INP(m0s14_data_i[19]), .ZN(n22428) );
  OA22X1 U21964 ( .IN1(n19640), .IN2(n22429), .IN3(n19617), .IN4(n22428), .Q(
        n19492) );
  INVX0 U21965 ( .INP(m0s11_data_i[19]), .ZN(n21549) );
  INVX0 U21966 ( .INP(m0s2_data_i[19]), .ZN(n21558) );
  OA22X1 U21967 ( .IN1(n19631), .IN2(n21549), .IN3(n19634), .IN4(n21558), .Q(
        n19491) );
  INVX0 U21968 ( .INP(m0s0_data_i[19]), .ZN(n22433) );
  INVX0 U21969 ( .INP(m0s10_data_i[19]), .ZN(n22432) );
  OA22X1 U21970 ( .IN1(n19630), .IN2(n22433), .IN3(n19642), .IN4(n22432), .Q(
        n19490) );
  INVX0 U21971 ( .INP(m0s3_data_i[19]), .ZN(n22431) );
  INVX0 U21972 ( .INP(m0s12_data_i[19]), .ZN(n22434) );
  OA22X1 U21973 ( .IN1(n19633), .IN2(n22431), .IN3(n19635), .IN4(n22434), .Q(
        n19489) );
  NAND4X0 U21974 ( .IN1(n19492), .IN2(n19491), .IN3(n19490), .IN4(n19489), 
        .QN(n19493) );
  NOR2X0 U21975 ( .IN1(n19494), .IN2(n19493), .QN(n19496) );
  NAND2X0 U21976 ( .IN1(s15_data_i[19]), .IN2(n19654), .QN(n19495) );
  NAND2X0 U21977 ( .IN1(n19496), .IN2(n19495), .QN(m4_data_o[19]) );
  INVX0 U21978 ( .INP(m0s12_data_i[20]), .ZN(n22449) );
  INVX0 U21979 ( .INP(m0s10_data_i[20]), .ZN(n21574) );
  OA22X1 U21980 ( .IN1(n19635), .IN2(n22449), .IN3(n19642), .IN4(n21574), .Q(
        n19500) );
  INVX0 U21981 ( .INP(m0s13_data_i[20]), .ZN(n21567) );
  INVX0 U21982 ( .INP(m0s5_data_i[20]), .ZN(n22448) );
  OA22X1 U21983 ( .IN1(n19641), .IN2(n21567), .IN3(n19647), .IN4(n22448), .Q(
        n19499) );
  INVX0 U21984 ( .INP(m0s4_data_i[20]), .ZN(n21577) );
  INVX0 U21985 ( .INP(m0s6_data_i[20]), .ZN(n22454) );
  OA22X1 U21986 ( .IN1(n19632), .IN2(n21577), .IN3(n19643), .IN4(n22454), .Q(
        n19498) );
  NAND2X0 U21987 ( .IN1(n29313), .IN2(m0s14_data_i[20]), .QN(n19497) );
  NAND4X0 U21988 ( .IN1(n19500), .IN2(n19499), .IN3(n19498), .IN4(n19497), 
        .QN(n19506) );
  INVX0 U21989 ( .INP(m0s3_data_i[20]), .ZN(n21568) );
  INVX0 U21990 ( .INP(m0s1_data_i[20]), .ZN(n21575) );
  OA22X1 U21991 ( .IN1(n19633), .IN2(n21568), .IN3(n19646), .IN4(n21575), .Q(
        n19504) );
  INVX0 U21992 ( .INP(m0s9_data_i[20]), .ZN(n22447) );
  INVX0 U21993 ( .INP(m0s7_data_i[20]), .ZN(n21576) );
  OA22X1 U21994 ( .IN1(n19640), .IN2(n22447), .IN3(n19645), .IN4(n21576), .Q(
        n19503) );
  INVX0 U21995 ( .INP(m0s11_data_i[20]), .ZN(n22450) );
  INVX0 U21996 ( .INP(m0s8_data_i[20]), .ZN(n21573) );
  OA22X1 U21997 ( .IN1(n19631), .IN2(n22450), .IN3(n19644), .IN4(n21573), .Q(
        n19502) );
  INVX0 U21998 ( .INP(m0s2_data_i[20]), .ZN(n22452) );
  INVX0 U21999 ( .INP(m0s0_data_i[20]), .ZN(n22451) );
  OA22X1 U22000 ( .IN1(n19634), .IN2(n22452), .IN3(n19630), .IN4(n22451), .Q(
        n19501) );
  NAND4X0 U22001 ( .IN1(n19504), .IN2(n19503), .IN3(n19502), .IN4(n19501), 
        .QN(n19505) );
  NOR2X0 U22002 ( .IN1(n19506), .IN2(n19505), .QN(n19508) );
  NAND2X0 U22003 ( .IN1(s15_data_i[20]), .IN2(n19654), .QN(n19507) );
  NAND2X0 U22004 ( .IN1(n19508), .IN2(n19507), .QN(m4_data_o[20]) );
  INVX0 U22005 ( .INP(m0s14_data_i[21]), .ZN(n21586) );
  INVX0 U22006 ( .INP(m0s7_data_i[21]), .ZN(n22857) );
  OA22X1 U22007 ( .IN1(n19617), .IN2(n21586), .IN3(n19645), .IN4(n22857), .Q(
        n19512) );
  INVX0 U22008 ( .INP(m0s3_data_i[21]), .ZN(n21593) );
  INVX0 U22009 ( .INP(m0s2_data_i[21]), .ZN(n22856) );
  OA22X1 U22010 ( .IN1(n19633), .IN2(n21593), .IN3(n19634), .IN4(n22856), .Q(
        n19511) );
  INVX0 U22011 ( .INP(m0s6_data_i[21]), .ZN(n22855) );
  INVX0 U22012 ( .INP(m0s1_data_i[21]), .ZN(n22466) );
  OA22X1 U22013 ( .IN1(n19643), .IN2(n22855), .IN3(n19646), .IN4(n22466), .Q(
        n19510) );
  NAND2X0 U22014 ( .IN1(n29323), .IN2(m0s4_data_i[21]), .QN(n19509) );
  NAND4X0 U22015 ( .IN1(n19512), .IN2(n19511), .IN3(n19510), .IN4(n19509), 
        .QN(n19518) );
  INVX0 U22016 ( .INP(m0s11_data_i[21]), .ZN(n20942) );
  INVX0 U22017 ( .INP(m0s13_data_i[21]), .ZN(n21587) );
  OA22X1 U22018 ( .IN1(n19631), .IN2(n20942), .IN3(n19641), .IN4(n21587), .Q(
        n19516) );
  INVX0 U22019 ( .INP(m0s12_data_i[21]), .ZN(n22852) );
  INVX0 U22020 ( .INP(m0s10_data_i[21]), .ZN(n22849) );
  OA22X1 U22021 ( .IN1(n19635), .IN2(n22852), .IN3(n19642), .IN4(n22849), .Q(
        n19515) );
  INVX0 U22022 ( .INP(m0s9_data_i[21]), .ZN(n21594) );
  INVX0 U22023 ( .INP(m0s8_data_i[21]), .ZN(n21592) );
  OA22X1 U22024 ( .IN1(n19640), .IN2(n21594), .IN3(n19644), .IN4(n21592), .Q(
        n19514) );
  INVX0 U22025 ( .INP(m0s5_data_i[21]), .ZN(n22851) );
  INVX0 U22026 ( .INP(m0s0_data_i[21]), .ZN(n22853) );
  OA22X1 U22027 ( .IN1(n19647), .IN2(n22851), .IN3(n19630), .IN4(n22853), .Q(
        n19513) );
  NAND4X0 U22028 ( .IN1(n19516), .IN2(n19515), .IN3(n19514), .IN4(n19513), 
        .QN(n19517) );
  NOR2X0 U22029 ( .IN1(n19518), .IN2(n19517), .QN(n19520) );
  NAND2X0 U22030 ( .IN1(s15_data_i[21]), .IN2(n19654), .QN(n19519) );
  NAND2X0 U22031 ( .IN1(n19520), .IN2(n19519), .QN(m4_data_o[21]) );
  INVX0 U22032 ( .INP(m0s11_data_i[22]), .ZN(n20951) );
  INVX0 U22033 ( .INP(m0s7_data_i[22]), .ZN(n22874) );
  OA22X1 U22034 ( .IN1(n19631), .IN2(n20951), .IN3(n19645), .IN4(n22874), .Q(
        n19524) );
  INVX0 U22035 ( .INP(m0s3_data_i[22]), .ZN(n22871) );
  INVX0 U22036 ( .INP(m0s2_data_i[22]), .ZN(n22870) );
  OA22X1 U22037 ( .IN1(n19633), .IN2(n22871), .IN3(n19634), .IN4(n22870), .Q(
        n19523) );
  INVX0 U22038 ( .INP(m0s4_data_i[22]), .ZN(n22876) );
  INVX0 U22039 ( .INP(m0s0_data_i[22]), .ZN(n21604) );
  OA22X1 U22040 ( .IN1(n19632), .IN2(n22876), .IN3(n19630), .IN4(n21604), .Q(
        n19522) );
  NAND2X0 U22041 ( .IN1(n29313), .IN2(m0s14_data_i[22]), .QN(n19521) );
  NAND4X0 U22042 ( .IN1(n19524), .IN2(n19523), .IN3(n19522), .IN4(n19521), 
        .QN(n19530) );
  INVX0 U22043 ( .INP(m0s13_data_i[22]), .ZN(n21611) );
  INVX0 U22044 ( .INP(m0s9_data_i[22]), .ZN(n21610) );
  OA22X1 U22045 ( .IN1(n19641), .IN2(n21611), .IN3(n19640), .IN4(n21610), .Q(
        n19528) );
  INVX0 U22046 ( .INP(m0s12_data_i[22]), .ZN(n22875) );
  INVX0 U22047 ( .INP(m0s1_data_i[22]), .ZN(n21612) );
  OA22X1 U22048 ( .IN1(n19635), .IN2(n22875), .IN3(n19646), .IN4(n21612), .Q(
        n19527) );
  INVX0 U22049 ( .INP(m0s10_data_i[22]), .ZN(n22869) );
  INVX0 U22050 ( .INP(m0s8_data_i[22]), .ZN(n22873) );
  OA22X1 U22051 ( .IN1(n19642), .IN2(n22869), .IN3(n19644), .IN4(n22873), .Q(
        n19526) );
  INVX0 U22052 ( .INP(m0s6_data_i[22]), .ZN(n22872) );
  INVX0 U22053 ( .INP(m0s5_data_i[22]), .ZN(n21609) );
  OA22X1 U22054 ( .IN1(n19643), .IN2(n22872), .IN3(n19647), .IN4(n21609), .Q(
        n19525) );
  NAND4X0 U22055 ( .IN1(n19528), .IN2(n19527), .IN3(n19526), .IN4(n19525), 
        .QN(n19529) );
  NOR2X0 U22056 ( .IN1(n19530), .IN2(n19529), .QN(n19532) );
  NAND2X0 U22057 ( .IN1(s15_data_i[22]), .IN2(n19654), .QN(n19531) );
  NAND2X0 U22058 ( .IN1(n19532), .IN2(n19531), .QN(m4_data_o[22]) );
  INVX0 U22059 ( .INP(m0s11_data_i[23]), .ZN(n21630) );
  INVX0 U22060 ( .INP(m0s2_data_i[23]), .ZN(n21623) );
  OA22X1 U22061 ( .IN1(n19631), .IN2(n21630), .IN3(n19634), .IN4(n21623), .Q(
        n19536) );
  INVX0 U22062 ( .INP(m0s5_data_i[23]), .ZN(n21624) );
  INVX0 U22063 ( .INP(m0s1_data_i[23]), .ZN(n22491) );
  OA22X1 U22064 ( .IN1(n19647), .IN2(n21624), .IN3(n19646), .IN4(n22491), .Q(
        n19535) );
  INVX0 U22065 ( .INP(m0s9_data_i[23]), .ZN(n21633) );
  INVX0 U22066 ( .INP(m0s6_data_i[23]), .ZN(n21625) );
  OA22X1 U22067 ( .IN1(n19640), .IN2(n21633), .IN3(n19643), .IN4(n21625), .Q(
        n19534) );
  NAND2X0 U22068 ( .IN1(n29328), .IN2(m0s0_data_i[23]), .QN(n19533) );
  NAND4X0 U22069 ( .IN1(n19536), .IN2(n19535), .IN3(n19534), .IN4(n19533), 
        .QN(n19542) );
  INVX0 U22070 ( .INP(m0s3_data_i[23]), .ZN(n21631) );
  INVX0 U22071 ( .INP(m0s10_data_i[23]), .ZN(n22494) );
  OA22X1 U22072 ( .IN1(n19633), .IN2(n21631), .IN3(n19642), .IN4(n22494), .Q(
        n19540) );
  INVX0 U22073 ( .INP(m0s4_data_i[23]), .ZN(n20968) );
  INVX0 U22074 ( .INP(m0s13_data_i[23]), .ZN(n21632) );
  OA22X1 U22075 ( .IN1(n19632), .IN2(n20968), .IN3(n19641), .IN4(n21632), .Q(
        n19539) );
  INVX0 U22076 ( .INP(m0s12_data_i[23]), .ZN(n21622) );
  INVX0 U22077 ( .INP(m0s8_data_i[23]), .ZN(n22492) );
  OA22X1 U22078 ( .IN1(n19635), .IN2(n21622), .IN3(n19644), .IN4(n22492), .Q(
        n19538) );
  INVX0 U22079 ( .INP(m0s14_data_i[23]), .ZN(n21621) );
  INVX0 U22080 ( .INP(m0s7_data_i[23]), .ZN(n22495) );
  OA22X1 U22081 ( .IN1(n19617), .IN2(n21621), .IN3(n19645), .IN4(n22495), .Q(
        n19537) );
  NAND4X0 U22082 ( .IN1(n19540), .IN2(n19539), .IN3(n19538), .IN4(n19537), 
        .QN(n19541) );
  NOR2X0 U22083 ( .IN1(n19542), .IN2(n19541), .QN(n19544) );
  NAND2X0 U22084 ( .IN1(s15_data_i[23]), .IN2(n19654), .QN(n19543) );
  NAND2X0 U22085 ( .IN1(n19544), .IN2(n19543), .QN(m4_data_o[23]) );
  INVX0 U22086 ( .INP(m0s9_data_i[24]), .ZN(n21650) );
  INVX0 U22087 ( .INP(m0s6_data_i[24]), .ZN(n22889) );
  OA22X1 U22088 ( .IN1(n19640), .IN2(n21650), .IN3(n19643), .IN4(n22889), .Q(
        n19548) );
  INVX0 U22089 ( .INP(m0s2_data_i[24]), .ZN(n22890) );
  INVX0 U22090 ( .INP(m0s14_data_i[24]), .ZN(n22893) );
  OA22X1 U22091 ( .IN1(n19634), .IN2(n22890), .IN3(n19617), .IN4(n22893), .Q(
        n19547) );
  INVX0 U22092 ( .INP(m0s4_data_i[24]), .ZN(n21644) );
  INVX0 U22093 ( .INP(m0s8_data_i[24]), .ZN(n21653) );
  OA22X1 U22094 ( .IN1(n19632), .IN2(n21644), .IN3(n19644), .IN4(n21653), .Q(
        n19546) );
  NAND2X0 U22095 ( .IN1(n29317), .IN2(m0s10_data_i[24]), .QN(n19545) );
  NAND4X0 U22096 ( .IN1(n19548), .IN2(n19547), .IN3(n19546), .IN4(n19545), 
        .QN(n19554) );
  INVX0 U22097 ( .INP(m0s3_data_i[24]), .ZN(n21643) );
  INVX0 U22098 ( .INP(m0s5_data_i[24]), .ZN(n22895) );
  OA22X1 U22099 ( .IN1(n19633), .IN2(n21643), .IN3(n19647), .IN4(n22895), .Q(
        n19552) );
  INVX0 U22100 ( .INP(m0s12_data_i[24]), .ZN(n21652) );
  INVX0 U22101 ( .INP(m0s1_data_i[24]), .ZN(n22896) );
  OA22X1 U22102 ( .IN1(n19635), .IN2(n21652), .IN3(n19646), .IN4(n22896), .Q(
        n19551) );
  INVX0 U22103 ( .INP(m0s13_data_i[24]), .ZN(n22888) );
  INVX0 U22104 ( .INP(m0s0_data_i[24]), .ZN(n21649) );
  OA22X1 U22105 ( .IN1(n19641), .IN2(n22888), .IN3(n19630), .IN4(n21649), .Q(
        n19550) );
  INVX0 U22106 ( .INP(m0s11_data_i[24]), .ZN(n21651) );
  INVX0 U22107 ( .INP(m0s7_data_i[24]), .ZN(n22891) );
  OA22X1 U22108 ( .IN1(n19631), .IN2(n21651), .IN3(n19645), .IN4(n22891), .Q(
        n19549) );
  NAND4X0 U22109 ( .IN1(n19552), .IN2(n19551), .IN3(n19550), .IN4(n19549), 
        .QN(n19553) );
  NOR2X0 U22110 ( .IN1(n19554), .IN2(n19553), .QN(n19556) );
  NAND2X0 U22111 ( .IN1(s15_data_i[24]), .IN2(n19654), .QN(n19555) );
  NAND2X0 U22112 ( .IN1(n19556), .IN2(n19555), .QN(m4_data_o[24]) );
  INVX0 U22113 ( .INP(m0s9_data_i[25]), .ZN(n22520) );
  INVX0 U22114 ( .INP(m0s1_data_i[25]), .ZN(n21662) );
  OA22X1 U22115 ( .IN1(n19640), .IN2(n22520), .IN3(n19646), .IN4(n21662), .Q(
        n19560) );
  INVX0 U22116 ( .INP(m0s0_data_i[25]), .ZN(n21664) );
  INVX0 U22117 ( .INP(m0s7_data_i[25]), .ZN(n21672) );
  OA22X1 U22118 ( .IN1(n19630), .IN2(n21664), .IN3(n19645), .IN4(n21672), .Q(
        n19559) );
  INVX0 U22119 ( .INP(m0s3_data_i[25]), .ZN(n22521) );
  INVX0 U22120 ( .INP(m0s2_data_i[25]), .ZN(n21663) );
  OA22X1 U22121 ( .IN1(n19633), .IN2(n22521), .IN3(n19634), .IN4(n21663), .Q(
        n19558) );
  NAND2X0 U22122 ( .IN1(n29322), .IN2(m0s5_data_i[25]), .QN(n19557) );
  NAND4X0 U22123 ( .IN1(n19560), .IN2(n19559), .IN3(n19558), .IN4(n19557), 
        .QN(n19566) );
  INVX0 U22124 ( .INP(m0s11_data_i[25]), .ZN(n21670) );
  INVX0 U22125 ( .INP(m0s8_data_i[25]), .ZN(n21671) );
  OA22X1 U22126 ( .IN1(n19631), .IN2(n21670), .IN3(n19644), .IN4(n21671), .Q(
        n19564) );
  INVX0 U22127 ( .INP(m0s13_data_i[25]), .ZN(n20993) );
  INVX0 U22128 ( .INP(m0s6_data_i[25]), .ZN(n22119) );
  OA22X1 U22129 ( .IN1(n19641), .IN2(n20993), .IN3(n19643), .IN4(n22119), .Q(
        n19563) );
  INVX0 U22130 ( .INP(m0s4_data_i[25]), .ZN(n21665) );
  INVX0 U22131 ( .INP(m0s14_data_i[25]), .ZN(n22524) );
  OA22X1 U22132 ( .IN1(n19632), .IN2(n21665), .IN3(n19617), .IN4(n22524), .Q(
        n19562) );
  INVX0 U22133 ( .INP(m0s12_data_i[25]), .ZN(n22522) );
  INVX0 U22134 ( .INP(m0s10_data_i[25]), .ZN(n22523) );
  OA22X1 U22135 ( .IN1(n19635), .IN2(n22522), .IN3(n19642), .IN4(n22523), .Q(
        n19561) );
  NAND4X0 U22136 ( .IN1(n19564), .IN2(n19563), .IN3(n19562), .IN4(n19561), 
        .QN(n19565) );
  NOR2X0 U22137 ( .IN1(n19566), .IN2(n19565), .QN(n19568) );
  NAND2X0 U22138 ( .IN1(s15_data_i[25]), .IN2(n19654), .QN(n19567) );
  NAND2X0 U22139 ( .IN1(n19568), .IN2(n19567), .QN(m4_data_o[25]) );
  INVX0 U22140 ( .INP(m0s13_data_i[26]), .ZN(n21691) );
  INVX0 U22141 ( .INP(m0s10_data_i[26]), .ZN(n22540) );
  OA22X1 U22142 ( .IN1(n19641), .IN2(n21691), .IN3(n19642), .IN4(n22540), .Q(
        n19572) );
  INVX0 U22143 ( .INP(m0s3_data_i[26]), .ZN(n21694) );
  INVX0 U22144 ( .INP(m0s12_data_i[26]), .ZN(n21686) );
  OA22X1 U22145 ( .IN1(n19633), .IN2(n21694), .IN3(n19635), .IN4(n21686), .Q(
        n19571) );
  INVX0 U22146 ( .INP(m0s11_data_i[26]), .ZN(n22541) );
  INVX0 U22147 ( .INP(m0s6_data_i[26]), .ZN(n22539) );
  OA22X1 U22148 ( .IN1(n19631), .IN2(n22541), .IN3(n19643), .IN4(n22539), .Q(
        n19570) );
  NAND2X0 U22149 ( .IN1(n29319), .IN2(m0s8_data_i[26]), .QN(n19569) );
  NAND4X0 U22150 ( .IN1(n19572), .IN2(n19571), .IN3(n19570), .IN4(n19569), 
        .QN(n19578) );
  INVX0 U22151 ( .INP(m0s14_data_i[26]), .ZN(n21681) );
  INVX0 U22152 ( .INP(m0s1_data_i[26]), .ZN(n21695) );
  OA22X1 U22153 ( .IN1(n19617), .IN2(n21681), .IN3(n19646), .IN4(n21695), .Q(
        n19576) );
  INVX0 U22154 ( .INP(m0s4_data_i[26]), .ZN(n21685) );
  INVX0 U22155 ( .INP(m0s0_data_i[26]), .ZN(n21692) );
  OA22X1 U22156 ( .IN1(n19632), .IN2(n21685), .IN3(n19630), .IN4(n21692), .Q(
        n19575) );
  INVX0 U22157 ( .INP(m0s9_data_i[26]), .ZN(n21693) );
  INVX0 U22158 ( .INP(m0s5_data_i[26]), .ZN(n21684) );
  OA22X1 U22159 ( .IN1(n19640), .IN2(n21693), .IN3(n19647), .IN4(n21684), .Q(
        n19574) );
  INVX0 U22160 ( .INP(m0s2_data_i[26]), .ZN(n21682) );
  INVX0 U22161 ( .INP(m0s7_data_i[26]), .ZN(n21683) );
  OA22X1 U22162 ( .IN1(n19634), .IN2(n21682), .IN3(n19645), .IN4(n21683), .Q(
        n19573) );
  NAND4X0 U22163 ( .IN1(n19576), .IN2(n19575), .IN3(n19574), .IN4(n19573), 
        .QN(n19577) );
  NOR2X0 U22164 ( .IN1(n19578), .IN2(n19577), .QN(n19580) );
  NAND2X0 U22165 ( .IN1(s15_data_i[26]), .IN2(n19654), .QN(n19579) );
  NAND2X0 U22166 ( .IN1(n19580), .IN2(n19579), .QN(m4_data_o[26]) );
  INVX0 U22167 ( .INP(m0s13_data_i[27]), .ZN(n22918) );
  INVX0 U22168 ( .INP(m0s1_data_i[27]), .ZN(n22910) );
  OA22X1 U22169 ( .IN1(n19641), .IN2(n22918), .IN3(n19646), .IN4(n22910), .Q(
        n19584) );
  INVX0 U22170 ( .INP(m0s2_data_i[27]), .ZN(n22916) );
  INVX0 U22171 ( .INP(m0s14_data_i[27]), .ZN(n21710) );
  OA22X1 U22172 ( .IN1(n19634), .IN2(n22916), .IN3(n19617), .IN4(n21710), .Q(
        n19583) );
  INVX0 U22173 ( .INP(m0s11_data_i[27]), .ZN(n21713) );
  INVX0 U22174 ( .INP(m0s6_data_i[27]), .ZN(n21715) );
  OA22X1 U22175 ( .IN1(n19631), .IN2(n21713), .IN3(n19643), .IN4(n21715), .Q(
        n19582) );
  NAND2X0 U22176 ( .IN1(n29324), .IN2(m0s3_data_i[27]), .QN(n19581) );
  NAND4X0 U22177 ( .IN1(n19584), .IN2(n19583), .IN3(n19582), .IN4(n19581), 
        .QN(n19590) );
  INVX0 U22178 ( .INP(m0s10_data_i[27]), .ZN(n22911) );
  INVX0 U22179 ( .INP(m0s7_data_i[27]), .ZN(n22908) );
  OA22X1 U22180 ( .IN1(n19642), .IN2(n22911), .IN3(n19645), .IN4(n22908), .Q(
        n19588) );
  INVX0 U22181 ( .INP(m0s12_data_i[27]), .ZN(n22915) );
  INVX0 U22182 ( .INP(m0s5_data_i[27]), .ZN(n21705) );
  OA22X1 U22183 ( .IN1(n19635), .IN2(n22915), .IN3(n19647), .IN4(n21705), .Q(
        n19587) );
  INVX0 U22184 ( .INP(m0s9_data_i[27]), .ZN(n21714) );
  INVX0 U22185 ( .INP(m0s0_data_i[27]), .ZN(n21018) );
  OA22X1 U22186 ( .IN1(n19640), .IN2(n21714), .IN3(n19630), .IN4(n21018), .Q(
        n19586) );
  INVX0 U22187 ( .INP(m0s4_data_i[27]), .ZN(n21711) );
  INVX0 U22188 ( .INP(m0s8_data_i[27]), .ZN(n22913) );
  OA22X1 U22189 ( .IN1(n19632), .IN2(n21711), .IN3(n19644), .IN4(n22913), .Q(
        n19585) );
  NAND4X0 U22190 ( .IN1(n19588), .IN2(n19587), .IN3(n19586), .IN4(n19585), 
        .QN(n19589) );
  NOR2X0 U22191 ( .IN1(n19590), .IN2(n19589), .QN(n19592) );
  NAND2X0 U22192 ( .IN1(s15_data_i[27]), .IN2(n19654), .QN(n19591) );
  NAND2X0 U22193 ( .IN1(n19592), .IN2(n19591), .QN(m4_data_o[27]) );
  INVX0 U22194 ( .INP(m0s6_data_i[28]), .ZN(n22940) );
  INVX0 U22195 ( .INP(m0s1_data_i[28]), .ZN(n22941) );
  OA22X1 U22196 ( .IN1(n19643), .IN2(n22940), .IN3(n19646), .IN4(n22941), .Q(
        n19596) );
  INVX0 U22197 ( .INP(m0s3_data_i[28]), .ZN(n21743) );
  INVX0 U22198 ( .INP(m0s9_data_i[28]), .ZN(n22934) );
  OA22X1 U22199 ( .IN1(n19633), .IN2(n21743), .IN3(n19640), .IN4(n22934), .Q(
        n19595) );
  INVX0 U22200 ( .INP(m0s13_data_i[28]), .ZN(n22932) );
  INVX0 U22201 ( .INP(m0s2_data_i[28]), .ZN(n21741) );
  OA22X1 U22202 ( .IN1(n19641), .IN2(n22932), .IN3(n19634), .IN4(n21741), .Q(
        n19594) );
  NAND2X0 U22203 ( .IN1(n29317), .IN2(m0s10_data_i[28]), .QN(n19593) );
  NAND4X0 U22204 ( .IN1(n19596), .IN2(n19595), .IN3(n19594), .IN4(n19593), 
        .QN(n19602) );
  INVX0 U22205 ( .INP(m0s11_data_i[28]), .ZN(n22930) );
  INVX0 U22206 ( .INP(m0s14_data_i[28]), .ZN(n21725) );
  OA22X1 U22207 ( .IN1(n19631), .IN2(n22930), .IN3(n19617), .IN4(n21725), .Q(
        n19600) );
  INVX0 U22208 ( .INP(m0s0_data_i[28]), .ZN(n22568) );
  INVX0 U22209 ( .INP(m0s8_data_i[28]), .ZN(n21739) );
  OA22X1 U22210 ( .IN1(n19630), .IN2(n22568), .IN3(n19644), .IN4(n21739), .Q(
        n19599) );
  INVX0 U22211 ( .INP(m0s12_data_i[28]), .ZN(n22935) );
  INVX0 U22212 ( .INP(m0s5_data_i[28]), .ZN(n22936) );
  OA22X1 U22213 ( .IN1(n19635), .IN2(n22935), .IN3(n19647), .IN4(n22936), .Q(
        n19598) );
  INVX0 U22214 ( .INP(m0s4_data_i[28]), .ZN(n22938) );
  INVX0 U22215 ( .INP(m0s7_data_i[28]), .ZN(n21737) );
  OA22X1 U22216 ( .IN1(n19632), .IN2(n22938), .IN3(n19645), .IN4(n21737), .Q(
        n19597) );
  NAND4X0 U22217 ( .IN1(n19600), .IN2(n19599), .IN3(n19598), .IN4(n19597), 
        .QN(n19601) );
  NOR2X0 U22218 ( .IN1(n19602), .IN2(n19601), .QN(n19604) );
  NAND2X0 U22219 ( .IN1(s15_data_i[28]), .IN2(n19654), .QN(n19603) );
  NAND2X0 U22220 ( .IN1(n19604), .IN2(n19603), .QN(m4_data_o[28]) );
  INVX0 U22221 ( .INP(m0s3_data_i[29]), .ZN(n22953) );
  INVX0 U22222 ( .INP(m0s4_data_i[29]), .ZN(n21051) );
  OA22X1 U22223 ( .IN1(n19633), .IN2(n22953), .IN3(n19632), .IN4(n21051), .Q(
        n19608) );
  INVX0 U22224 ( .INP(m0s9_data_i[29]), .ZN(n22955) );
  INVX0 U22225 ( .INP(m0s2_data_i[29]), .ZN(n21049) );
  OA22X1 U22226 ( .IN1(n19640), .IN2(n22955), .IN3(n19634), .IN4(n21049), .Q(
        n19607) );
  INVX0 U22227 ( .INP(m0s11_data_i[29]), .ZN(n21042) );
  INVX0 U22228 ( .INP(m0s6_data_i[29]), .ZN(n22963) );
  OA22X1 U22229 ( .IN1(n19631), .IN2(n21042), .IN3(n19643), .IN4(n22963), .Q(
        n19606) );
  NAND2X0 U22230 ( .IN1(n29322), .IN2(m0s5_data_i[29]), .QN(n19605) );
  NAND4X0 U22231 ( .IN1(n19608), .IN2(n19607), .IN3(n19606), .IN4(n19605), 
        .QN(n19614) );
  INVX0 U22232 ( .INP(m0s12_data_i[29]), .ZN(n22957) );
  INVX0 U22233 ( .INP(m0s1_data_i[29]), .ZN(n22959) );
  OA22X1 U22234 ( .IN1(n19635), .IN2(n22957), .IN3(n19646), .IN4(n22959), .Q(
        n19612) );
  INVX0 U22235 ( .INP(m0s13_data_i[29]), .ZN(n21041) );
  INVX0 U22236 ( .INP(m0s10_data_i[29]), .ZN(n22961) );
  OA22X1 U22237 ( .IN1(n19641), .IN2(n21041), .IN3(n19642), .IN4(n22961), .Q(
        n19611) );
  INVX0 U22238 ( .INP(m0s14_data_i[29]), .ZN(n21050) );
  INVX0 U22239 ( .INP(m0s7_data_i[29]), .ZN(n22583) );
  OA22X1 U22240 ( .IN1(n19617), .IN2(n21050), .IN3(n19645), .IN4(n22583), .Q(
        n19610) );
  INVX0 U22241 ( .INP(m0s0_data_i[29]), .ZN(n21043) );
  INVX0 U22242 ( .INP(m0s8_data_i[29]), .ZN(n21048) );
  OA22X1 U22243 ( .IN1(n19630), .IN2(n21043), .IN3(n19644), .IN4(n21048), .Q(
        n19609) );
  NAND4X0 U22244 ( .IN1(n19612), .IN2(n19611), .IN3(n19610), .IN4(n19609), 
        .QN(n19613) );
  NOR2X0 U22245 ( .IN1(n19614), .IN2(n19613), .QN(n19616) );
  NAND2X0 U22246 ( .IN1(s15_data_i[29]), .IN2(n19654), .QN(n19615) );
  NAND2X0 U22247 ( .IN1(n19616), .IN2(n19615), .QN(m4_data_o[29]) );
  OA22X1 U22248 ( .IN1(n19632), .IN2(n21069), .IN3(n19641), .IN4(n22602), .Q(
        n19621) );
  OA22X1 U22249 ( .IN1(n19633), .IN2(n21070), .IN3(n19643), .IN4(n21071), .Q(
        n19620) );
  OA22X1 U22250 ( .IN1(n19634), .IN2(n22603), .IN3(n19617), .IN4(n22597), .Q(
        n19619) );
  NAND2X0 U22251 ( .IN1(n29318), .IN2(m0s9_data_i[30]), .QN(n19618) );
  NAND4X0 U22252 ( .IN1(n19621), .IN2(n19620), .IN3(n19619), .IN4(n19618), 
        .QN(n19627) );
  OA22X1 U22253 ( .IN1(n19635), .IN2(n22600), .IN3(n19642), .IN4(n22598), .Q(
        n19625) );
  OA22X1 U22254 ( .IN1(n19647), .IN2(n21072), .IN3(n19644), .IN4(n21061), .Q(
        n19624) );
  OA22X1 U22255 ( .IN1(n19645), .IN2(n21060), .IN3(n19646), .IN4(n22601), .Q(
        n19623) );
  OA22X1 U22256 ( .IN1(n19631), .IN2(n21062), .IN3(n19630), .IN4(n22177), .Q(
        n19622) );
  NAND4X0 U22257 ( .IN1(n19625), .IN2(n19624), .IN3(n19623), .IN4(n19622), 
        .QN(n19626) );
  NOR2X0 U22258 ( .IN1(n19627), .IN2(n19626), .QN(n19629) );
  NAND2X0 U22259 ( .IN1(s15_data_i[30]), .IN2(n19654), .QN(n19628) );
  NAND2X0 U22260 ( .IN1(n19629), .IN2(n19628), .QN(m4_data_o[30]) );
  OA22X1 U22261 ( .IN1(n19631), .IN2(n21086), .IN3(n19630), .IN4(n21107), .Q(
        n19639) );
  OA22X1 U22262 ( .IN1(n19633), .IN2(n22617), .IN3(n19632), .IN4(n21105), .Q(
        n19638) );
  INVX0 U22263 ( .INP(m0s12_data_i[31]), .ZN(n21097) );
  OA22X1 U22264 ( .IN1(n19635), .IN2(n21097), .IN3(n19634), .IN4(n22619), .Q(
        n19637) );
  NAND2X0 U22265 ( .IN1(n29313), .IN2(m0s14_data_i[31]), .QN(n19636) );
  NAND4X0 U22266 ( .IN1(n19639), .IN2(n19638), .IN3(n19637), .IN4(n19636), 
        .QN(n19653) );
  OA22X1 U22267 ( .IN1(n19641), .IN2(n22618), .IN3(n19640), .IN4(n21102), .Q(
        n19651) );
  OA22X1 U22268 ( .IN1(n19643), .IN2(n21081), .IN3(n19642), .IN4(n21088), .Q(
        n19650) );
  OA22X1 U22269 ( .IN1(n19645), .IN2(n21090), .IN3(n19644), .IN4(n21083), .Q(
        n19649) );
  OA22X1 U22270 ( .IN1(n19647), .IN2(n22616), .IN3(n19646), .IN4(n21099), .Q(
        n19648) );
  NAND4X0 U22271 ( .IN1(n19651), .IN2(n19650), .IN3(n19649), .IN4(n19648), 
        .QN(n19652) );
  NOR2X0 U22272 ( .IN1(n19653), .IN2(n19652), .QN(n19656) );
  NAND2X0 U22273 ( .IN1(s15_data_i[31]), .IN2(n19654), .QN(n19655) );
  NAND2X0 U22274 ( .IN1(n19656), .IN2(n19655), .QN(m4_data_o[31]) );
  NOR2X0 U22275 ( .IN1(m3s0_addr[31]), .IN2(m3s0_addr[30]), .QN(n19657) );
  INVX0 U22276 ( .INP(m3s0_addr[29]), .ZN(n28919) );
  NOR2X0 U22277 ( .IN1(m3s0_addr[28]), .IN2(n28919), .QN(n19668) );
  AND2X1 U22278 ( .IN1(n19657), .IN2(n19668), .Q(n29306) );
  INVX0 U22279 ( .INP(n23114), .ZN(n23210) );
  NAND2X0 U22280 ( .IN1(n21133), .IN2(n23113), .QN(n19999) );
  NOR2X0 U22281 ( .IN1(n23210), .IN2(n19999), .QN(n29011) );
  NAND2X0 U22282 ( .IN1(n29306), .IN2(n29011), .QN(n27500) );
  INVX0 U22283 ( .INP(m3s0_addr[28]), .ZN(n28908) );
  NOR2X0 U22284 ( .IN1(m3s0_addr[29]), .IN2(n28908), .QN(n19662) );
  INVX0 U22285 ( .INP(m3s0_addr[30]), .ZN(n28940) );
  NOR2X0 U22286 ( .IN1(m3s0_addr[31]), .IN2(n28940), .QN(n19663) );
  AND2X1 U22287 ( .IN1(n19662), .IN2(n19663), .Q(n29303) );
  INVX0 U22288 ( .INP(n23227), .ZN(n23134) );
  NAND2X0 U22289 ( .IN1(n21143), .IN2(n23132), .QN(n20015) );
  NOR2X0 U22290 ( .IN1(n23134), .IN2(n20015), .QN(n29064) );
  NAND2X0 U22291 ( .IN1(n29303), .IN2(n29064), .QN(n26589) );
  OA22X1 U22292 ( .IN1(n23214), .IN2(n27500), .IN3(n21144), .IN4(n26589), .Q(
        n19661) );
  INVX0 U22293 ( .INP(m3s0_addr[31]), .ZN(n28958) );
  NOR2X0 U22294 ( .IN1(m3s0_addr[30]), .IN2(n28958), .QN(n19669) );
  AND2X1 U22295 ( .IN1(n19662), .IN2(n19669), .Q(n29299) );
  INVX0 U22296 ( .INP(n23117), .ZN(n23249) );
  NAND2X0 U22297 ( .IN1(n21142), .IN2(n23116), .QN(n19998) );
  NOR2X0 U22298 ( .IN1(n23249), .IN2(n19998), .QN(n29127) );
  NAND2X0 U22299 ( .IN1(n29299), .IN2(n29127), .QN(n25369) );
  NOR2X0 U22300 ( .IN1(n28908), .IN2(n28919), .QN(n19666) );
  AND2X1 U22301 ( .IN1(n19666), .IN2(n19657), .Q(n29305) );
  INVX0 U22302 ( .INP(n23233), .ZN(n23166) );
  NAND2X0 U22303 ( .IN1(n21118), .IN2(n23164), .QN(n19997) );
  NOR2X0 U22304 ( .IN1(n23166), .IN2(n19997), .QN(n29028) );
  NAND2X0 U22305 ( .IN1(n29305), .IN2(n29028), .QN(n27198) );
  OA22X1 U22306 ( .IN1(n23253), .IN2(n25369), .IN3(n21120), .IN4(n27198), .Q(
        n19660) );
  NOR2X0 U22307 ( .IN1(n28958), .IN2(n28940), .QN(n19667) );
  NOR2X0 U22308 ( .IN1(m3s0_addr[28]), .IN2(m3s0_addr[29]), .QN(n19664) );
  AND2X1 U22309 ( .IN1(n19667), .IN2(n19664), .Q(n29296) );
  INVX0 U22310 ( .INP(n23224), .ZN(n23152) );
  NAND2X0 U22311 ( .IN1(n23151), .IN2(n21139), .QN(n20018) );
  NOR2X0 U22312 ( .IN1(n23152), .IN2(n20018), .QN(n29184) );
  NAND2X0 U22313 ( .IN1(n29296), .IN2(n29184), .QN(n24455) );
  AND2X1 U22314 ( .IN1(n19664), .IN2(n19657), .Q(n29309) );
  INVX0 U22315 ( .INP(n23251), .ZN(n23156) );
  NAND2X0 U22316 ( .IN1(n23154), .IN2(n21140), .QN(n20006) );
  NOR2X0 U22317 ( .IN1(n23156), .IN2(n20006), .QN(n28967) );
  NAND2X0 U22318 ( .IN1(n29309), .IN2(n28967), .QN(n28110) );
  OA22X1 U22319 ( .IN1(n21141), .IN2(n24455), .IN3(n23252), .IN4(n28110), .Q(
        n19659) );
  AND2X1 U22320 ( .IN1(n19662), .IN2(n19657), .Q(n29307) );
  NAND3X0 U22321 ( .IN1(n23236), .IN2(n23140), .IN3(n21135), .QN(n28090) );
  NAND2X0 U22322 ( .IN1(n29307), .IN2(n28986), .QN(n27802) );
  OR2X1 U22323 ( .IN1(n21138), .IN2(n27802), .Q(n19658) );
  NAND4X0 U22324 ( .IN1(n19661), .IN2(n19660), .IN3(n19659), .IN4(n19658), 
        .QN(n19675) );
  AND2X1 U22325 ( .IN1(n19663), .IN2(n19668), .Q(n29302) );
  INVX0 U22326 ( .INP(n23230), .ZN(n23138) );
  NAND2X0 U22327 ( .IN1(n21125), .IN2(n23136), .QN(n19993) );
  NOR2X0 U22328 ( .IN1(n23138), .IN2(n19993), .QN(n29073) );
  NAND2X0 U22329 ( .IN1(n29302), .IN2(n29073), .QN(n26279) );
  AND2X1 U22330 ( .IN1(n19667), .IN2(n19662), .Q(n29295) );
  INVX0 U22331 ( .INP(n23212), .ZN(n23130) );
  NAND2X0 U22332 ( .IN1(n21127), .IN2(n23129), .QN(n20004) );
  NOR2X0 U22333 ( .IN1(n23130), .IN2(n20004), .QN(n29210) );
  NAND2X0 U22334 ( .IN1(n29295), .IN2(n29210), .QN(n24152) );
  OA22X1 U22335 ( .IN1(n21126), .IN2(n26279), .IN3(n23213), .IN4(n24152), .Q(
        n19673) );
  AND2X1 U22336 ( .IN1(n19664), .IN2(n19663), .Q(n29304) );
  INVX0 U22337 ( .INP(n23120), .ZN(n23243) );
  NAND2X0 U22338 ( .IN1(n21124), .IN2(n23118), .QN(n19994) );
  NOR2X0 U22339 ( .IN1(n23243), .IN2(n19994), .QN(n29046) );
  NAND2X0 U22340 ( .IN1(n29304), .IN2(n29046), .QN(n26893) );
  AND2X1 U22341 ( .IN1(n19666), .IN2(n19663), .Q(n29301) );
  INVX0 U22342 ( .INP(n23215), .ZN(n23145) );
  NAND2X0 U22343 ( .IN1(n21119), .IN2(n23143), .QN(n20008) );
  NOR2X0 U22344 ( .IN1(n23145), .IN2(n20008), .QN(n29092) );
  NAND2X0 U22345 ( .IN1(n29301), .IN2(n29092), .QN(n25977) );
  OA22X1 U22346 ( .IN1(n23247), .IN2(n26893), .IN3(n23220), .IN4(n25977), .Q(
        n19672) );
  NAND2X0 U22347 ( .IN1(n19669), .IN2(n19664), .QN(n23091) );
  INVX0 U22348 ( .INP(n23091), .ZN(n29300) );
  NAND2X0 U22349 ( .IN1(n19665), .IN2(n23122), .QN(n19995) );
  NOR2X0 U22350 ( .IN1(n23245), .IN2(n19995), .QN(n29119) );
  NAND2X0 U22351 ( .IN1(n29300), .IN2(n29119), .QN(n25671) );
  AND2X1 U22352 ( .IN1(n19666), .IN2(n19669), .Q(n29297) );
  INVX0 U22353 ( .INP(n23221), .ZN(n23148) );
  NAND2X0 U22354 ( .IN1(n23147), .IN2(n21136), .QN(n19996) );
  NOR2X0 U22355 ( .IN1(n23148), .IN2(n19996), .QN(n29166) );
  NAND2X0 U22356 ( .IN1(n29297), .IN2(n29166), .QN(n24762) );
  OA22X1 U22357 ( .IN1(n23246), .IN2(n25671), .IN3(n21137), .IN4(n24762), .Q(
        n19671) );
  AND2X1 U22358 ( .IN1(n19667), .IN2(n19668), .Q(n29294) );
  INVX0 U22359 ( .INP(n23240), .ZN(n23126) );
  NAND2X0 U22360 ( .IN1(n23124), .IN2(n21122), .QN(n20005) );
  NOR2X0 U22361 ( .IN1(n23126), .IN2(n20005), .QN(n29225) );
  NAND2X0 U22362 ( .IN1(n29294), .IN2(n29225), .QN(n23850) );
  AND2X1 U22363 ( .IN1(n19669), .IN2(n19668), .Q(n29298) );
  INVX0 U22364 ( .INP(n23217), .ZN(n23160) );
  NAND2X0 U22365 ( .IN1(n21134), .IN2(n23158), .QN(n20011) );
  NOR2X0 U22366 ( .IN1(n23160), .IN2(n20011), .QN(n29147) );
  NAND2X0 U22367 ( .IN1(n29298), .IN2(n29147), .QN(n25065) );
  OA22X1 U22368 ( .IN1(n21123), .IN2(n23850), .IN3(n23219), .IN4(n25065), .Q(
        n19670) );
  NAND4X0 U22369 ( .IN1(n19673), .IN2(n19672), .IN3(n19671), .IN4(n19670), 
        .QN(n19674) );
  NOR2X0 U22370 ( .IN1(n19675), .IN2(n19674), .QN(n19677) );
  NAND2X0 U22371 ( .IN1(n23314), .IN2(n23261), .QN(n19676) );
  NAND2X0 U22372 ( .IN1(n19677), .IN2(n19676), .QN(m3_ack_o) );
  INVX0 U22373 ( .INP(n29294), .ZN(n23069) );
  INVX0 U22374 ( .INP(n29307), .ZN(n23085) );
  OA22X1 U22375 ( .IN1(n21154), .IN2(n23069), .IN3(n21161), .IN4(n23085), .Q(
        n19681) );
  INVX0 U22376 ( .INP(n29298), .ZN(n23083) );
  INVX0 U22377 ( .INP(n29295), .ZN(n19979) );
  OA22X1 U22378 ( .IN1(n22207), .IN2(n23083), .IN3(n21823), .IN4(n19979), .Q(
        n19680) );
  INVX0 U22379 ( .INP(m0s5_data_i[0]), .ZN(n21160) );
  INVX0 U22380 ( .INP(n29303), .ZN(n22982) );
  INVX0 U22381 ( .INP(n29304), .ZN(n23063) );
  OA22X1 U22382 ( .IN1(n21160), .IN2(n22982), .IN3(n22203), .IN4(n23063), .Q(
        n19679) );
  NAND2X0 U22383 ( .IN1(m0s2_data_i[0]), .IN2(n29306), .QN(n19678) );
  NAND4X0 U22384 ( .IN1(n19681), .IN2(n19680), .IN3(n19679), .IN4(n19678), 
        .QN(n19687) );
  INVX0 U22385 ( .INP(n29305), .ZN(n23089) );
  INVX0 U22386 ( .INP(n29301), .ZN(n23093) );
  OA22X1 U22387 ( .IN1(n22206), .IN2(n23089), .IN3(n21162), .IN4(n23093), .Q(
        n19685) );
  OA22X1 U22388 ( .IN1(n21163), .IN2(n23091), .IN3(n21159), .IN4(n23021), .Q(
        n19684) );
  INVX0 U22389 ( .INP(n29297), .ZN(n23067) );
  INVX0 U22390 ( .INP(n29309), .ZN(n23065) );
  OA22X1 U22391 ( .IN1(n22208), .IN2(n23067), .IN3(n22204), .IN4(n23065), .Q(
        n19683) );
  INVX0 U22392 ( .INP(n29302), .ZN(n23003) );
  OA22X1 U22393 ( .IN1(n20251), .IN2(n23087), .IN3(n21153), .IN4(n23003), .Q(
        n19682) );
  NAND4X0 U22394 ( .IN1(n19685), .IN2(n19684), .IN3(n19683), .IN4(n19682), 
        .QN(n19686) );
  NOR2X0 U22395 ( .IN1(n19687), .IN2(n19686), .QN(n19689) );
  INVX0 U22396 ( .INP(n19808), .ZN(n29293) );
  NAND2X0 U22397 ( .IN1(n29293), .IN2(n22218), .QN(n19688) );
  NAND2X0 U22398 ( .IN1(n19689), .IN2(n19688), .QN(m3_data_o[0]) );
  OA22X1 U22399 ( .IN1(n21182), .IN2(n23085), .IN3(n21186), .IN4(n23083), .Q(
        n19693) );
  OA22X1 U22400 ( .IN1(n21184), .IN2(n19979), .IN3(n21173), .IN4(n23063), .Q(
        n19692) );
  OA22X1 U22401 ( .IN1(n21176), .IN2(n23089), .IN3(n22224), .IN4(n23069), .Q(
        n19691) );
  NAND2X0 U22402 ( .IN1(m0s0_data_i[1]), .IN2(n29309), .QN(n19690) );
  NAND4X0 U22403 ( .IN1(n19693), .IN2(n19692), .IN3(n19691), .IN4(n19690), 
        .QN(n19699) );
  OA22X1 U22404 ( .IN1(n22226), .IN2(n23093), .IN3(n21174), .IN4(n23091), .Q(
        n19697) );
  OA22X1 U22405 ( .IN1(n21175), .IN2(n23003), .IN3(n21183), .IN4(n23021), .Q(
        n19696) );
  INVX0 U22406 ( .INP(m0s11_data_i[1]), .ZN(n20689) );
  OA22X1 U22407 ( .IN1(n21185), .IN2(n23087), .IN3(n20689), .IN4(n23067), .Q(
        n19695) );
  INVX0 U22408 ( .INP(n29306), .ZN(n23059) );
  OA22X1 U22409 ( .IN1(n21177), .IN2(n22982), .IN3(n22225), .IN4(n23059), .Q(
        n19694) );
  NAND4X0 U22410 ( .IN1(n19697), .IN2(n19696), .IN3(n19695), .IN4(n19694), 
        .QN(n19698) );
  NOR2X0 U22411 ( .IN1(n19699), .IN2(n19698), .QN(n19701) );
  NAND2X0 U22412 ( .IN1(n29293), .IN2(n22235), .QN(n19700) );
  NAND2X0 U22413 ( .IN1(n19701), .IN2(n19700), .QN(m3_data_o[1]) );
  OA22X1 U22414 ( .IN1(n21205), .IN2(n23065), .IN3(n21208), .IN4(n23003), .Q(
        n19705) );
  INVX0 U22415 ( .INP(n29299), .ZN(n23021) );
  OA22X1 U22416 ( .IN1(n21210), .IN2(n23021), .IN3(n21207), .IN4(n23059), .Q(
        n19704) );
  OA22X1 U22417 ( .IN1(n21211), .IN2(n22982), .IN3(n21199), .IN4(n23085), .Q(
        n19703) );
  NAND2X0 U22418 ( .IN1(m0s14_data_i[2]), .IN2(n29294), .QN(n19702) );
  NAND4X0 U22419 ( .IN1(n19705), .IN2(n19704), .IN3(n19703), .IN4(n19702), 
        .QN(n19711) );
  OA22X1 U22420 ( .IN1(n21196), .IN2(n23091), .IN3(n21206), .IN4(n23083), .Q(
        n19709) );
  INVX0 U22421 ( .INP(m0s3_data_i[2]), .ZN(n21200) );
  OA22X1 U22422 ( .IN1(n21200), .IN2(n23089), .IN3(n21197), .IN4(n23063), .Q(
        n19708) );
  OA22X1 U22423 ( .IN1(n21212), .IN2(n19979), .IN3(n20702), .IN4(n23067), .Q(
        n19707) );
  OA22X1 U22424 ( .IN1(n21198), .IN2(n23087), .IN3(n21209), .IN4(n23093), .Q(
        n19706) );
  NAND4X0 U22425 ( .IN1(n19709), .IN2(n19708), .IN3(n19707), .IN4(n19706), 
        .QN(n19710) );
  NOR2X0 U22426 ( .IN1(n19711), .IN2(n19710), .QN(n19713) );
  NAND2X0 U22427 ( .IN1(n29293), .IN2(n22247), .QN(n19712) );
  NAND2X0 U22428 ( .IN1(n19713), .IN2(n19712), .QN(m3_data_o[2]) );
  INVX0 U22429 ( .INP(m0s5_data_i[3]), .ZN(n22637) );
  OA22X1 U22430 ( .IN1(n21222), .IN2(n23093), .IN3(n22637), .IN4(n22982), .Q(
        n19717) );
  OA22X1 U22431 ( .IN1(n22635), .IN2(n23087), .IN3(n21235), .IN4(n23065), .Q(
        n19716) );
  OA22X1 U22432 ( .IN1(n21226), .IN2(n23085), .IN3(n21224), .IN4(n23003), .Q(
        n19715) );
  NAND2X0 U22433 ( .IN1(m0s3_data_i[3]), .IN2(n29305), .QN(n19714) );
  NAND4X0 U22434 ( .IN1(n19717), .IN2(n19716), .IN3(n19715), .IN4(n19714), 
        .QN(n19723) );
  OA22X1 U22435 ( .IN1(n21234), .IN2(n23067), .IN3(n21231), .IN4(n23069), .Q(
        n19721) );
  OA22X1 U22436 ( .IN1(n22634), .IN2(n23063), .IN3(n21232), .IN4(n23083), .Q(
        n19720) );
  OA22X1 U22437 ( .IN1(n22636), .IN2(n19979), .IN3(n21223), .IN4(n23021), .Q(
        n19719) );
  OA22X1 U22438 ( .IN1(n21225), .IN2(n23059), .IN3(n21233), .IN4(n23091), .Q(
        n19718) );
  NAND4X0 U22439 ( .IN1(n19721), .IN2(n19720), .IN3(n19719), .IN4(n19718), 
        .QN(n19722) );
  NOR2X0 U22440 ( .IN1(n19723), .IN2(n19722), .QN(n19725) );
  NAND2X0 U22441 ( .IN1(n29293), .IN2(n22646), .QN(n19724) );
  NAND2X0 U22442 ( .IN1(n19725), .IN2(n19724), .QN(m3_data_o[3]) );
  OA22X1 U22443 ( .IN1(n21246), .IN2(n23085), .IN3(n22653), .IN4(n19979), .Q(
        n19729) );
  OA22X1 U22444 ( .IN1(n22654), .IN2(n23087), .IN3(n22651), .IN4(n23063), .Q(
        n19728) );
  OA22X1 U22445 ( .IN1(n22652), .IN2(n23059), .IN3(n21245), .IN4(n23083), .Q(
        n19727) );
  NAND2X0 U22446 ( .IN1(m0s5_data_i[4]), .IN2(n29303), .QN(n19726) );
  NAND4X0 U22447 ( .IN1(n19729), .IN2(n19728), .IN3(n19727), .IN4(n19726), 
        .QN(n19735) );
  OA22X1 U22448 ( .IN1(n20727), .IN2(n23089), .IN3(n21257), .IN4(n23093), .Q(
        n19733) );
  OA22X1 U22449 ( .IN1(n21255), .IN2(n23067), .IN3(n21244), .IN4(n23069), .Q(
        n19732) );
  OA22X1 U22450 ( .IN1(n21248), .IN2(n23003), .IN3(n21247), .IN4(n23021), .Q(
        n19731) );
  INVX0 U22451 ( .INP(m0s8_data_i[4]), .ZN(n21256) );
  OA22X1 U22452 ( .IN1(n21256), .IN2(n23091), .IN3(n21254), .IN4(n23065), .Q(
        n19730) );
  NAND4X0 U22453 ( .IN1(n19733), .IN2(n19732), .IN3(n19731), .IN4(n19730), 
        .QN(n19734) );
  NOR2X0 U22454 ( .IN1(n19735), .IN2(n19734), .QN(n19737) );
  NAND2X0 U22455 ( .IN1(n29293), .IN2(n22663), .QN(n19736) );
  NAND2X0 U22456 ( .IN1(n19737), .IN2(n19736), .QN(m3_data_o[4]) );
  OA22X1 U22457 ( .IN1(n21279), .IN2(n23003), .IN3(n21267), .IN4(n23021), .Q(
        n19741) );
  OA22X1 U22458 ( .IN1(n21269), .IN2(n23063), .IN3(n22671), .IN4(n19979), .Q(
        n19740) );
  INVX0 U22459 ( .INP(m0s10_data_i[5]), .ZN(n21278) );
  OA22X1 U22460 ( .IN1(n21278), .IN2(n23083), .IN3(n22668), .IN4(n23089), .Q(
        n19739) );
  NAND2X0 U22461 ( .IN1(m0s11_data_i[5]), .IN2(n29297), .QN(n19738) );
  NAND4X0 U22462 ( .IN1(n19741), .IN2(n19740), .IN3(n19739), .IN4(n19738), 
        .QN(n19747) );
  INVX0 U22463 ( .INP(n29296), .ZN(n23087) );
  OA22X1 U22464 ( .IN1(n21277), .IN2(n23065), .IN3(n21266), .IN4(n23087), .Q(
        n19745) );
  OA22X1 U22465 ( .IN1(n20736), .IN2(n22982), .IN3(n21276), .IN4(n23091), .Q(
        n19744) );
  OA22X1 U22466 ( .IN1(n22669), .IN2(n23059), .IN3(n22670), .IN4(n23093), .Q(
        n19743) );
  OA22X1 U22467 ( .IN1(n21275), .IN2(n23069), .IN3(n21274), .IN4(n23085), .Q(
        n19742) );
  NAND4X0 U22468 ( .IN1(n19745), .IN2(n19744), .IN3(n19743), .IN4(n19742), 
        .QN(n19746) );
  NOR2X0 U22469 ( .IN1(n19747), .IN2(n19746), .QN(n19749) );
  NAND2X0 U22470 ( .IN1(n29293), .IN2(n22680), .QN(n19748) );
  NAND2X0 U22471 ( .IN1(n19749), .IN2(n19748), .QN(m3_data_o[5]) );
  OA22X1 U22472 ( .IN1(n21291), .IN2(n23087), .IN3(n21301), .IN4(n23085), .Q(
        n19753) );
  OA22X1 U22473 ( .IN1(n22686), .IN2(n23083), .IN3(n22685), .IN4(n23089), .Q(
        n19752) );
  OA22X1 U22474 ( .IN1(n22688), .IN2(n23091), .IN3(n20753), .IN4(n23067), .Q(
        n19751) );
  NAND2X0 U22475 ( .IN1(m0s0_data_i[6]), .IN2(n29309), .QN(n19750) );
  NAND4X0 U22476 ( .IN1(n19753), .IN2(n19752), .IN3(n19751), .IN4(n19750), 
        .QN(n19759) );
  OA22X1 U22477 ( .IN1(n21297), .IN2(n23059), .IN3(n21288), .IN4(n23069), .Q(
        n19757) );
  OA22X1 U22478 ( .IN1(n21298), .IN2(n23003), .IN3(n21290), .IN4(n23063), .Q(
        n19756) );
  OA22X1 U22479 ( .IN1(n21292), .IN2(n22982), .IN3(n21300), .IN4(n23021), .Q(
        n19755) );
  INVX0 U22480 ( .INP(m0s7_data_i[6]), .ZN(n21289) );
  OA22X1 U22481 ( .IN1(n21289), .IN2(n23093), .IN3(n22687), .IN4(n19979), .Q(
        n19754) );
  NAND4X0 U22482 ( .IN1(n19757), .IN2(n19756), .IN3(n19755), .IN4(n19754), 
        .QN(n19758) );
  NOR2X0 U22483 ( .IN1(n19759), .IN2(n19758), .QN(n19761) );
  NAND2X0 U22484 ( .IN1(n29293), .IN2(n22697), .QN(n19760) );
  NAND2X0 U22485 ( .IN1(n19761), .IN2(n19760), .QN(m3_data_o[6]) );
  OA22X1 U22486 ( .IN1(n22705), .IN2(n23063), .IN3(n21319), .IN4(n23091), .Q(
        n19765) );
  OA22X1 U22487 ( .IN1(n21311), .IN2(n23085), .IN3(n21310), .IN4(n23067), .Q(
        n19764) );
  OA22X1 U22488 ( .IN1(n21312), .IN2(n22982), .IN3(n22704), .IN4(n23087), .Q(
        n19763) );
  NAND2X0 U22489 ( .IN1(m0s9_data_i[7]), .IN2(n29299), .QN(n19762) );
  NAND4X0 U22490 ( .IN1(n19765), .IN2(n19764), .IN3(n19763), .IN4(n19762), 
        .QN(n19771) );
  OA22X1 U22491 ( .IN1(n20766), .IN2(n23093), .IN3(n22702), .IN4(n23059), .Q(
        n19769) );
  INVX0 U22492 ( .INP(m0s0_data_i[7]), .ZN(n22703) );
  OA22X1 U22493 ( .IN1(n22703), .IN2(n23065), .IN3(n21323), .IN4(n23069), .Q(
        n19768) );
  OA22X1 U22494 ( .IN1(n21314), .IN2(n23083), .IN3(n21320), .IN4(n23089), .Q(
        n19767) );
  OA22X1 U22495 ( .IN1(n21321), .IN2(n23003), .IN3(n21313), .IN4(n19979), .Q(
        n19766) );
  NAND4X0 U22496 ( .IN1(n19769), .IN2(n19768), .IN3(n19767), .IN4(n19766), 
        .QN(n19770) );
  NOR2X0 U22497 ( .IN1(n19771), .IN2(n19770), .QN(n19773) );
  NAND2X0 U22498 ( .IN1(n29293), .IN2(n22714), .QN(n19772) );
  NAND2X0 U22499 ( .IN1(n19773), .IN2(n19772), .QN(m3_data_o[7]) );
  INVX0 U22500 ( .INP(m0s11_data_i[8]), .ZN(n21333) );
  OA22X1 U22501 ( .IN1(n21333), .IN2(n23067), .IN3(n21345), .IN4(n23003), .Q(
        n19777) );
  OA22X1 U22502 ( .IN1(n21346), .IN2(n19979), .IN3(n21343), .IN4(n23069), .Q(
        n19776) );
  OA22X1 U22503 ( .IN1(n21342), .IN2(n22982), .IN3(n22722), .IN4(n23085), .Q(
        n19775) );
  NAND2X0 U22504 ( .IN1(m0s8_data_i[8]), .IN2(n29300), .QN(n19774) );
  NAND4X0 U22505 ( .IN1(n19777), .IN2(n19776), .IN3(n19775), .IN4(n19774), 
        .QN(n19783) );
  OA22X1 U22506 ( .IN1(n21344), .IN2(n23087), .IN3(n22720), .IN4(n23093), .Q(
        n19781) );
  OA22X1 U22507 ( .IN1(n21335), .IN2(n23063), .IN3(n21337), .IN4(n23083), .Q(
        n19780) );
  OA22X1 U22508 ( .IN1(n21334), .IN2(n23089), .IN3(n21332), .IN4(n23021), .Q(
        n19779) );
  OA22X1 U22509 ( .IN1(n22721), .IN2(n23065), .IN3(n21336), .IN4(n23059), .Q(
        n19778) );
  NAND4X0 U22510 ( .IN1(n19781), .IN2(n19780), .IN3(n19779), .IN4(n19778), 
        .QN(n19782) );
  NOR2X0 U22511 ( .IN1(n19783), .IN2(n19782), .QN(n19785) );
  NAND2X0 U22512 ( .IN1(n29293), .IN2(n22731), .QN(n19784) );
  NAND2X0 U22513 ( .IN1(n19785), .IN2(n19784), .QN(m3_data_o[8]) );
  OA22X1 U22514 ( .IN1(n22754), .IN2(n23087), .IN3(n22751), .IN4(n23083), .Q(
        n19789) );
  OA22X1 U22515 ( .IN1(n22750), .IN2(n23093), .IN3(n22753), .IN4(n23063), .Q(
        n19788) );
  OA22X1 U22516 ( .IN1(n21385), .IN2(n23021), .IN3(n21376), .IN4(n22982), .Q(
        n19787) );
  NAND2X0 U22517 ( .IN1(m0s13_data_i[10]), .IN2(n29295), .QN(n19786) );
  NAND4X0 U22518 ( .IN1(n19789), .IN2(n19788), .IN3(n19787), .IN4(n19786), 
        .QN(n19795) );
  INVX0 U22519 ( .INP(m0s2_data_i[10]), .ZN(n22749) );
  OA22X1 U22520 ( .IN1(n21382), .IN2(n23067), .IN3(n22749), .IN4(n23059), .Q(
        n19793) );
  OA22X1 U22521 ( .IN1(n22329), .IN2(n23069), .IN3(n21377), .IN4(n23091), .Q(
        n19792) );
  OA22X1 U22522 ( .IN1(n21374), .IN2(n23003), .IN3(n21384), .IN4(n23085), .Q(
        n19791) );
  OA22X1 U22523 ( .IN1(n22752), .IN2(n23089), .IN3(n21375), .IN4(n23065), .Q(
        n19790) );
  NAND4X0 U22524 ( .IN1(n19793), .IN2(n19792), .IN3(n19791), .IN4(n19790), 
        .QN(n19794) );
  NOR2X0 U22525 ( .IN1(n19795), .IN2(n19794), .QN(n19797) );
  NAND2X0 U22526 ( .IN1(n29293), .IN2(n22763), .QN(n19796) );
  NAND2X0 U22527 ( .IN1(n19797), .IN2(n19796), .QN(m3_data_o[10]) );
  INVX0 U22528 ( .INP(m0s13_data_i[16]), .ZN(n22010) );
  OA22X1 U22529 ( .IN1(n23069), .IN2(n21492), .IN3(n19979), .IN4(n22010), .Q(
        n19801) );
  OA22X1 U22530 ( .IN1(n23089), .IN2(n21491), .IN3(n23059), .IN4(n21490), .Q(
        n19800) );
  OA22X1 U22531 ( .IN1(n23085), .IN2(n21503), .IN3(n22982), .IN4(n22009), .Q(
        n19799) );
  NAND2X0 U22532 ( .IN1(n29309), .IN2(m0s0_data_i[16]), .QN(n19798) );
  NAND4X0 U22533 ( .IN1(n19801), .IN2(n19800), .IN3(n19799), .IN4(n19798), 
        .QN(n19807) );
  OA22X1 U22534 ( .IN1(n23021), .IN2(n21493), .IN3(n23087), .IN4(n22012), .Q(
        n19805) );
  OA22X1 U22535 ( .IN1(n23093), .IN2(n21500), .IN3(n23003), .IN4(n21502), .Q(
        n19804) );
  OA22X1 U22536 ( .IN1(n23083), .IN2(n21501), .IN3(n23063), .IN4(n21494), .Q(
        n19803) );
  OA22X1 U22537 ( .IN1(n23091), .IN2(n21499), .IN3(n23067), .IN4(n22011), .Q(
        n19802) );
  NAND4X0 U22538 ( .IN1(n19805), .IN2(n19804), .IN3(n19803), .IN4(n19802), 
        .QN(n19806) );
  NOR2X0 U22539 ( .IN1(n19807), .IN2(n19806), .QN(n19810) );
  NOR2X0 U22540 ( .IN1(n23501), .IN2(n19808), .QN(n19990) );
  NAND2X0 U22541 ( .IN1(s15_data_i[16]), .IN2(n19990), .QN(n19809) );
  NAND2X0 U22542 ( .IN1(n19810), .IN2(n19809), .QN(m3_data_o[16]) );
  OA22X1 U22543 ( .IN1(n23091), .IN2(n22397), .IN3(n23067), .IN4(n22832), .Q(
        n19814) );
  OA22X1 U22544 ( .IN1(n23083), .IN2(n22834), .IN3(n23063), .IN4(n22833), .Q(
        n19813) );
  OA22X1 U22545 ( .IN1(n23065), .IN2(n21520), .IN3(n22982), .IN4(n21513), .Q(
        n19812) );
  NAND2X0 U22546 ( .IN1(n29295), .IN2(m0s13_data_i[17]), .QN(n19811) );
  NAND4X0 U22547 ( .IN1(n19814), .IN2(n19813), .IN3(n19812), .IN4(n19811), 
        .QN(n19820) );
  OA22X1 U22548 ( .IN1(n23089), .IN2(n22830), .IN3(n23069), .IN4(n21519), .Q(
        n19818) );
  OA22X1 U22549 ( .IN1(n23021), .IN2(n22835), .IN3(n23059), .IN4(n21512), .Q(
        n19817) );
  OA22X1 U22550 ( .IN1(n23003), .IN2(n21521), .IN3(n23085), .IN4(n21518), .Q(
        n19816) );
  INVX0 U22551 ( .INP(m0s12_data_i[17]), .ZN(n22837) );
  OA22X1 U22552 ( .IN1(n23093), .IN2(n22831), .IN3(n23087), .IN4(n22837), .Q(
        n19815) );
  NAND4X0 U22553 ( .IN1(n19818), .IN2(n19817), .IN3(n19816), .IN4(n19815), 
        .QN(n19819) );
  NOR2X0 U22554 ( .IN1(n19820), .IN2(n19819), .QN(n19822) );
  NAND2X0 U22555 ( .IN1(s15_data_i[17]), .IN2(n19990), .QN(n19821) );
  NAND2X0 U22556 ( .IN1(n19822), .IN2(n19821), .QN(m3_data_o[17]) );
  OA22X1 U22557 ( .IN1(n23067), .IN2(n21537), .IN3(n23085), .IN4(n22037), .Q(
        n19826) );
  OA22X1 U22558 ( .IN1(n19979), .IN2(n21539), .IN3(n23063), .IN4(n21536), .Q(
        n19825) );
  OA22X1 U22559 ( .IN1(n23091), .IN2(n21531), .IN3(n23065), .IN4(n22415), .Q(
        n19824) );
  NAND2X0 U22560 ( .IN1(n29302), .IN2(m0s6_data_i[18]), .QN(n19823) );
  NAND4X0 U22561 ( .IN1(n19826), .IN2(n19825), .IN3(n19824), .IN4(n19823), 
        .QN(n19832) );
  OA22X1 U22562 ( .IN1(n23021), .IN2(n21530), .IN3(n23087), .IN4(n22410), .Q(
        n19830) );
  OA22X1 U22563 ( .IN1(n23089), .IN2(n22413), .IN3(n22982), .IN4(n22414), .Q(
        n19829) );
  OA22X1 U22564 ( .IN1(n23059), .IN2(n21538), .IN3(n23083), .IN4(n21540), .Q(
        n19828) );
  OA22X1 U22565 ( .IN1(n23093), .IN2(n22411), .IN3(n23069), .IN4(n20901), .Q(
        n19827) );
  NAND4X0 U22566 ( .IN1(n19830), .IN2(n19829), .IN3(n19828), .IN4(n19827), 
        .QN(n19831) );
  NOR2X0 U22567 ( .IN1(n19832), .IN2(n19831), .QN(n19834) );
  NAND2X0 U22568 ( .IN1(s15_data_i[18]), .IN2(n19990), .QN(n19833) );
  NAND2X0 U22569 ( .IN1(n19834), .IN2(n19833), .QN(m3_data_o[18]) );
  OA22X1 U22570 ( .IN1(n23089), .IN2(n22431), .IN3(n22982), .IN4(n22050), .Q(
        n19838) );
  OA22X1 U22571 ( .IN1(n23021), .IN2(n22429), .IN3(n23091), .IN4(n21550), .Q(
        n19837) );
  OA22X1 U22572 ( .IN1(n23059), .IN2(n21558), .IN3(n23069), .IN4(n22428), .Q(
        n19836) );
  NAND2X0 U22573 ( .IN1(n29304), .IN2(m0s4_data_i[19]), .QN(n19835) );
  NAND4X0 U22574 ( .IN1(n19838), .IN2(n19837), .IN3(n19836), .IN4(n19835), 
        .QN(n19844) );
  OA22X1 U22575 ( .IN1(n23093), .IN2(n22435), .IN3(n23087), .IN4(n22434), .Q(
        n19842) );
  OA22X1 U22576 ( .IN1(n23067), .IN2(n21549), .IN3(n23083), .IN4(n22432), .Q(
        n19841) );
  INVX0 U22577 ( .INP(m0s13_data_i[19]), .ZN(n22430) );
  OA22X1 U22578 ( .IN1(n23085), .IN2(n21557), .IN3(n19979), .IN4(n22430), .Q(
        n19840) );
  OA22X1 U22579 ( .IN1(n23003), .IN2(n21551), .IN3(n23065), .IN4(n22433), .Q(
        n19839) );
  NAND4X0 U22580 ( .IN1(n19842), .IN2(n19841), .IN3(n19840), .IN4(n19839), 
        .QN(n19843) );
  NOR2X0 U22581 ( .IN1(n19844), .IN2(n19843), .QN(n19846) );
  NAND2X0 U22582 ( .IN1(s15_data_i[19]), .IN2(n19990), .QN(n19845) );
  NAND2X0 U22583 ( .IN1(n19846), .IN2(n19845), .QN(m3_data_o[19]) );
  INVX0 U22584 ( .INP(m0s14_data_i[20]), .ZN(n22453) );
  OA22X1 U22585 ( .IN1(n23091), .IN2(n21573), .IN3(n23069), .IN4(n22453), .Q(
        n19850) );
  OA22X1 U22586 ( .IN1(n23021), .IN2(n22447), .IN3(n23083), .IN4(n21574), .Q(
        n19849) );
  OA22X1 U22587 ( .IN1(n23089), .IN2(n21568), .IN3(n23003), .IN4(n22454), .Q(
        n19848) );
  NAND2X0 U22588 ( .IN1(n29301), .IN2(m0s7_data_i[20]), .QN(n19847) );
  NAND4X0 U22589 ( .IN1(n19850), .IN2(n19849), .IN3(n19848), .IN4(n19847), 
        .QN(n19856) );
  OA22X1 U22590 ( .IN1(n23059), .IN2(n22452), .IN3(n19979), .IN4(n21567), .Q(
        n19854) );
  OA22X1 U22591 ( .IN1(n23067), .IN2(n22450), .IN3(n22982), .IN4(n22448), .Q(
        n19853) );
  OA22X1 U22592 ( .IN1(n23085), .IN2(n21575), .IN3(n23063), .IN4(n21577), .Q(
        n19852) );
  OA22X1 U22593 ( .IN1(n23087), .IN2(n22449), .IN3(n23065), .IN4(n22451), .Q(
        n19851) );
  NAND4X0 U22594 ( .IN1(n19854), .IN2(n19853), .IN3(n19852), .IN4(n19851), 
        .QN(n19855) );
  NOR2X0 U22595 ( .IN1(n19856), .IN2(n19855), .QN(n19858) );
  NAND2X0 U22596 ( .IN1(s15_data_i[20]), .IN2(n19990), .QN(n19857) );
  NAND2X0 U22597 ( .IN1(n19858), .IN2(n19857), .QN(m3_data_o[20]) );
  OA22X1 U22598 ( .IN1(n23091), .IN2(n21592), .IN3(n23085), .IN4(n22466), .Q(
        n19862) );
  OA22X1 U22599 ( .IN1(n23083), .IN2(n22849), .IN3(n22982), .IN4(n22851), .Q(
        n19861) );
  OA22X1 U22600 ( .IN1(n23093), .IN2(n22857), .IN3(n23067), .IN4(n20942), .Q(
        n19860) );
  NAND2X0 U22601 ( .IN1(n29295), .IN2(m0s13_data_i[21]), .QN(n19859) );
  NAND4X0 U22602 ( .IN1(n19862), .IN2(n19861), .IN3(n19860), .IN4(n19859), 
        .QN(n19868) );
  OA22X1 U22603 ( .IN1(n23089), .IN2(n21593), .IN3(n23065), .IN4(n22853), .Q(
        n19866) );
  OA22X1 U22604 ( .IN1(n23021), .IN2(n21594), .IN3(n23059), .IN4(n22856), .Q(
        n19865) );
  INVX0 U22605 ( .INP(m0s4_data_i[21]), .ZN(n22850) );
  OA22X1 U22606 ( .IN1(n23003), .IN2(n22855), .IN3(n23063), .IN4(n22850), .Q(
        n19864) );
  OA22X1 U22607 ( .IN1(n23087), .IN2(n22852), .IN3(n23069), .IN4(n21586), .Q(
        n19863) );
  NAND4X0 U22608 ( .IN1(n19866), .IN2(n19865), .IN3(n19864), .IN4(n19863), 
        .QN(n19867) );
  NOR2X0 U22609 ( .IN1(n19868), .IN2(n19867), .QN(n19870) );
  NAND2X0 U22610 ( .IN1(s15_data_i[21]), .IN2(n19990), .QN(n19869) );
  NAND2X0 U22611 ( .IN1(n19870), .IN2(n19869), .QN(m3_data_o[21]) );
  OA22X1 U22612 ( .IN1(n23093), .IN2(n22874), .IN3(n23059), .IN4(n22870), .Q(
        n19874) );
  OA22X1 U22613 ( .IN1(n23085), .IN2(n21612), .IN3(n19979), .IN4(n21611), .Q(
        n19873) );
  INVX0 U22614 ( .INP(m0s14_data_i[22]), .ZN(n21603) );
  OA22X1 U22615 ( .IN1(n23091), .IN2(n22873), .IN3(n23069), .IN4(n21603), .Q(
        n19872) );
  NAND2X0 U22616 ( .IN1(n29298), .IN2(m0s10_data_i[22]), .QN(n19871) );
  NAND4X0 U22617 ( .IN1(n19874), .IN2(n19873), .IN3(n19872), .IN4(n19871), 
        .QN(n19880) );
  OA22X1 U22618 ( .IN1(n23087), .IN2(n22875), .IN3(n23065), .IN4(n21604), .Q(
        n19878) );
  OA22X1 U22619 ( .IN1(n23003), .IN2(n22872), .IN3(n23067), .IN4(n20951), .Q(
        n19877) );
  OA22X1 U22620 ( .IN1(n23063), .IN2(n22876), .IN3(n22982), .IN4(n21609), .Q(
        n19876) );
  OA22X1 U22621 ( .IN1(n23021), .IN2(n21610), .IN3(n23089), .IN4(n22871), .Q(
        n19875) );
  NAND4X0 U22622 ( .IN1(n19878), .IN2(n19877), .IN3(n19876), .IN4(n19875), 
        .QN(n19879) );
  NOR2X0 U22623 ( .IN1(n19880), .IN2(n19879), .QN(n19882) );
  NAND2X0 U22624 ( .IN1(s15_data_i[22]), .IN2(n19990), .QN(n19881) );
  NAND2X0 U22625 ( .IN1(n19882), .IN2(n19881), .QN(m3_data_o[22]) );
  OA22X1 U22626 ( .IN1(n23021), .IN2(n21633), .IN3(n23083), .IN4(n22494), .Q(
        n19886) );
  INVX0 U22627 ( .INP(m0s0_data_i[23]), .ZN(n21634) );
  OA22X1 U22628 ( .IN1(n23065), .IN2(n21634), .IN3(n23069), .IN4(n21621), .Q(
        n19885) );
  OA22X1 U22629 ( .IN1(n23003), .IN2(n21625), .IN3(n23087), .IN4(n21622), .Q(
        n19884) );
  NAND2X0 U22630 ( .IN1(n29305), .IN2(m0s3_data_i[23]), .QN(n19883) );
  NAND4X0 U22631 ( .IN1(n19886), .IN2(n19885), .IN3(n19884), .IN4(n19883), 
        .QN(n19892) );
  OA22X1 U22632 ( .IN1(n23091), .IN2(n22492), .IN3(n23063), .IN4(n20968), .Q(
        n19890) );
  OA22X1 U22633 ( .IN1(n23059), .IN2(n21623), .IN3(n19979), .IN4(n21632), .Q(
        n19889) );
  OA22X1 U22634 ( .IN1(n23085), .IN2(n22491), .IN3(n22982), .IN4(n21624), .Q(
        n19888) );
  OA22X1 U22635 ( .IN1(n23093), .IN2(n22495), .IN3(n23067), .IN4(n21630), .Q(
        n19887) );
  NAND4X0 U22636 ( .IN1(n19890), .IN2(n19889), .IN3(n19888), .IN4(n19887), 
        .QN(n19891) );
  NOR2X0 U22637 ( .IN1(n19892), .IN2(n19891), .QN(n19894) );
  NAND2X0 U22638 ( .IN1(s15_data_i[23]), .IN2(n19990), .QN(n19893) );
  NAND2X0 U22639 ( .IN1(n19894), .IN2(n19893), .QN(m3_data_o[23]) );
  OA22X1 U22640 ( .IN1(n23003), .IN2(n22889), .IN3(n19979), .IN4(n22888), .Q(
        n19898) );
  OA22X1 U22641 ( .IN1(n23093), .IN2(n22891), .IN3(n23065), .IN4(n21649), .Q(
        n19897) );
  OA22X1 U22642 ( .IN1(n23091), .IN2(n21653), .IN3(n23069), .IN4(n22893), .Q(
        n19896) );
  NAND2X0 U22643 ( .IN1(n29306), .IN2(m0s2_data_i[24]), .QN(n19895) );
  NAND4X0 U22644 ( .IN1(n19898), .IN2(n19897), .IN3(n19896), .IN4(n19895), 
        .QN(n19904) );
  OA22X1 U22645 ( .IN1(n23089), .IN2(n21643), .IN3(n23087), .IN4(n21652), .Q(
        n19902) );
  INVX0 U22646 ( .INP(m0s10_data_i[24]), .ZN(n22892) );
  OA22X1 U22647 ( .IN1(n23083), .IN2(n22892), .IN3(n22982), .IN4(n22895), .Q(
        n19901) );
  OA22X1 U22648 ( .IN1(n23085), .IN2(n22896), .IN3(n23063), .IN4(n21644), .Q(
        n19900) );
  OA22X1 U22649 ( .IN1(n23021), .IN2(n21650), .IN3(n23067), .IN4(n21651), .Q(
        n19899) );
  NAND4X0 U22650 ( .IN1(n19902), .IN2(n19901), .IN3(n19900), .IN4(n19899), 
        .QN(n19903) );
  NOR2X0 U22651 ( .IN1(n19904), .IN2(n19903), .QN(n19906) );
  NAND2X0 U22652 ( .IN1(s15_data_i[24]), .IN2(n19990), .QN(n19905) );
  NAND2X0 U22653 ( .IN1(n19906), .IN2(n19905), .QN(m3_data_o[24]) );
  OA22X1 U22654 ( .IN1(n23093), .IN2(n21672), .IN3(n23067), .IN4(n21670), .Q(
        n19910) );
  OA22X1 U22655 ( .IN1(n23091), .IN2(n21671), .IN3(n23069), .IN4(n22524), .Q(
        n19909) );
  INVX0 U22656 ( .INP(m0s5_data_i[25]), .ZN(n22525) );
  OA22X1 U22657 ( .IN1(n23059), .IN2(n21663), .IN3(n22982), .IN4(n22525), .Q(
        n19908) );
  NAND2X0 U22658 ( .IN1(n29299), .IN2(m0s9_data_i[25]), .QN(n19907) );
  NAND4X0 U22659 ( .IN1(n19910), .IN2(n19909), .IN3(n19908), .IN4(n19907), 
        .QN(n19916) );
  OA22X1 U22660 ( .IN1(n19979), .IN2(n20993), .IN3(n23063), .IN4(n21665), .Q(
        n19914) );
  OA22X1 U22661 ( .IN1(n23003), .IN2(n22119), .IN3(n23085), .IN4(n21662), .Q(
        n19913) );
  OA22X1 U22662 ( .IN1(n23089), .IN2(n22521), .IN3(n23087), .IN4(n22522), .Q(
        n19912) );
  OA22X1 U22663 ( .IN1(n23065), .IN2(n21664), .IN3(n23083), .IN4(n22523), .Q(
        n19911) );
  NAND4X0 U22664 ( .IN1(n19914), .IN2(n19913), .IN3(n19912), .IN4(n19911), 
        .QN(n19915) );
  NOR2X0 U22665 ( .IN1(n19916), .IN2(n19915), .QN(n19918) );
  NAND2X0 U22666 ( .IN1(s15_data_i[25]), .IN2(n19990), .QN(n19917) );
  NAND2X0 U22667 ( .IN1(n19918), .IN2(n19917), .QN(m3_data_o[25]) );
  OA22X1 U22668 ( .IN1(n23003), .IN2(n22539), .IN3(n23083), .IN4(n22540), .Q(
        n19922) );
  OA22X1 U22669 ( .IN1(n23021), .IN2(n21693), .IN3(n23087), .IN4(n21686), .Q(
        n19921) );
  OA22X1 U22670 ( .IN1(n23089), .IN2(n21694), .IN3(n23067), .IN4(n22541), .Q(
        n19920) );
  NAND2X0 U22671 ( .IN1(n29294), .IN2(m0s14_data_i[26]), .QN(n19919) );
  NAND4X0 U22672 ( .IN1(n19922), .IN2(n19921), .IN3(n19920), .IN4(n19919), 
        .QN(n19928) );
  INVX0 U22673 ( .INP(m0s8_data_i[26]), .ZN(n22538) );
  OA22X1 U22674 ( .IN1(n23091), .IN2(n22538), .IN3(n23065), .IN4(n21692), .Q(
        n19926) );
  OA22X1 U22675 ( .IN1(n23059), .IN2(n21682), .IN3(n23085), .IN4(n21695), .Q(
        n19925) );
  OA22X1 U22676 ( .IN1(n19979), .IN2(n21691), .IN3(n22982), .IN4(n21684), .Q(
        n19924) );
  OA22X1 U22677 ( .IN1(n23093), .IN2(n21683), .IN3(n23063), .IN4(n21685), .Q(
        n19923) );
  NAND4X0 U22678 ( .IN1(n19926), .IN2(n19925), .IN3(n19924), .IN4(n19923), 
        .QN(n19927) );
  NOR2X0 U22679 ( .IN1(n19928), .IN2(n19927), .QN(n19930) );
  NAND2X0 U22680 ( .IN1(s15_data_i[26]), .IN2(n19990), .QN(n19929) );
  NAND2X0 U22681 ( .IN1(n19930), .IN2(n19929), .QN(m3_data_o[26]) );
  OA22X1 U22682 ( .IN1(n23003), .IN2(n21715), .IN3(n23085), .IN4(n22910), .Q(
        n19934) );
  OA22X1 U22683 ( .IN1(n23021), .IN2(n21714), .IN3(n23093), .IN4(n22908), .Q(
        n19933) );
  OA22X1 U22684 ( .IN1(n23069), .IN2(n21710), .IN3(n23063), .IN4(n21711), .Q(
        n19932) );
  NAND2X0 U22685 ( .IN1(n29297), .IN2(m0s11_data_i[27]), .QN(n19931) );
  NAND4X0 U22686 ( .IN1(n19934), .IN2(n19933), .IN3(n19932), .IN4(n19931), 
        .QN(n19940) );
  OA22X1 U22687 ( .IN1(n23065), .IN2(n21018), .IN3(n19979), .IN4(n22918), .Q(
        n19938) );
  INVX0 U22688 ( .INP(m0s3_data_i[27]), .ZN(n22912) );
  OA22X1 U22689 ( .IN1(n23091), .IN2(n22913), .IN3(n23089), .IN4(n22912), .Q(
        n19937) );
  OA22X1 U22690 ( .IN1(n23087), .IN2(n22915), .IN3(n23083), .IN4(n22911), .Q(
        n19936) );
  OA22X1 U22691 ( .IN1(n23059), .IN2(n22916), .IN3(n22982), .IN4(n21705), .Q(
        n19935) );
  NAND4X0 U22692 ( .IN1(n19938), .IN2(n19937), .IN3(n19936), .IN4(n19935), 
        .QN(n19939) );
  NOR2X0 U22693 ( .IN1(n19940), .IN2(n19939), .QN(n19942) );
  NAND2X0 U22694 ( .IN1(s15_data_i[27]), .IN2(n19990), .QN(n19941) );
  NAND2X0 U22695 ( .IN1(n19942), .IN2(n19941), .QN(m3_data_o[27]) );
  OA22X1 U22696 ( .IN1(n23069), .IN2(n21725), .IN3(n23063), .IN4(n22938), .Q(
        n19946) );
  OA22X1 U22697 ( .IN1(n23087), .IN2(n22935), .IN3(n23085), .IN4(n22941), .Q(
        n19945) );
  OA22X1 U22698 ( .IN1(n23089), .IN2(n21743), .IN3(n23003), .IN4(n22940), .Q(
        n19944) );
  NAND2X0 U22699 ( .IN1(n29309), .IN2(m0s0_data_i[28]), .QN(n19943) );
  NAND4X0 U22700 ( .IN1(n19946), .IN2(n19945), .IN3(n19944), .IN4(n19943), 
        .QN(n19952) );
  INVX0 U22701 ( .INP(m0s10_data_i[28]), .ZN(n21729) );
  OA22X1 U22702 ( .IN1(n23093), .IN2(n21737), .IN3(n23083), .IN4(n21729), .Q(
        n19950) );
  OA22X1 U22703 ( .IN1(n23091), .IN2(n21739), .IN3(n22982), .IN4(n22936), .Q(
        n19949) );
  OA22X1 U22704 ( .IN1(n23067), .IN2(n22930), .IN3(n23059), .IN4(n21741), .Q(
        n19948) );
  OA22X1 U22705 ( .IN1(n23021), .IN2(n22934), .IN3(n19979), .IN4(n22932), .Q(
        n19947) );
  NAND4X0 U22706 ( .IN1(n19950), .IN2(n19949), .IN3(n19948), .IN4(n19947), 
        .QN(n19951) );
  NOR2X0 U22707 ( .IN1(n19952), .IN2(n19951), .QN(n19954) );
  NAND2X0 U22708 ( .IN1(s15_data_i[28]), .IN2(n19990), .QN(n19953) );
  NAND2X0 U22709 ( .IN1(n19954), .IN2(n19953), .QN(m3_data_o[28]) );
  INVX0 U22710 ( .INP(m0s5_data_i[29]), .ZN(n21040) );
  OA22X1 U22711 ( .IN1(n23065), .IN2(n21043), .IN3(n22982), .IN4(n21040), .Q(
        n19958) );
  OA22X1 U22712 ( .IN1(n23091), .IN2(n21048), .IN3(n23085), .IN4(n22959), .Q(
        n19957) );
  OA22X1 U22713 ( .IN1(n23083), .IN2(n22961), .IN3(n23063), .IN4(n21051), .Q(
        n19956) );
  NAND2X0 U22714 ( .IN1(n29296), .IN2(m0s12_data_i[29]), .QN(n19955) );
  NAND4X0 U22715 ( .IN1(n19958), .IN2(n19957), .IN3(n19956), .IN4(n19955), 
        .QN(n19964) );
  OA22X1 U22716 ( .IN1(n23021), .IN2(n22955), .IN3(n23003), .IN4(n22963), .Q(
        n19962) );
  OA22X1 U22717 ( .IN1(n23089), .IN2(n22953), .IN3(n23069), .IN4(n21050), .Q(
        n19961) );
  OA22X1 U22718 ( .IN1(n23093), .IN2(n22583), .IN3(n23059), .IN4(n21049), .Q(
        n19960) );
  OA22X1 U22719 ( .IN1(n23067), .IN2(n21042), .IN3(n19979), .IN4(n21041), .Q(
        n19959) );
  NAND4X0 U22720 ( .IN1(n19962), .IN2(n19961), .IN3(n19960), .IN4(n19959), 
        .QN(n19963) );
  NOR2X0 U22721 ( .IN1(n19964), .IN2(n19963), .QN(n19966) );
  NAND2X0 U22722 ( .IN1(s15_data_i[29]), .IN2(n19990), .QN(n19965) );
  NAND2X0 U22723 ( .IN1(n19966), .IN2(n19965), .QN(m3_data_o[29]) );
  OA22X1 U22724 ( .IN1(n23085), .IN2(n22601), .IN3(n22982), .IN4(n21072), .Q(
        n19970) );
  INVX0 U22725 ( .INP(m0s9_data_i[30]), .ZN(n21067) );
  OA22X1 U22726 ( .IN1(n23021), .IN2(n21067), .IN3(n23093), .IN4(n21060), .Q(
        n19969) );
  OA22X1 U22727 ( .IN1(n23067), .IN2(n21062), .IN3(n19979), .IN4(n22602), .Q(
        n19968) );
  NAND2X0 U22728 ( .IN1(n29298), .IN2(m0s10_data_i[30]), .QN(n19967) );
  NAND4X0 U22729 ( .IN1(n19970), .IN2(n19969), .IN3(n19968), .IN4(n19967), 
        .QN(n19976) );
  OA22X1 U22730 ( .IN1(n23003), .IN2(n21071), .IN3(n23059), .IN4(n22603), .Q(
        n19974) );
  OA22X1 U22731 ( .IN1(n23089), .IN2(n21070), .IN3(n23065), .IN4(n22177), .Q(
        n19973) );
  OA22X1 U22732 ( .IN1(n23087), .IN2(n22600), .IN3(n23069), .IN4(n22597), .Q(
        n19972) );
  OA22X1 U22733 ( .IN1(n23091), .IN2(n21061), .IN3(n23063), .IN4(n21069), .Q(
        n19971) );
  NAND4X0 U22734 ( .IN1(n19974), .IN2(n19973), .IN3(n19972), .IN4(n19971), 
        .QN(n19975) );
  NOR2X0 U22735 ( .IN1(n19976), .IN2(n19975), .QN(n19978) );
  NAND2X0 U22736 ( .IN1(s15_data_i[30]), .IN2(n19990), .QN(n19977) );
  NAND2X0 U22737 ( .IN1(n19978), .IN2(n19977), .QN(m3_data_o[30]) );
  OA22X1 U22738 ( .IN1(n23085), .IN2(n21099), .IN3(n23063), .IN4(n21105), .Q(
        n19983) );
  OA22X1 U22739 ( .IN1(n23093), .IN2(n21090), .IN3(n19979), .IN4(n22618), .Q(
        n19982) );
  OA22X1 U22740 ( .IN1(n23021), .IN2(n21102), .IN3(n23083), .IN4(n21088), .Q(
        n19981) );
  NAND2X0 U22741 ( .IN1(n29309), .IN2(m0s0_data_i[31]), .QN(n19980) );
  NAND4X0 U22742 ( .IN1(n19983), .IN2(n19982), .IN3(n19981), .IN4(n19980), 
        .QN(n19989) );
  OA22X1 U22743 ( .IN1(n23087), .IN2(n21097), .IN3(n23069), .IN4(n21096), .Q(
        n19987) );
  OA22X1 U22744 ( .IN1(n23091), .IN2(n21083), .IN3(n23067), .IN4(n21086), .Q(
        n19986) );
  OA22X1 U22745 ( .IN1(n23003), .IN2(n21081), .IN3(n22982), .IN4(n22616), .Q(
        n19985) );
  OA22X1 U22746 ( .IN1(n23089), .IN2(n22617), .IN3(n23059), .IN4(n22619), .Q(
        n19984) );
  NAND4X0 U22747 ( .IN1(n19987), .IN2(n19986), .IN3(n19985), .IN4(n19984), 
        .QN(n19988) );
  NOR2X0 U22748 ( .IN1(n19989), .IN2(n19988), .QN(n19992) );
  NAND2X0 U22749 ( .IN1(s15_data_i[31]), .IN2(n19990), .QN(n19991) );
  NAND2X0 U22750 ( .IN1(n19992), .IN2(n19991), .QN(m3_data_o[31]) );
  INVX0 U22751 ( .INP(m2s0_addr[30]), .ZN(n28932) );
  NOR2X0 U22752 ( .IN1(m2s0_addr[31]), .IN2(n28932), .QN(n20013) );
  INVX0 U22753 ( .INP(m2s0_addr[29]), .ZN(n28926) );
  NOR2X0 U22754 ( .IN1(m2s0_addr[28]), .IN2(n28926), .QN(n20010) );
  NAND2X0 U22755 ( .IN1(n20013), .IN2(n20010), .QN(n22964) );
  INVX0 U22756 ( .INP(n22964), .ZN(n29283) );
  NOR2X0 U22757 ( .IN1(n23230), .IN2(n19993), .QN(n29082) );
  NAND2X0 U22758 ( .IN1(n29283), .IN2(n29082), .QN(n26282) );
  INVX0 U22759 ( .INP(s6_rty_i), .ZN(n23429) );
  NOR2X0 U22760 ( .IN1(m2s0_addr[29]), .IN2(m2s0_addr[28]), .QN(n20016) );
  NAND2X0 U22761 ( .IN1(n20016), .IN2(n20013), .QN(n22939) );
  INVX0 U22762 ( .INP(n22939), .ZN(n29285) );
  NOR2X0 U22763 ( .IN1(n23120), .IN2(n19994), .QN(n29037) );
  NAND2X0 U22764 ( .IN1(n29285), .IN2(n29037), .QN(n26894) );
  INVX0 U22765 ( .INP(s4_rty_i), .ZN(n23436) );
  OA22X1 U22766 ( .IN1(n26282), .IN2(n23429), .IN3(n26894), .IN4(n23436), .Q(
        n20003) );
  INVX0 U22767 ( .INP(m2s0_addr[31]), .ZN(n28948) );
  NOR2X0 U22768 ( .IN1(m2s0_addr[30]), .IN2(n28948), .QN(n20009) );
  NAND2X0 U22769 ( .IN1(n20016), .IN2(n20009), .QN(n22914) );
  INVX0 U22770 ( .INP(n22914), .ZN(n29281) );
  NOR2X0 U22771 ( .IN1(n23123), .IN2(n19995), .QN(n29112) );
  NAND2X0 U22772 ( .IN1(n29281), .IN2(n29112), .QN(n25676) );
  INVX0 U22773 ( .INP(s8_rty_i), .ZN(n23428) );
  INVX0 U22774 ( .INP(m2s0_addr[28]), .ZN(n28909) );
  NOR2X0 U22775 ( .IN1(n28926), .IN2(n28909), .QN(n20007) );
  NAND2X0 U22776 ( .IN1(n20007), .IN2(n20009), .QN(n22931) );
  INVX0 U22777 ( .INP(n22931), .ZN(n29278) );
  NOR2X0 U22778 ( .IN1(n23221), .IN2(n19996), .QN(n29164) );
  NAND2X0 U22779 ( .IN1(n29278), .IN2(n29164), .QN(n24765) );
  INVX0 U22780 ( .INP(s11_rty_i), .ZN(n23426) );
  OA22X1 U22781 ( .IN1(n25676), .IN2(n23428), .IN3(n24765), .IN4(n23426), .Q(
        n20002) );
  NOR2X0 U22782 ( .IN1(m2s0_addr[31]), .IN2(m2s0_addr[30]), .QN(n20012) );
  AND2X1 U22783 ( .IN1(n20007), .IN2(n20012), .Q(n29286) );
  NOR2X0 U22784 ( .IN1(n23233), .IN2(n19997), .QN(n29021) );
  NAND2X0 U22785 ( .IN1(n29286), .IN2(n29021), .QN(n27194) );
  INVX0 U22786 ( .INP(s3_rty_i), .ZN(n23427) );
  NOR2X0 U22787 ( .IN1(m2s0_addr[29]), .IN2(n28909), .QN(n20014) );
  NAND2X0 U22788 ( .IN1(n20014), .IN2(n20009), .QN(n22956) );
  INVX0 U22789 ( .INP(n22956), .ZN(n29280) );
  NOR2X0 U22790 ( .IN1(n23117), .IN2(n19998), .QN(n29135) );
  NAND2X0 U22791 ( .IN1(n29280), .IN2(n29135), .QN(n25372) );
  INVX0 U22792 ( .INP(s9_rty_i), .ZN(n23431) );
  OA22X1 U22793 ( .IN1(n27194), .IN2(n23427), .IN3(n25372), .IN4(n23431), .Q(
        n20001) );
  NAND2X0 U22794 ( .IN1(n20012), .IN2(n20010), .QN(n22917) );
  INVX0 U22795 ( .INP(n22917), .ZN(n29287) );
  NOR2X0 U22796 ( .IN1(n23114), .IN2(n19999), .QN(n29003) );
  NAND2X0 U22797 ( .IN1(n29287), .IN2(n29003), .QN(n27503) );
  INVX0 U22798 ( .INP(s2_rty_i), .ZN(n23435) );
  OR2X1 U22799 ( .IN1(n27503), .IN2(n23435), .Q(n20000) );
  NAND4X0 U22800 ( .IN1(n20003), .IN2(n20002), .IN3(n20001), .IN4(n20000), 
        .QN(n20024) );
  NOR2X0 U22801 ( .IN1(n28948), .IN2(n28932), .QN(n20017) );
  NAND2X0 U22802 ( .IN1(n20017), .IN2(n20014), .QN(n22933) );
  INVX0 U22803 ( .INP(n22933), .ZN(n29276) );
  NOR2X0 U22804 ( .IN1(n23212), .IN2(n20004), .QN(n29207) );
  NAND2X0 U22805 ( .IN1(n29276), .IN2(n29207), .QN(n24151) );
  INVX0 U22806 ( .INP(s13_rty_i), .ZN(n23430) );
  NAND2X0 U22807 ( .IN1(n20017), .IN2(n20010), .QN(n22894) );
  INVX0 U22808 ( .INP(n22894), .ZN(n29275) );
  NOR2X0 U22809 ( .IN1(n23240), .IN2(n20005), .QN(n29217) );
  NAND2X0 U22810 ( .IN1(n29275), .IN2(n29217), .QN(n23844) );
  INVX0 U22811 ( .INP(s14_rty_i), .ZN(n23433) );
  OA22X1 U22812 ( .IN1(n24151), .IN2(n23430), .IN3(n23844), .IN4(n23433), .Q(
        n20022) );
  NAND2X0 U22813 ( .IN1(n20012), .IN2(n20016), .QN(n22854) );
  INVX0 U22814 ( .INP(n22854), .ZN(n29290) );
  NOR2X0 U22815 ( .IN1(n23251), .IN2(n20006), .QN(n28975) );
  NAND2X0 U22816 ( .IN1(n29290), .IN2(n28975), .QN(n28109) );
  INVX0 U22817 ( .INP(s0_rty_i), .ZN(n23432) );
  NAND2X0 U22818 ( .IN1(n20007), .IN2(n20013), .QN(n22909) );
  INVX0 U22819 ( .INP(n22909), .ZN(n29282) );
  NOR2X0 U22820 ( .IN1(n23215), .IN2(n20008), .QN(n29091) );
  NAND2X0 U22821 ( .IN1(n29282), .IN2(n29091), .QN(n25982) );
  INVX0 U22822 ( .INP(s7_rty_i), .ZN(n23421) );
  OA22X1 U22823 ( .IN1(n28109), .IN2(n23432), .IN3(n25982), .IN4(n23421), .Q(
        n20021) );
  NAND2X0 U22824 ( .IN1(n20010), .IN2(n20009), .QN(n22962) );
  INVX0 U22825 ( .INP(n22962), .ZN(n29279) );
  NOR2X0 U22826 ( .IN1(n23217), .IN2(n20011), .QN(n29148) );
  NAND2X0 U22827 ( .IN1(n29279), .IN2(n29148), .QN(n25063) );
  INVX0 U22828 ( .INP(s10_rty_i), .ZN(n23422) );
  NAND2X0 U22829 ( .IN1(n20012), .IN2(n20014), .QN(n22960) );
  INVX0 U22830 ( .INP(n23236), .ZN(n23142) );
  AND3X1 U22831 ( .IN1(n23142), .IN2(n23140), .IN3(n21135), .Q(n28985) );
  INVX0 U22832 ( .INP(n28985), .ZN(n28089) );
  NOR2X0 U22833 ( .IN1(n22960), .IN2(n28089), .QN(n20040) );
  INVX0 U22834 ( .INP(n20040), .ZN(n27811) );
  INVX0 U22835 ( .INP(s1_rty_i), .ZN(n23424) );
  OA22X1 U22836 ( .IN1(n25063), .IN2(n23422), .IN3(n27811), .IN4(n23424), .Q(
        n20020) );
  NAND2X0 U22837 ( .IN1(n20014), .IN2(n20013), .QN(n22937) );
  INVX0 U22838 ( .INP(n22937), .ZN(n29284) );
  NOR2X0 U22839 ( .IN1(n23227), .IN2(n20015), .QN(n29055) );
  NAND2X0 U22840 ( .IN1(n29284), .IN2(n29055), .QN(n26592) );
  INVX0 U22841 ( .INP(s5_rty_i), .ZN(n23423) );
  AND2X1 U22842 ( .IN1(n20017), .IN2(n20016), .Q(n29277) );
  NOR2X0 U22843 ( .IN1(n23224), .IN2(n20018), .QN(n29192) );
  NAND2X0 U22844 ( .IN1(n29277), .IN2(n29192), .QN(n24458) );
  INVX0 U22845 ( .INP(s12_rty_i), .ZN(n23425) );
  OA22X1 U22846 ( .IN1(n26592), .IN2(n23423), .IN3(n24458), .IN4(n23425), .Q(
        n20019) );
  NAND4X0 U22847 ( .IN1(n20022), .IN2(n20021), .IN3(n20020), .IN4(n20019), 
        .QN(n20023) );
  NOR2X0 U22848 ( .IN1(n20024), .IN2(n20023), .QN(n20026) );
  AND2X1 U22849 ( .IN1(n20051), .IN2(n23445), .Q(n20037) );
  NAND2X0 U22850 ( .IN1(s15_rty_i), .IN2(n20037), .QN(n20025) );
  NAND2X0 U22851 ( .IN1(n20026), .IN2(n20025), .QN(m2_rty_o) );
  INVX0 U22852 ( .INP(s0_err_i), .ZN(n23405) );
  INVX0 U22853 ( .INP(s3_err_i), .ZN(n23399) );
  OA22X1 U22854 ( .IN1(n28109), .IN2(n23405), .IN3(n27194), .IN4(n23399), .Q(
        n20030) );
  INVX0 U22855 ( .INP(s9_err_i), .ZN(n23401) );
  INVX0 U22856 ( .INP(s11_err_i), .ZN(n23397) );
  OA22X1 U22857 ( .IN1(n25372), .IN2(n23401), .IN3(n24765), .IN4(n23397), .Q(
        n20029) );
  INVX0 U22858 ( .INP(s5_err_i), .ZN(n23404) );
  INVX0 U22859 ( .INP(s14_err_i), .ZN(n23398) );
  OA22X1 U22860 ( .IN1(n26592), .IN2(n23404), .IN3(n23844), .IN4(n23398), .Q(
        n20028) );
  NAND2X0 U22861 ( .IN1(n20040), .IN2(s1_err_i), .QN(n20027) );
  NAND4X0 U22862 ( .IN1(n20030), .IN2(n20029), .IN3(n20028), .IN4(n20027), 
        .QN(n20036) );
  INVX0 U22863 ( .INP(s8_err_i), .ZN(n23394) );
  INVX0 U22864 ( .INP(s10_err_i), .ZN(n23408) );
  OA22X1 U22865 ( .IN1(n25676), .IN2(n23394), .IN3(n25063), .IN4(n23408), .Q(
        n20034) );
  INVX0 U22866 ( .INP(s13_err_i), .ZN(n23402) );
  INVX0 U22867 ( .INP(s12_err_i), .ZN(n23407) );
  OA22X1 U22868 ( .IN1(n24151), .IN2(n23402), .IN3(n24458), .IN4(n23407), .Q(
        n20033) );
  INVX0 U22869 ( .INP(s7_err_i), .ZN(n23406) );
  INVX0 U22870 ( .INP(s6_err_i), .ZN(n23400) );
  OA22X1 U22871 ( .IN1(n25982), .IN2(n23406), .IN3(n26282), .IN4(n23400), .Q(
        n20032) );
  INVX0 U22872 ( .INP(s2_err_i), .ZN(n23396) );
  INVX0 U22873 ( .INP(s4_err_i), .ZN(n23395) );
  OA22X1 U22874 ( .IN1(n27503), .IN2(n23396), .IN3(n26894), .IN4(n23395), .Q(
        n20031) );
  NAND4X0 U22875 ( .IN1(n20034), .IN2(n20033), .IN3(n20032), .IN4(n20031), 
        .QN(n20035) );
  NOR2X0 U22876 ( .IN1(n20036), .IN2(n20035), .QN(n20039) );
  NAND2X0 U22877 ( .IN1(s15_err_i), .IN2(n20037), .QN(n20038) );
  NAND2X0 U22878 ( .IN1(n20039), .IN2(n20038), .QN(m2_err_o) );
  OA22X1 U22879 ( .IN1(n21144), .IN2(n26592), .IN3(n23213), .IN4(n24151), .Q(
        n20044) );
  OA22X1 U22880 ( .IN1(n23253), .IN2(n25372), .IN3(n21123), .IN4(n23844), .Q(
        n20043) );
  OA22X1 U22881 ( .IN1(n21137), .IN2(n24765), .IN3(n21141), .IN4(n24458), .Q(
        n20042) );
  NAND2X0 U22882 ( .IN1(s1_ack_i), .IN2(n20040), .QN(n20041) );
  NAND4X0 U22883 ( .IN1(n20044), .IN2(n20043), .IN3(n20042), .IN4(n20041), 
        .QN(n20050) );
  OA22X1 U22884 ( .IN1(n23252), .IN2(n28109), .IN3(n23219), .IN4(n25063), .Q(
        n20048) );
  OA22X1 U22885 ( .IN1(n23246), .IN2(n25676), .IN3(n23214), .IN4(n27503), .Q(
        n20047) );
  OA22X1 U22886 ( .IN1(n23247), .IN2(n26894), .IN3(n21120), .IN4(n27194), .Q(
        n20046) );
  OA22X1 U22887 ( .IN1(n21126), .IN2(n26282), .IN3(n23220), .IN4(n25982), .Q(
        n20045) );
  NAND4X0 U22888 ( .IN1(n20048), .IN2(n20047), .IN3(n20046), .IN4(n20045), 
        .QN(n20049) );
  NOR2X0 U22889 ( .IN1(n20050), .IN2(n20049), .QN(n20053) );
  NAND2X0 U22890 ( .IN1(n20051), .IN2(n23261), .QN(n20052) );
  NAND2X0 U22891 ( .IN1(n20053), .IN2(n20052), .QN(m2_ack_o) );
  OA22X1 U22892 ( .IN1(n22205), .IN2(n22917), .IN3(n21160), .IN4(n22937), .Q(
        n20057) );
  INVX0 U22893 ( .INP(n29286), .ZN(n22954) );
  OA22X1 U22894 ( .IN1(n21154), .IN2(n22894), .IN3(n22206), .IN4(n22954), .Q(
        n20056) );
  OA22X1 U22895 ( .IN1(n22207), .IN2(n22962), .IN3(n22204), .IN4(n22854), .Q(
        n20055) );
  NAND2X0 U22896 ( .IN1(m0s8_data_i[0]), .IN2(n29281), .QN(n20054) );
  NAND4X0 U22897 ( .IN1(n20057), .IN2(n20056), .IN3(n20055), .IN4(n20054), 
        .QN(n20063) );
  INVX0 U22898 ( .INP(n29277), .ZN(n22958) );
  OA22X1 U22899 ( .IN1(n20251), .IN2(n22958), .IN3(n21162), .IN4(n22909), .Q(
        n20061) );
  OA22X1 U22900 ( .IN1(n21161), .IN2(n22960), .IN3(n22203), .IN4(n22939), .Q(
        n20060) );
  OA22X1 U22901 ( .IN1(n22208), .IN2(n22931), .IN3(n21823), .IN4(n22933), .Q(
        n20059) );
  OA22X1 U22902 ( .IN1(n21153), .IN2(n22964), .IN3(n21159), .IN4(n22956), .Q(
        n20058) );
  NAND4X0 U22903 ( .IN1(n20061), .IN2(n20060), .IN3(n20059), .IN4(n20058), 
        .QN(n20062) );
  NOR2X0 U22904 ( .IN1(n20063), .IN2(n20062), .QN(n20065) );
  INVX0 U22905 ( .INP(n20112), .ZN(n29274) );
  NAND2X0 U22906 ( .IN1(n29274), .IN2(n22218), .QN(n20064) );
  NAND2X0 U22907 ( .IN1(n20065), .IN2(n20064), .QN(m2_data_o[0]) );
  OA22X1 U22908 ( .IN1(n21183), .IN2(n22956), .IN3(n20689), .IN4(n22931), .Q(
        n20069) );
  OA22X1 U22909 ( .IN1(n21186), .IN2(n22962), .IN3(n21173), .IN4(n22939), .Q(
        n20068) );
  OA22X1 U22910 ( .IN1(n22225), .IN2(n22917), .IN3(n21174), .IN4(n22914), .Q(
        n20067) );
  NAND2X0 U22911 ( .IN1(m0s6_data_i[1]), .IN2(n29283), .QN(n20066) );
  NAND4X0 U22912 ( .IN1(n20069), .IN2(n20068), .IN3(n20067), .IN4(n20066), 
        .QN(n20075) );
  OA22X1 U22913 ( .IN1(n21176), .IN2(n22954), .IN3(n22226), .IN4(n22909), .Q(
        n20073) );
  OA22X1 U22914 ( .IN1(n21177), .IN2(n22937), .IN3(n21184), .IN4(n22933), .Q(
        n20072) );
  OA22X1 U22915 ( .IN1(n22224), .IN2(n22894), .IN3(n22223), .IN4(n22854), .Q(
        n20071) );
  OA22X1 U22916 ( .IN1(n21185), .IN2(n22958), .IN3(n21182), .IN4(n22960), .Q(
        n20070) );
  NAND4X0 U22917 ( .IN1(n20073), .IN2(n20072), .IN3(n20071), .IN4(n20070), 
        .QN(n20074) );
  NOR2X0 U22918 ( .IN1(n20075), .IN2(n20074), .QN(n20077) );
  NAND2X0 U22919 ( .IN1(n29274), .IN2(n22235), .QN(n20076) );
  NAND2X0 U22920 ( .IN1(n20077), .IN2(n20076), .QN(m2_data_o[1]) );
  OA22X1 U22921 ( .IN1(n21200), .IN2(n22954), .IN3(n21208), .IN4(n22964), .Q(
        n20081) );
  OA22X1 U22922 ( .IN1(n21212), .IN2(n22933), .IN3(n21207), .IN4(n22917), .Q(
        n20080) );
  OA22X1 U22923 ( .IN1(n21210), .IN2(n22956), .IN3(n21205), .IN4(n22854), .Q(
        n20079) );
  NAND2X0 U22924 ( .IN1(m0s8_data_i[2]), .IN2(n29281), .QN(n20078) );
  NAND4X0 U22925 ( .IN1(n20081), .IN2(n20080), .IN3(n20079), .IN4(n20078), 
        .QN(n20087) );
  OA22X1 U22926 ( .IN1(n21211), .IN2(n22937), .IN3(n21195), .IN4(n22894), .Q(
        n20085) );
  OA22X1 U22927 ( .IN1(n21198), .IN2(n22958), .IN3(n21199), .IN4(n22960), .Q(
        n20084) );
  OA22X1 U22928 ( .IN1(n21197), .IN2(n22939), .IN3(n21206), .IN4(n22962), .Q(
        n20083) );
  OA22X1 U22929 ( .IN1(n21209), .IN2(n22909), .IN3(n20702), .IN4(n22931), .Q(
        n20082) );
  NAND4X0 U22930 ( .IN1(n20085), .IN2(n20084), .IN3(n20083), .IN4(n20082), 
        .QN(n20086) );
  NOR2X0 U22931 ( .IN1(n20087), .IN2(n20086), .QN(n20089) );
  NAND2X0 U22932 ( .IN1(n29274), .IN2(n22247), .QN(n20088) );
  NAND2X0 U22933 ( .IN1(n20089), .IN2(n20088), .QN(m2_data_o[2]) );
  OA22X1 U22934 ( .IN1(n21735), .IN2(n22957), .IN3(n21742), .IN4(n21049), .Q(
        n20093) );
  OA22X1 U22935 ( .IN1(n21736), .IN2(n21040), .IN3(n21745), .IN4(n22963), .Q(
        n20092) );
  OA22X1 U22936 ( .IN1(n21740), .IN2(n21048), .IN3(n21726), .IN4(n21050), .Q(
        n20091) );
  NAND2X0 U22937 ( .IN1(n29343), .IN2(m0s3_data_i[29]), .QN(n20090) );
  NAND4X0 U22938 ( .IN1(n20093), .IN2(n20092), .IN3(n20091), .IN4(n20090), 
        .QN(n20099) );
  OA22X1 U22939 ( .IN1(n21727), .IN2(n22959), .IN3(n21746), .IN4(n22955), .Q(
        n20097) );
  OA22X1 U22940 ( .IN1(n21730), .IN2(n22961), .IN3(n21724), .IN4(n21043), .Q(
        n20096) );
  OA22X1 U22941 ( .IN1(n21738), .IN2(n22583), .IN3(n21704), .IN4(n21041), .Q(
        n20095) );
  OA22X1 U22942 ( .IN1(n21728), .IN2(n21042), .IN3(n21712), .IN4(n21051), .Q(
        n20094) );
  NAND4X0 U22943 ( .IN1(n20097), .IN2(n20096), .IN3(n20095), .IN4(n20094), 
        .QN(n20098) );
  NOR2X0 U22944 ( .IN1(n20099), .IN2(n20098), .QN(n20101) );
  NAND2X0 U22945 ( .IN1(s15_data_i[29]), .IN2(n21753), .QN(n20100) );
  NAND2X0 U22946 ( .IN1(n20101), .IN2(n20100), .QN(m5_data_o[29]) );
  OA22X1 U22947 ( .IN1(n22956), .IN2(n21493), .IN3(n22954), .IN4(n21491), .Q(
        n20105) );
  OA22X1 U22948 ( .IN1(n22909), .IN2(n21500), .IN3(n22937), .IN4(n22009), .Q(
        n20104) );
  OA22X1 U22949 ( .IN1(n22958), .IN2(n22012), .IN3(n22933), .IN4(n22010), .Q(
        n20103) );
  NAND2X0 U22950 ( .IN1(n29290), .IN2(m0s0_data_i[16]), .QN(n20102) );
  NAND4X0 U22951 ( .IN1(n20105), .IN2(n20104), .IN3(n20103), .IN4(n20102), 
        .QN(n20111) );
  OA22X1 U22952 ( .IN1(n22960), .IN2(n21503), .IN3(n22894), .IN4(n21492), .Q(
        n20109) );
  OA22X1 U22953 ( .IN1(n22939), .IN2(n21494), .IN3(n22917), .IN4(n21490), .Q(
        n20108) );
  OA22X1 U22954 ( .IN1(n22931), .IN2(n22011), .IN3(n22914), .IN4(n21499), .Q(
        n20107) );
  OA22X1 U22955 ( .IN1(n22964), .IN2(n21502), .IN3(n22962), .IN4(n21501), .Q(
        n20106) );
  NAND4X0 U22956 ( .IN1(n20109), .IN2(n20108), .IN3(n20107), .IN4(n20106), 
        .QN(n20110) );
  NOR2X0 U22957 ( .IN1(n20111), .IN2(n20110), .QN(n20114) );
  NOR2X0 U22958 ( .IN1(n23501), .IN2(n20112), .QN(n22973) );
  NAND2X0 U22959 ( .IN1(s15_data_i[16]), .IN2(n22973), .QN(n20113) );
  NAND2X0 U22960 ( .IN1(n20114), .IN2(n20113), .QN(m2_data_o[16]) );
  OA22X1 U22961 ( .IN1(n22958), .IN2(n22410), .IN3(n22914), .IN4(n21531), .Q(
        n20118) );
  INVX0 U22962 ( .INP(m0s6_data_i[18]), .ZN(n22412) );
  OA22X1 U22963 ( .IN1(n22964), .IN2(n22412), .IN3(n22954), .IN4(n22413), .Q(
        n20117) );
  OA22X1 U22964 ( .IN1(n22909), .IN2(n22411), .IN3(n22917), .IN4(n21538), .Q(
        n20116) );
  NAND2X0 U22965 ( .IN1(n29278), .IN2(m0s11_data_i[18]), .QN(n20115) );
  NAND4X0 U22966 ( .IN1(n20118), .IN2(n20117), .IN3(n20116), .IN4(n20115), 
        .QN(n20124) );
  OA22X1 U22967 ( .IN1(n22956), .IN2(n21530), .IN3(n22962), .IN4(n21540), .Q(
        n20122) );
  OA22X1 U22968 ( .IN1(n22939), .IN2(n21536), .IN3(n22937), .IN4(n22414), .Q(
        n20121) );
  OA22X1 U22969 ( .IN1(n22933), .IN2(n21539), .IN3(n22894), .IN4(n20901), .Q(
        n20120) );
  OA22X1 U22970 ( .IN1(n22960), .IN2(n22037), .IN3(n22854), .IN4(n22415), .Q(
        n20119) );
  NAND4X0 U22971 ( .IN1(n20122), .IN2(n20121), .IN3(n20120), .IN4(n20119), 
        .QN(n20123) );
  NOR2X0 U22972 ( .IN1(n20124), .IN2(n20123), .QN(n20126) );
  NAND2X0 U22973 ( .IN1(s15_data_i[18]), .IN2(n22973), .QN(n20125) );
  NAND2X0 U22974 ( .IN1(n20126), .IN2(n20125), .QN(m2_data_o[18]) );
  OA22X1 U22975 ( .IN1(n22960), .IN2(n21557), .IN3(n22962), .IN4(n22432), .Q(
        n20130) );
  OA22X1 U22976 ( .IN1(n22958), .IN2(n22434), .IN3(n22937), .IN4(n22050), .Q(
        n20129) );
  OA22X1 U22977 ( .IN1(n22939), .IN2(n21556), .IN3(n22931), .IN4(n21549), .Q(
        n20128) );
  NAND2X0 U22978 ( .IN1(n29283), .IN2(m0s6_data_i[19]), .QN(n20127) );
  NAND4X0 U22979 ( .IN1(n20130), .IN2(n20129), .IN3(n20128), .IN4(n20127), 
        .QN(n20136) );
  OA22X1 U22980 ( .IN1(n22909), .IN2(n22435), .IN3(n22854), .IN4(n22433), .Q(
        n20134) );
  OA22X1 U22981 ( .IN1(n22956), .IN2(n22429), .IN3(n22917), .IN4(n21558), .Q(
        n20133) );
  OA22X1 U22982 ( .IN1(n22933), .IN2(n22430), .IN3(n22954), .IN4(n22431), .Q(
        n20132) );
  OA22X1 U22983 ( .IN1(n22914), .IN2(n21550), .IN3(n22894), .IN4(n22428), .Q(
        n20131) );
  NAND4X0 U22984 ( .IN1(n20134), .IN2(n20133), .IN3(n20132), .IN4(n20131), 
        .QN(n20135) );
  NOR2X0 U22985 ( .IN1(n20136), .IN2(n20135), .QN(n20138) );
  NAND2X0 U22986 ( .IN1(s15_data_i[19]), .IN2(n22973), .QN(n20137) );
  NAND2X0 U22987 ( .IN1(n20138), .IN2(n20137), .QN(m2_data_o[19]) );
  OA22X1 U22988 ( .IN1(n22933), .IN2(n21567), .IN3(n22854), .IN4(n22451), .Q(
        n20142) );
  OA22X1 U22989 ( .IN1(n22958), .IN2(n22449), .IN3(n22962), .IN4(n21574), .Q(
        n20141) );
  OA22X1 U22990 ( .IN1(n22909), .IN2(n21576), .IN3(n22937), .IN4(n22448), .Q(
        n20140) );
  NAND2X0 U22991 ( .IN1(n29275), .IN2(m0s14_data_i[20]), .QN(n20139) );
  NAND4X0 U22992 ( .IN1(n20142), .IN2(n20141), .IN3(n20140), .IN4(n20139), 
        .QN(n20148) );
  OA22X1 U22993 ( .IN1(n22960), .IN2(n21575), .IN3(n22931), .IN4(n22450), .Q(
        n20146) );
  OA22X1 U22994 ( .IN1(n22964), .IN2(n22454), .IN3(n22954), .IN4(n21568), .Q(
        n20145) );
  OA22X1 U22995 ( .IN1(n22956), .IN2(n22447), .IN3(n22914), .IN4(n21573), .Q(
        n20144) );
  OA22X1 U22996 ( .IN1(n22939), .IN2(n21577), .IN3(n22917), .IN4(n22452), .Q(
        n20143) );
  NAND4X0 U22997 ( .IN1(n20146), .IN2(n20145), .IN3(n20144), .IN4(n20143), 
        .QN(n20147) );
  NOR2X0 U22998 ( .IN1(n20148), .IN2(n20147), .QN(n20150) );
  NAND2X0 U22999 ( .IN1(s15_data_i[20]), .IN2(n22973), .QN(n20149) );
  NAND2X0 U23000 ( .IN1(n20150), .IN2(n20149), .QN(m2_data_o[20]) );
  OA22X1 U23001 ( .IN1(n22956), .IN2(n21633), .IN3(n22914), .IN4(n22492), .Q(
        n20154) );
  OA22X1 U23002 ( .IN1(n22939), .IN2(n20968), .IN3(n22962), .IN4(n22494), .Q(
        n20153) );
  OA22X1 U23003 ( .IN1(n22933), .IN2(n21632), .IN3(n22894), .IN4(n21621), .Q(
        n20152) );
  NAND2X0 U23004 ( .IN1(n29284), .IN2(m0s5_data_i[23]), .QN(n20151) );
  NAND4X0 U23005 ( .IN1(n20154), .IN2(n20153), .IN3(n20152), .IN4(n20151), 
        .QN(n20160) );
  OA22X1 U23006 ( .IN1(n22958), .IN2(n21622), .IN3(n22964), .IN4(n21625), .Q(
        n20158) );
  OA22X1 U23007 ( .IN1(n22909), .IN2(n22495), .IN3(n22917), .IN4(n21623), .Q(
        n20157) );
  OA22X1 U23008 ( .IN1(n22960), .IN2(n22491), .IN3(n22954), .IN4(n21631), .Q(
        n20156) );
  OA22X1 U23009 ( .IN1(n22931), .IN2(n21630), .IN3(n22854), .IN4(n21634), .Q(
        n20155) );
  NAND4X0 U23010 ( .IN1(n20158), .IN2(n20157), .IN3(n20156), .IN4(n20155), 
        .QN(n20159) );
  NOR2X0 U23011 ( .IN1(n20160), .IN2(n20159), .QN(n20162) );
  NAND2X0 U23012 ( .IN1(s15_data_i[23]), .IN2(n22973), .QN(n20161) );
  NAND2X0 U23013 ( .IN1(n20162), .IN2(n20161), .QN(m2_data_o[23]) );
  OA22X1 U23014 ( .IN1(n22960), .IN2(n21662), .IN3(n22914), .IN4(n21671), .Q(
        n20166) );
  OA22X1 U23015 ( .IN1(n22909), .IN2(n21672), .IN3(n22937), .IN4(n22525), .Q(
        n20165) );
  OA22X1 U23016 ( .IN1(n22939), .IN2(n21665), .IN3(n22958), .IN4(n22522), .Q(
        n20164) );
  NAND2X0 U23017 ( .IN1(n29279), .IN2(m0s10_data_i[25]), .QN(n20163) );
  NAND4X0 U23018 ( .IN1(n20166), .IN2(n20165), .IN3(n20164), .IN4(n20163), 
        .QN(n20172) );
  OA22X1 U23019 ( .IN1(n22956), .IN2(n22520), .IN3(n22917), .IN4(n21663), .Q(
        n20170) );
  OA22X1 U23020 ( .IN1(n22894), .IN2(n22524), .IN3(n22954), .IN4(n22521), .Q(
        n20169) );
  OA22X1 U23021 ( .IN1(n22931), .IN2(n21670), .IN3(n22854), .IN4(n21664), .Q(
        n20168) );
  OA22X1 U23022 ( .IN1(n22964), .IN2(n22119), .IN3(n22933), .IN4(n20993), .Q(
        n20167) );
  NAND4X0 U23023 ( .IN1(n20170), .IN2(n20169), .IN3(n20168), .IN4(n20167), 
        .QN(n20171) );
  NOR2X0 U23024 ( .IN1(n20172), .IN2(n20171), .QN(n20174) );
  NAND2X0 U23025 ( .IN1(s15_data_i[25]), .IN2(n22973), .QN(n20173) );
  NAND2X0 U23026 ( .IN1(n20174), .IN2(n20173), .QN(m2_data_o[25]) );
  OA22X1 U23027 ( .IN1(n22964), .IN2(n22539), .IN3(n22937), .IN4(n21684), .Q(
        n20178) );
  OA22X1 U23028 ( .IN1(n22960), .IN2(n21695), .IN3(n22954), .IN4(n21694), .Q(
        n20177) );
  OA22X1 U23029 ( .IN1(n22939), .IN2(n21685), .IN3(n22914), .IN4(n22538), .Q(
        n20176) );
  NAND2X0 U23030 ( .IN1(n29287), .IN2(m0s2_data_i[26]), .QN(n20175) );
  NAND4X0 U23031 ( .IN1(n20178), .IN2(n20177), .IN3(n20176), .IN4(n20175), 
        .QN(n20184) );
  OA22X1 U23032 ( .IN1(n22933), .IN2(n21691), .IN3(n22854), .IN4(n21692), .Q(
        n20182) );
  OA22X1 U23033 ( .IN1(n22958), .IN2(n21686), .IN3(n22931), .IN4(n22541), .Q(
        n20181) );
  OA22X1 U23034 ( .IN1(n22956), .IN2(n21693), .IN3(n22962), .IN4(n22540), .Q(
        n20180) );
  OA22X1 U23035 ( .IN1(n22909), .IN2(n21683), .IN3(n22894), .IN4(n21681), .Q(
        n20179) );
  NAND4X0 U23036 ( .IN1(n20182), .IN2(n20181), .IN3(n20180), .IN4(n20179), 
        .QN(n20183) );
  NOR2X0 U23037 ( .IN1(n20184), .IN2(n20183), .QN(n20186) );
  NAND2X0 U23038 ( .IN1(s15_data_i[26]), .IN2(n22973), .QN(n20185) );
  NAND2X0 U23039 ( .IN1(n20186), .IN2(n20185), .QN(m2_data_o[26]) );
  OA22X1 U23040 ( .IN1(n22939), .IN2(n21069), .IN3(n22958), .IN4(n22600), .Q(
        n20190) );
  OA22X1 U23041 ( .IN1(n22933), .IN2(n22602), .IN3(n22914), .IN4(n21061), .Q(
        n20189) );
  OA22X1 U23042 ( .IN1(n22956), .IN2(n21067), .IN3(n22931), .IN4(n21062), .Q(
        n20188) );
  NAND2X0 U23043 ( .IN1(n29287), .IN2(m0s2_data_i[30]), .QN(n20187) );
  NAND4X0 U23044 ( .IN1(n20190), .IN2(n20189), .IN3(n20188), .IN4(n20187), 
        .QN(n20196) );
  OA22X1 U23045 ( .IN1(n22954), .IN2(n21070), .IN3(n22854), .IN4(n22177), .Q(
        n20194) );
  OA22X1 U23046 ( .IN1(n22960), .IN2(n22601), .IN3(n22894), .IN4(n22597), .Q(
        n20193) );
  OA22X1 U23047 ( .IN1(n22909), .IN2(n21060), .IN3(n22964), .IN4(n21071), .Q(
        n20192) );
  OA22X1 U23048 ( .IN1(n22937), .IN2(n21072), .IN3(n22962), .IN4(n22598), .Q(
        n20191) );
  NAND4X0 U23049 ( .IN1(n20194), .IN2(n20193), .IN3(n20192), .IN4(n20191), 
        .QN(n20195) );
  NOR2X0 U23050 ( .IN1(n20196), .IN2(n20195), .QN(n20198) );
  NAND2X0 U23051 ( .IN1(s15_data_i[30]), .IN2(n22973), .QN(n20197) );
  NAND2X0 U23052 ( .IN1(n20198), .IN2(n20197), .QN(m2_data_o[30]) );
  OA22X1 U23053 ( .IN1(n22937), .IN2(n22616), .IN3(n22962), .IN4(n21088), .Q(
        n20202) );
  OA22X1 U23054 ( .IN1(n22956), .IN2(n21102), .IN3(n22933), .IN4(n22618), .Q(
        n20201) );
  OA22X1 U23055 ( .IN1(n22909), .IN2(n21090), .IN3(n22894), .IN4(n21096), .Q(
        n20200) );
  NAND2X0 U23056 ( .IN1(n29281), .IN2(m0s8_data_i[31]), .QN(n20199) );
  NAND4X0 U23057 ( .IN1(n20202), .IN2(n20201), .IN3(n20200), .IN4(n20199), 
        .QN(n20208) );
  OA22X1 U23058 ( .IN1(n22939), .IN2(n21105), .IN3(n22958), .IN4(n21097), .Q(
        n20206) );
  OA22X1 U23059 ( .IN1(n22960), .IN2(n21099), .IN3(n22917), .IN4(n22619), .Q(
        n20205) );
  OA22X1 U23060 ( .IN1(n22964), .IN2(n21081), .IN3(n22954), .IN4(n22617), .Q(
        n20204) );
  OA22X1 U23061 ( .IN1(n22931), .IN2(n21086), .IN3(n22854), .IN4(n21107), .Q(
        n20203) );
  NAND4X0 U23062 ( .IN1(n20206), .IN2(n20205), .IN3(n20204), .IN4(n20203), 
        .QN(n20207) );
  NOR2X0 U23063 ( .IN1(n20208), .IN2(n20207), .QN(n20210) );
  NAND2X0 U23064 ( .IN1(s15_data_i[31]), .IN2(n22973), .QN(n20209) );
  NAND2X0 U23065 ( .IN1(n20210), .IN2(n20209), .QN(m2_data_o[31]) );
  NAND2X0 U23066 ( .IN1(m1s0_addr[31]), .IN2(m1s0_addr[30]), .QN(n20215) );
  INVX0 U23067 ( .INP(m1s0_addr[29]), .ZN(n28924) );
  NAND2X0 U23068 ( .IN1(m1s0_addr[28]), .IN2(n28924), .QN(n20219) );
  NOR2X0 U23069 ( .IN1(n20215), .IN2(n20219), .QN(n29257) );
  INVX0 U23070 ( .INP(n29257), .ZN(n22554) );
  INVX0 U23071 ( .INP(m1s0_addr[30]), .ZN(n28935) );
  NAND2X0 U23072 ( .IN1(m1s0_addr[31]), .IN2(n28935), .QN(n20221) );
  OR2X1 U23073 ( .IN1(n20219), .IN2(n20221), .Q(n22582) );
  OA22X1 U23074 ( .IN1(n22554), .IN2(n22010), .IN3(n22582), .IN4(n21493), .Q(
        n20214) );
  INVX0 U23075 ( .INP(m1s0_addr[28]), .ZN(n28911) );
  NAND2X0 U23076 ( .IN1(n28924), .IN2(n28911), .QN(n20218) );
  INVX0 U23077 ( .INP(m1s0_addr[31]), .ZN(n28952) );
  NAND2X0 U23078 ( .IN1(n28952), .IN2(m1s0_addr[30]), .QN(n20216) );
  OR2X1 U23079 ( .IN1(n20218), .IN2(n20216), .Q(n22567) );
  NAND2X0 U23080 ( .IN1(m1s0_addr[29]), .IN2(m1s0_addr[28]), .QN(n20222) );
  OR2X1 U23081 ( .IN1(n20222), .IN2(n20216), .Q(n22584) );
  OA22X1 U23082 ( .IN1(n22567), .IN2(n21494), .IN3(n22584), .IN4(n21500), .Q(
        n20213) );
  NAND2X0 U23083 ( .IN1(n28952), .IN2(n28935), .QN(n20220) );
  NAND2X0 U23084 ( .IN1(n28911), .IN2(m1s0_addr[29]), .QN(n20217) );
  OR2X1 U23085 ( .IN1(n20220), .IN2(n20217), .Q(n22620) );
  OR2X1 U23086 ( .IN1(n20215), .IN2(n20218), .Q(n23226) );
  OA22X1 U23087 ( .IN1(n22620), .IN2(n21490), .IN3(n23226), .IN4(n22012), .Q(
        n20212) );
  NOR2X0 U23088 ( .IN1(n20220), .IN2(n20218), .QN(n29271) );
  NAND2X0 U23089 ( .IN1(n29271), .IN2(m0s0_data_i[16]), .QN(n20211) );
  NAND4X0 U23090 ( .IN1(n20214), .IN2(n20213), .IN3(n20212), .IN4(n20211), 
        .QN(n20228) );
  NOR2X0 U23091 ( .IN1(n20222), .IN2(n20220), .QN(n29267) );
  INVX0 U23092 ( .INP(n29267), .ZN(n23235) );
  OR2X1 U23093 ( .IN1(n20215), .IN2(n20217), .Q(n23241) );
  OA22X1 U23094 ( .IN1(n23235), .IN2(n21491), .IN3(n23241), .IN4(n21492), .Q(
        n20226) );
  NOR2X0 U23095 ( .IN1(n20216), .IN2(n20219), .QN(n29265) );
  INVX0 U23096 ( .INP(n29265), .ZN(n23229) );
  OR2X1 U23097 ( .IN1(n20217), .IN2(n20221), .Q(n22599) );
  OA22X1 U23098 ( .IN1(n23229), .IN2(n22009), .IN3(n22599), .IN4(n21501), .Q(
        n20225) );
  OR2X1 U23099 ( .IN1(n20217), .IN2(n20216), .Q(n23232) );
  NOR2X0 U23100 ( .IN1(n20218), .IN2(n20221), .QN(n29262) );
  OA22X1 U23101 ( .IN1(n23232), .IN2(n21502), .IN3(n22493), .IN4(n21499), .Q(
        n20224) );
  OR2X1 U23102 ( .IN1(n20220), .IN2(n20219), .Q(n23238) );
  NOR2X0 U23103 ( .IN1(n20222), .IN2(n20221), .QN(n29259) );
  INVX0 U23104 ( .INP(n29259), .ZN(n23223) );
  OA22X1 U23105 ( .IN1(n23238), .IN2(n21503), .IN3(n23223), .IN4(n22011), .Q(
        n20223) );
  NAND4X0 U23106 ( .IN1(n20226), .IN2(n20225), .IN3(n20224), .IN4(n20223), 
        .QN(n20227) );
  NOR2X0 U23107 ( .IN1(n20228), .IN2(n20227), .QN(n20230) );
  NOR2X0 U23108 ( .IN1(n23501), .IN2(n22217), .QN(n22629) );
  NAND2X0 U23109 ( .IN1(s15_data_i[16]), .IN2(n22629), .QN(n20229) );
  NAND2X0 U23110 ( .IN1(n20230), .IN2(n20229), .QN(m1_data_o[16]) );
  INVX0 U23111 ( .INP(m7s0_addr[28]), .ZN(n28913) );
  NOR2X0 U23112 ( .IN1(m7s0_addr[29]), .IN2(n28913), .QN(n20237) );
  INVX0 U23113 ( .INP(m7s0_addr[30]), .ZN(n28933) );
  NOR2X0 U23114 ( .IN1(m7s0_addr[31]), .IN2(n28933), .QN(n20241) );
  AND2X1 U23115 ( .IN1(n20237), .IN2(n20241), .Q(n29379) );
  NAND3X0 U23116 ( .IN1(n23133), .IN2(n23227), .IN3(n23132), .QN(n26833) );
  NAND2X0 U23117 ( .IN1(n29379), .IN2(n29065), .QN(n26587) );
  INVX0 U23118 ( .INP(m7s0_addr[31]), .ZN(n28960) );
  NOR2X0 U23119 ( .IN1(n28960), .IN2(n28933), .QN(n20231) );
  AND2X1 U23120 ( .IN1(n20231), .IN2(n20237), .Q(n29371) );
  NAND3X0 U23121 ( .IN1(n23212), .IN2(n23129), .IN3(n23128), .QN(n24397) );
  NAND2X0 U23122 ( .IN1(n29371), .IN2(n29201), .QN(n24149) );
  OA22X1 U23123 ( .IN1(n21144), .IN2(n26587), .IN3(n23213), .IN4(n24149), .Q(
        n20235) );
  INVX0 U23124 ( .INP(m7s0_addr[29]), .ZN(n28921) );
  NOR2X0 U23125 ( .IN1(m7s0_addr[28]), .IN2(n28921), .QN(n20236) );
  AND2X1 U23126 ( .IN1(n20236), .IN2(n20241), .Q(n29378) );
  NAND3X0 U23127 ( .IN1(n23230), .IN2(n23137), .IN3(n23136), .QN(n26527) );
  NAND2X0 U23128 ( .IN1(n29378), .IN2(n29075), .QN(n26286) );
  NOR2X0 U23129 ( .IN1(m7s0_addr[28]), .IN2(m7s0_addr[29]), .QN(n20240) );
  AND2X1 U23130 ( .IN1(n20231), .IN2(n20240), .Q(n29372) );
  NAND3X0 U23131 ( .IN1(n23151), .IN2(n23224), .IN3(n23150), .QN(n24701) );
  NAND2X0 U23132 ( .IN1(n29372), .IN2(n29190), .QN(n24460) );
  OA22X1 U23133 ( .IN1(n21126), .IN2(n26286), .IN3(n21141), .IN4(n24460), .Q(
        n20234) );
  NOR2X0 U23134 ( .IN1(m7s0_addr[31]), .IN2(m7s0_addr[30]), .QN(n20238) );
  AND2X1 U23135 ( .IN1(n20238), .IN2(n20236), .Q(n29382) );
  NAND3X0 U23136 ( .IN1(n23114), .IN2(n23113), .IN3(n23112), .QN(n27747) );
  NAND2X0 U23137 ( .IN1(n29382), .IN2(n29004), .QN(n27505) );
  AND2X1 U23138 ( .IN1(n20238), .IN2(n20240), .Q(n29385) );
  NAND3X0 U23139 ( .IN1(n23251), .IN2(n23155), .IN3(n23154), .QN(n28830) );
  NAND2X0 U23140 ( .IN1(n29385), .IN2(n28976), .QN(n28111) );
  OA22X1 U23141 ( .IN1(n23214), .IN2(n27505), .IN3(n23252), .IN4(n28111), .Q(
        n20233) );
  AND2X1 U23142 ( .IN1(n20231), .IN2(n20236), .Q(n29370) );
  INVX0 U23143 ( .INP(n29370), .ZN(n20614) );
  AND3X1 U23144 ( .IN1(n23240), .IN2(n23125), .IN3(n23124), .Q(n29228) );
  INVX0 U23145 ( .INP(n29228), .ZN(n24136) );
  NOR2X0 U23146 ( .IN1(n20614), .IN2(n24136), .QN(n23845) );
  NAND2X0 U23147 ( .IN1(s14_ack_i), .IN2(n23845), .QN(n20232) );
  NAND4X0 U23148 ( .IN1(n20235), .IN2(n20234), .IN3(n20233), .IN4(n20232), 
        .QN(n20248) );
  AND2X1 U23149 ( .IN1(n20240), .IN2(n20241), .Q(n29380) );
  NAND3X0 U23150 ( .IN1(n23120), .IN2(n23119), .IN3(n23118), .QN(n27137) );
  NAND2X0 U23151 ( .IN1(n29380), .IN2(n29047), .QN(n26890) );
  NOR2X0 U23152 ( .IN1(n28913), .IN2(n28921), .QN(n20242) );
  NOR2X0 U23153 ( .IN1(m7s0_addr[30]), .IN2(n28960), .QN(n20239) );
  AND2X1 U23154 ( .IN1(n20242), .IN2(n20239), .Q(n29373) );
  NAND3X0 U23155 ( .IN1(n23147), .IN2(n23146), .IN3(n23221), .QN(n25006) );
  NAND2X0 U23156 ( .IN1(n29373), .IN2(n29174), .QN(n24763) );
  OA22X1 U23157 ( .IN1(n23247), .IN2(n26890), .IN3(n21137), .IN4(n24763), .Q(
        n20246) );
  AND2X1 U23158 ( .IN1(n20238), .IN2(n20237), .Q(n29383) );
  NAND3X0 U23159 ( .IN1(n23141), .IN2(n23236), .IN3(n23140), .QN(n28057) );
  NAND2X0 U23160 ( .IN1(n29383), .IN2(n28994), .QN(n27809) );
  NAND2X0 U23161 ( .IN1(n20236), .IN2(n20239), .QN(n20630) );
  INVX0 U23162 ( .INP(n20630), .ZN(n29374) );
  AND3X1 U23163 ( .IN1(n23159), .IN2(n23217), .IN3(n23158), .Q(n29146) );
  NAND2X0 U23164 ( .IN1(n29374), .IN2(n29146), .QN(n25070) );
  OA22X1 U23165 ( .IN1(n21138), .IN2(n27809), .IN3(n23219), .IN4(n25070), .Q(
        n20245) );
  AND2X1 U23166 ( .IN1(n20237), .IN2(n20239), .Q(n29375) );
  NAND3X0 U23167 ( .IN1(n23116), .IN2(n23117), .IN3(n23115), .QN(n25619) );
  NAND2X0 U23168 ( .IN1(n29375), .IN2(n29129), .QN(n25368) );
  AND2X1 U23169 ( .IN1(n20242), .IN2(n20238), .Q(n29381) );
  NAND3X0 U23170 ( .IN1(n23233), .IN2(n23165), .IN3(n23164), .QN(n27443) );
  NAND2X0 U23171 ( .IN1(n29381), .IN2(n29020), .QN(n27201) );
  OA22X1 U23172 ( .IN1(n23253), .IN2(n25368), .IN3(n21120), .IN4(n27201), .Q(
        n20244) );
  NAND2X0 U23173 ( .IN1(n20240), .IN2(n20239), .QN(n20628) );
  INVX0 U23174 ( .INP(n20628), .ZN(n29376) );
  AND3X1 U23175 ( .IN1(n23123), .IN2(n23122), .IN3(n23121), .Q(n29111) );
  NAND2X0 U23176 ( .IN1(n29376), .IN2(n29111), .QN(n25674) );
  NAND2X0 U23177 ( .IN1(n20242), .IN2(n20241), .QN(n20636) );
  INVX0 U23178 ( .INP(n20636), .ZN(n29377) );
  AND3X1 U23179 ( .IN1(n23144), .IN2(n23215), .IN3(n23143), .Q(n29102) );
  NAND2X0 U23180 ( .IN1(n29377), .IN2(n29102), .QN(n25981) );
  OA22X1 U23181 ( .IN1(n23246), .IN2(n25674), .IN3(n23220), .IN4(n25981), .Q(
        n20243) );
  NAND4X0 U23182 ( .IN1(n20246), .IN2(n20245), .IN3(n20244), .IN4(n20243), 
        .QN(n20247) );
  NOR2X0 U23183 ( .IN1(n20248), .IN2(n20247), .QN(n20250) );
  NAND2X0 U23184 ( .IN1(n23446), .IN2(n23261), .QN(n20249) );
  NAND2X0 U23185 ( .IN1(n20250), .IN2(n20249), .QN(m7_ack_o) );
  INVX0 U23186 ( .INP(n29375), .ZN(n20629) );
  OA22X1 U23187 ( .IN1(n22207), .IN2(n20630), .IN3(n21159), .IN4(n20629), .Q(
        n20255) );
  INVX0 U23188 ( .INP(n29372), .ZN(n20643) );
  OA22X1 U23189 ( .IN1(n20251), .IN2(n20643), .IN3(n21154), .IN4(n20614), .Q(
        n20254) );
  INVX0 U23190 ( .INP(n29378), .ZN(n20642) );
  OA22X1 U23191 ( .IN1(n21153), .IN2(n20642), .IN3(n21163), .IN4(n20628), .Q(
        n20253) );
  NAND2X0 U23192 ( .IN1(m0s0_data_i[0]), .IN2(n29385), .QN(n20252) );
  NAND4X0 U23193 ( .IN1(n20255), .IN2(n20254), .IN3(n20253), .IN4(n20252), 
        .QN(n20261) );
  INVX0 U23194 ( .INP(n29383), .ZN(n20639) );
  INVX0 U23195 ( .INP(n29380), .ZN(n20637) );
  OA22X1 U23196 ( .IN1(n21161), .IN2(n20639), .IN3(n22203), .IN4(n20637), .Q(
        n20259) );
  INVX0 U23197 ( .INP(n29371), .ZN(n20640) );
  INVX0 U23198 ( .INP(n29382), .ZN(n20641) );
  OA22X1 U23199 ( .IN1(n21823), .IN2(n20640), .IN3(n22205), .IN4(n20641), .Q(
        n20258) );
  INVX0 U23200 ( .INP(n29373), .ZN(n20627) );
  INVX0 U23201 ( .INP(n29379), .ZN(n20631) );
  OA22X1 U23202 ( .IN1(n22208), .IN2(n20627), .IN3(n21160), .IN4(n20631), .Q(
        n20257) );
  INVX0 U23203 ( .INP(n29381), .ZN(n20638) );
  OA22X1 U23204 ( .IN1(n22206), .IN2(n20638), .IN3(n21162), .IN4(n20636), .Q(
        n20256) );
  NAND4X0 U23205 ( .IN1(n20259), .IN2(n20258), .IN3(n20257), .IN4(n20256), 
        .QN(n20260) );
  NOR2X0 U23206 ( .IN1(n20261), .IN2(n20260), .QN(n20263) );
  INVX0 U23207 ( .INP(n20454), .ZN(n29369) );
  NAND2X0 U23208 ( .IN1(n29369), .IN2(n22218), .QN(n20262) );
  NAND2X0 U23209 ( .IN1(n20263), .IN2(n20262), .QN(m7_data_o[0]) );
  INVX0 U23210 ( .INP(n29385), .ZN(n20553) );
  OA22X1 U23211 ( .IN1(n21174), .IN2(n20628), .IN3(n22223), .IN4(n20553), .Q(
        n20267) );
  OA22X1 U23212 ( .IN1(n22226), .IN2(n20636), .IN3(n21184), .IN4(n20640), .Q(
        n20266) );
  OA22X1 U23213 ( .IN1(n21182), .IN2(n20639), .IN3(n21173), .IN4(n20637), .Q(
        n20265) );
  NAND2X0 U23214 ( .IN1(m0s3_data_i[1]), .IN2(n29381), .QN(n20264) );
  NAND4X0 U23215 ( .IN1(n20267), .IN2(n20266), .IN3(n20265), .IN4(n20264), 
        .QN(n20273) );
  OA22X1 U23216 ( .IN1(n21175), .IN2(n20642), .IN3(n21186), .IN4(n20630), .Q(
        n20271) );
  OA22X1 U23217 ( .IN1(n22224), .IN2(n20614), .IN3(n21183), .IN4(n20629), .Q(
        n20270) );
  OA22X1 U23218 ( .IN1(n21177), .IN2(n20631), .IN3(n21185), .IN4(n20643), .Q(
        n20269) );
  OA22X1 U23219 ( .IN1(n22225), .IN2(n20641), .IN3(n20689), .IN4(n20627), .Q(
        n20268) );
  NAND4X0 U23220 ( .IN1(n20271), .IN2(n20270), .IN3(n20269), .IN4(n20268), 
        .QN(n20272) );
  NOR2X0 U23221 ( .IN1(n20273), .IN2(n20272), .QN(n20275) );
  NAND2X0 U23222 ( .IN1(n29369), .IN2(n22235), .QN(n20274) );
  NAND2X0 U23223 ( .IN1(n20275), .IN2(n20274), .QN(m7_data_o[1]) );
  OA22X1 U23224 ( .IN1(n21208), .IN2(n20642), .IN3(n21199), .IN4(n20639), .Q(
        n20279) );
  OA22X1 U23225 ( .IN1(n21196), .IN2(n20628), .IN3(n21205), .IN4(n20553), .Q(
        n20278) );
  OA22X1 U23226 ( .IN1(n21198), .IN2(n20643), .IN3(n21200), .IN4(n20638), .Q(
        n20277) );
  NAND2X0 U23227 ( .IN1(m0s2_data_i[2]), .IN2(n29382), .QN(n20276) );
  NAND4X0 U23228 ( .IN1(n20279), .IN2(n20278), .IN3(n20277), .IN4(n20276), 
        .QN(n20285) );
  OA22X1 U23229 ( .IN1(n21212), .IN2(n20640), .IN3(n21211), .IN4(n20631), .Q(
        n20283) );
  OA22X1 U23230 ( .IN1(n21210), .IN2(n20629), .IN3(n21195), .IN4(n20614), .Q(
        n20282) );
  OA22X1 U23231 ( .IN1(n21206), .IN2(n20630), .IN3(n20702), .IN4(n20627), .Q(
        n20281) );
  OA22X1 U23232 ( .IN1(n21209), .IN2(n20636), .IN3(n21197), .IN4(n20637), .Q(
        n20280) );
  NAND4X0 U23233 ( .IN1(n20283), .IN2(n20282), .IN3(n20281), .IN4(n20280), 
        .QN(n20284) );
  NOR2X0 U23234 ( .IN1(n20285), .IN2(n20284), .QN(n20287) );
  NAND2X0 U23235 ( .IN1(n29369), .IN2(n22247), .QN(n20286) );
  NAND2X0 U23236 ( .IN1(n20287), .IN2(n20286), .QN(m7_data_o[2]) );
  OA22X1 U23237 ( .IN1(n22636), .IN2(n20640), .IN3(n21235), .IN4(n20553), .Q(
        n20291) );
  OA22X1 U23238 ( .IN1(n21234), .IN2(n20627), .IN3(n21233), .IN4(n20628), .Q(
        n20290) );
  OA22X1 U23239 ( .IN1(n21221), .IN2(n20638), .IN3(n21226), .IN4(n20639), .Q(
        n20289) );
  NAND2X0 U23240 ( .IN1(m0s10_data_i[3]), .IN2(n29374), .QN(n20288) );
  NAND4X0 U23241 ( .IN1(n20291), .IN2(n20290), .IN3(n20289), .IN4(n20288), 
        .QN(n20297) );
  OA22X1 U23242 ( .IN1(n21223), .IN2(n20629), .IN3(n21231), .IN4(n20614), .Q(
        n20295) );
  OA22X1 U23243 ( .IN1(n22637), .IN2(n20631), .IN3(n21225), .IN4(n20641), .Q(
        n20294) );
  OA22X1 U23244 ( .IN1(n22635), .IN2(n20643), .IN3(n22634), .IN4(n20637), .Q(
        n20293) );
  OA22X1 U23245 ( .IN1(n21222), .IN2(n20636), .IN3(n21224), .IN4(n20642), .Q(
        n20292) );
  NAND4X0 U23246 ( .IN1(n20295), .IN2(n20294), .IN3(n20293), .IN4(n20292), 
        .QN(n20296) );
  NOR2X0 U23247 ( .IN1(n20297), .IN2(n20296), .QN(n20299) );
  NAND2X0 U23248 ( .IN1(n29369), .IN2(n22646), .QN(n20298) );
  NAND2X0 U23249 ( .IN1(n20299), .IN2(n20298), .QN(m7_data_o[3]) );
  OA22X1 U23250 ( .IN1(n20727), .IN2(n20638), .IN3(n21244), .IN4(n20614), .Q(
        n20303) );
  OA22X1 U23251 ( .IN1(n21248), .IN2(n20642), .IN3(n22653), .IN4(n20640), .Q(
        n20302) );
  OA22X1 U23252 ( .IN1(n21256), .IN2(n20628), .IN3(n21245), .IN4(n20630), .Q(
        n20301) );
  NAND2X0 U23253 ( .IN1(m0s4_data_i[4]), .IN2(n29380), .QN(n20300) );
  NAND4X0 U23254 ( .IN1(n20303), .IN2(n20302), .IN3(n20301), .IN4(n20300), 
        .QN(n20309) );
  OA22X1 U23255 ( .IN1(n22654), .IN2(n20643), .IN3(n21246), .IN4(n20639), .Q(
        n20307) );
  OA22X1 U23256 ( .IN1(n21257), .IN2(n20636), .IN3(n21247), .IN4(n20629), .Q(
        n20306) );
  OA22X1 U23257 ( .IN1(n22652), .IN2(n20641), .IN3(n21254), .IN4(n20553), .Q(
        n20305) );
  OA22X1 U23258 ( .IN1(n21253), .IN2(n20631), .IN3(n21255), .IN4(n20627), .Q(
        n20304) );
  NAND4X0 U23259 ( .IN1(n20307), .IN2(n20306), .IN3(n20305), .IN4(n20304), 
        .QN(n20308) );
  NOR2X0 U23260 ( .IN1(n20309), .IN2(n20308), .QN(n20311) );
  NAND2X0 U23261 ( .IN1(n29369), .IN2(n22663), .QN(n20310) );
  NAND2X0 U23262 ( .IN1(n20311), .IN2(n20310), .QN(m7_data_o[4]) );
  OA22X1 U23263 ( .IN1(n22669), .IN2(n20641), .IN3(n21268), .IN4(n20627), .Q(
        n20315) );
  OA22X1 U23264 ( .IN1(n22668), .IN2(n20638), .IN3(n21276), .IN4(n20628), .Q(
        n20314) );
  OA22X1 U23265 ( .IN1(n21274), .IN2(n20639), .IN3(n21266), .IN4(n20643), .Q(
        n20313) );
  NAND2X0 U23266 ( .IN1(m0s7_data_i[5]), .IN2(n29377), .QN(n20312) );
  NAND4X0 U23267 ( .IN1(n20315), .IN2(n20314), .IN3(n20313), .IN4(n20312), 
        .QN(n20321) );
  OA22X1 U23268 ( .IN1(n21279), .IN2(n20642), .IN3(n20736), .IN4(n20631), .Q(
        n20319) );
  OA22X1 U23269 ( .IN1(n21278), .IN2(n20630), .IN3(n21277), .IN4(n20553), .Q(
        n20318) );
  OA22X1 U23270 ( .IN1(n21269), .IN2(n20637), .IN3(n21275), .IN4(n20614), .Q(
        n20317) );
  OA22X1 U23271 ( .IN1(n22671), .IN2(n20640), .IN3(n21267), .IN4(n20629), .Q(
        n20316) );
  NAND4X0 U23272 ( .IN1(n20319), .IN2(n20318), .IN3(n20317), .IN4(n20316), 
        .QN(n20320) );
  NOR2X0 U23273 ( .IN1(n20321), .IN2(n20320), .QN(n20323) );
  NAND2X0 U23274 ( .IN1(n29369), .IN2(n22680), .QN(n20322) );
  NAND2X0 U23275 ( .IN1(n20323), .IN2(n20322), .QN(m7_data_o[5]) );
  OA22X1 U23276 ( .IN1(n21298), .IN2(n20642), .IN3(n21290), .IN4(n20637), .Q(
        n20327) );
  OA22X1 U23277 ( .IN1(n21289), .IN2(n20636), .IN3(n22688), .IN4(n20628), .Q(
        n20326) );
  OA22X1 U23278 ( .IN1(n21297), .IN2(n20641), .IN3(n21288), .IN4(n20614), .Q(
        n20325) );
  NAND2X0 U23279 ( .IN1(m0s3_data_i[6]), .IN2(n29381), .QN(n20324) );
  NAND4X0 U23280 ( .IN1(n20327), .IN2(n20326), .IN3(n20325), .IN4(n20324), 
        .QN(n20333) );
  OA22X1 U23281 ( .IN1(n22686), .IN2(n20630), .IN3(n21301), .IN4(n20639), .Q(
        n20331) );
  OA22X1 U23282 ( .IN1(n21300), .IN2(n20629), .IN3(n21299), .IN4(n20553), .Q(
        n20330) );
  OA22X1 U23283 ( .IN1(n21291), .IN2(n20643), .IN3(n22687), .IN4(n20640), .Q(
        n20329) );
  OA22X1 U23284 ( .IN1(n21292), .IN2(n20631), .IN3(n20753), .IN4(n20627), .Q(
        n20328) );
  NAND4X0 U23285 ( .IN1(n20331), .IN2(n20330), .IN3(n20329), .IN4(n20328), 
        .QN(n20332) );
  NOR2X0 U23286 ( .IN1(n20333), .IN2(n20332), .QN(n20335) );
  NAND2X0 U23287 ( .IN1(n29369), .IN2(n22697), .QN(n20334) );
  NAND2X0 U23288 ( .IN1(n20335), .IN2(n20334), .QN(m7_data_o[6]) );
  OA22X1 U23289 ( .IN1(n22703), .IN2(n20553), .IN3(n21313), .IN4(n20640), .Q(
        n20339) );
  OA22X1 U23290 ( .IN1(n21312), .IN2(n20631), .IN3(n21321), .IN4(n20642), .Q(
        n20338) );
  OA22X1 U23291 ( .IN1(n22705), .IN2(n20637), .IN3(n20766), .IN4(n20636), .Q(
        n20337) );
  NAND2X0 U23292 ( .IN1(m0s2_data_i[7]), .IN2(n29382), .QN(n20336) );
  NAND4X0 U23293 ( .IN1(n20339), .IN2(n20338), .IN3(n20337), .IN4(n20336), 
        .QN(n20345) );
  OA22X1 U23294 ( .IN1(n21319), .IN2(n20628), .IN3(n21314), .IN4(n20630), .Q(
        n20343) );
  OA22X1 U23295 ( .IN1(n21322), .IN2(n20629), .IN3(n21320), .IN4(n20638), .Q(
        n20342) );
  OA22X1 U23296 ( .IN1(n21323), .IN2(n20614), .IN3(n21310), .IN4(n20627), .Q(
        n20341) );
  OA22X1 U23297 ( .IN1(n22704), .IN2(n20643), .IN3(n21311), .IN4(n20639), .Q(
        n20340) );
  NAND4X0 U23298 ( .IN1(n20343), .IN2(n20342), .IN3(n20341), .IN4(n20340), 
        .QN(n20344) );
  NOR2X0 U23299 ( .IN1(n20345), .IN2(n20344), .QN(n20347) );
  NAND2X0 U23300 ( .IN1(n29369), .IN2(n22714), .QN(n20346) );
  NAND2X0 U23301 ( .IN1(n20347), .IN2(n20346), .QN(m7_data_o[7]) );
  OA22X1 U23302 ( .IN1(n22722), .IN2(n20639), .IN3(n22719), .IN4(n20628), .Q(
        n20351) );
  OA22X1 U23303 ( .IN1(n21335), .IN2(n20637), .IN3(n21336), .IN4(n20641), .Q(
        n20350) );
  OA22X1 U23304 ( .IN1(n21333), .IN2(n20627), .IN3(n21342), .IN4(n20631), .Q(
        n20349) );
  NAND2X0 U23305 ( .IN1(m0s0_data_i[8]), .IN2(n29385), .QN(n20348) );
  NAND4X0 U23306 ( .IN1(n20351), .IN2(n20350), .IN3(n20349), .IN4(n20348), 
        .QN(n20357) );
  OA22X1 U23307 ( .IN1(n22720), .IN2(n20636), .IN3(n21337), .IN4(n20630), .Q(
        n20355) );
  OA22X1 U23308 ( .IN1(n21345), .IN2(n20642), .IN3(n21346), .IN4(n20640), .Q(
        n20354) );
  OA22X1 U23309 ( .IN1(n21344), .IN2(n20643), .IN3(n21334), .IN4(n20638), .Q(
        n20353) );
  OA22X1 U23310 ( .IN1(n21343), .IN2(n20614), .IN3(n21332), .IN4(n20629), .Q(
        n20352) );
  NAND4X0 U23311 ( .IN1(n20355), .IN2(n20354), .IN3(n20353), .IN4(n20352), 
        .QN(n20356) );
  NOR2X0 U23312 ( .IN1(n20357), .IN2(n20356), .QN(n20359) );
  NAND2X0 U23313 ( .IN1(n29369), .IN2(n22731), .QN(n20358) );
  NAND2X0 U23314 ( .IN1(n20359), .IN2(n20358), .QN(m7_data_o[8]) );
  OA22X1 U23315 ( .IN1(n20787), .IN2(n20639), .IN3(n21365), .IN4(n20614), .Q(
        n20363) );
  OA22X1 U23316 ( .IN1(n22984), .IN2(n20629), .IN3(n22736), .IN4(n20636), .Q(
        n20362) );
  INVX0 U23317 ( .INP(m0s13_data_i[9]), .ZN(n21363) );
  OA22X1 U23318 ( .IN1(n22978), .IN2(n20628), .IN3(n21363), .IN4(n20640), .Q(
        n20361) );
  NAND2X0 U23319 ( .IN1(m0s11_data_i[9]), .IN2(n29373), .QN(n20360) );
  NAND4X0 U23320 ( .IN1(n20363), .IN2(n20362), .IN3(n20361), .IN4(n20360), 
        .QN(n20369) );
  OA22X1 U23321 ( .IN1(n22979), .IN2(n20643), .IN3(n21362), .IN4(n20553), .Q(
        n20367) );
  OA22X1 U23322 ( .IN1(n21364), .IN2(n20630), .IN3(n21356), .IN4(n20642), .Q(
        n20366) );
  OA22X1 U23323 ( .IN1(n21357), .IN2(n20641), .IN3(n22983), .IN4(n20631), .Q(
        n20365) );
  OA22X1 U23324 ( .IN1(n22981), .IN2(n20638), .IN3(n22980), .IN4(n20637), .Q(
        n20364) );
  NAND4X0 U23325 ( .IN1(n20367), .IN2(n20366), .IN3(n20365), .IN4(n20364), 
        .QN(n20368) );
  NOR2X0 U23326 ( .IN1(n20369), .IN2(n20368), .QN(n20371) );
  NAND2X0 U23327 ( .IN1(n29369), .IN2(n22993), .QN(n20370) );
  NAND2X0 U23328 ( .IN1(n20371), .IN2(n20370), .QN(m7_data_o[9]) );
  OA22X1 U23329 ( .IN1(n21384), .IN2(n20639), .IN3(n22749), .IN4(n20641), .Q(
        n20375) );
  OA22X1 U23330 ( .IN1(n21385), .IN2(n20629), .IN3(n21376), .IN4(n20631), .Q(
        n20374) );
  OA22X1 U23331 ( .IN1(n21375), .IN2(n20553), .IN3(n22751), .IN4(n20630), .Q(
        n20373) );
  NAND2X0 U23332 ( .IN1(m0s8_data_i[10]), .IN2(n29376), .QN(n20372) );
  NAND4X0 U23333 ( .IN1(n20375), .IN2(n20374), .IN3(n20373), .IN4(n20372), 
        .QN(n20381) );
  OA22X1 U23334 ( .IN1(n21383), .IN2(n20640), .IN3(n22752), .IN4(n20638), .Q(
        n20379) );
  OA22X1 U23335 ( .IN1(n22750), .IN2(n20636), .IN3(n22754), .IN4(n20643), .Q(
        n20378) );
  OA22X1 U23336 ( .IN1(n21374), .IN2(n20642), .IN3(n22753), .IN4(n20637), .Q(
        n20377) );
  OA22X1 U23337 ( .IN1(n21382), .IN2(n20627), .IN3(n22329), .IN4(n20614), .Q(
        n20376) );
  NAND4X0 U23338 ( .IN1(n20379), .IN2(n20378), .IN3(n20377), .IN4(n20376), 
        .QN(n20380) );
  NOR2X0 U23339 ( .IN1(n20381), .IN2(n20380), .QN(n20383) );
  NAND2X0 U23340 ( .IN1(n29369), .IN2(n22763), .QN(n20382) );
  NAND2X0 U23341 ( .IN1(n20383), .IN2(n20382), .QN(m7_data_o[10]) );
  OA22X1 U23342 ( .IN1(n23002), .IN2(n20638), .IN3(n21399), .IN4(n20641), .Q(
        n20387) );
  OA22X1 U23343 ( .IN1(n21397), .IN2(n20643), .IN3(n21405), .IN4(n20636), .Q(
        n20386) );
  OA22X1 U23344 ( .IN1(n23004), .IN2(n20642), .IN3(n21398), .IN4(n20553), .Q(
        n20385) );
  NAND2X0 U23345 ( .IN1(m0s14_data_i[11]), .IN2(n29370), .QN(n20384) );
  NAND4X0 U23346 ( .IN1(n20387), .IN2(n20386), .IN3(n20385), .IN4(n20384), 
        .QN(n20393) );
  OA22X1 U23347 ( .IN1(n21396), .IN2(n20629), .IN3(n23000), .IN4(n20628), .Q(
        n20391) );
  OA22X1 U23348 ( .IN1(n22998), .IN2(n20637), .IN3(n21395), .IN4(n20630), .Q(
        n20390) );
  INVX0 U23349 ( .INP(m0s5_data_i[11]), .ZN(n21394) );
  OA22X1 U23350 ( .IN1(n23001), .IN2(n20627), .IN3(n21394), .IN4(n20631), .Q(
        n20389) );
  OA22X1 U23351 ( .IN1(n21406), .IN2(n20640), .IN3(n21404), .IN4(n20639), .Q(
        n20388) );
  NAND4X0 U23352 ( .IN1(n20391), .IN2(n20390), .IN3(n20389), .IN4(n20388), 
        .QN(n20392) );
  NOR2X0 U23353 ( .IN1(n20393), .IN2(n20392), .QN(n20395) );
  NAND2X0 U23354 ( .IN1(n29369), .IN2(n23013), .QN(n20394) );
  NAND2X0 U23355 ( .IN1(n20395), .IN2(n20394), .QN(m7_data_o[11]) );
  OA22X1 U23356 ( .IN1(n21422), .IN2(n20636), .IN3(n23020), .IN4(n20639), .Q(
        n20399) );
  OA22X1 U23357 ( .IN1(n21423), .IN2(n20630), .IN3(n23026), .IN4(n20641), .Q(
        n20398) );
  OA22X1 U23358 ( .IN1(n23022), .IN2(n20629), .IN3(n23025), .IN4(n20643), .Q(
        n20397) );
  NAND2X0 U23359 ( .IN1(m0s14_data_i[12]), .IN2(n29370), .QN(n20396) );
  NAND4X0 U23360 ( .IN1(n20399), .IN2(n20398), .IN3(n20397), .IN4(n20396), 
        .QN(n20405) );
  INVX0 U23361 ( .INP(m0s5_data_i[12]), .ZN(n21415) );
  OA22X1 U23362 ( .IN1(n21416), .IN2(n20628), .IN3(n21415), .IN4(n20631), .Q(
        n20403) );
  OA22X1 U23363 ( .IN1(n23018), .IN2(n20627), .IN3(n21421), .IN4(n20637), .Q(
        n20402) );
  OA22X1 U23364 ( .IN1(n20824), .IN2(n20642), .IN3(n23023), .IN4(n20638), .Q(
        n20401) );
  OA22X1 U23365 ( .IN1(n23019), .IN2(n20553), .IN3(n22780), .IN4(n20640), .Q(
        n20400) );
  NAND4X0 U23366 ( .IN1(n20403), .IN2(n20402), .IN3(n20401), .IN4(n20400), 
        .QN(n20404) );
  NOR2X0 U23367 ( .IN1(n20405), .IN2(n20404), .QN(n20407) );
  NAND2X0 U23368 ( .IN1(n29369), .IN2(n23034), .QN(n20406) );
  NAND2X0 U23369 ( .IN1(n20407), .IN2(n20406), .QN(m7_data_o[12]) );
  OA22X1 U23370 ( .IN1(n21434), .IN2(n20640), .IN3(n23039), .IN4(n20614), .Q(
        n20411) );
  OA22X1 U23371 ( .IN1(n23042), .IN2(n20553), .IN3(n23040), .IN4(n20641), .Q(
        n20410) );
  OA22X1 U23372 ( .IN1(n21435), .IN2(n20643), .IN3(n21432), .IN4(n20631), .Q(
        n20409) );
  NAND2X0 U23373 ( .IN1(m0s3_data_i[13]), .IN2(n29381), .QN(n20408) );
  NAND4X0 U23374 ( .IN1(n20411), .IN2(n20410), .IN3(n20409), .IN4(n20408), 
        .QN(n20417) );
  OA22X1 U23375 ( .IN1(n21441), .IN2(n20637), .IN3(n23043), .IN4(n20629), .Q(
        n20415) );
  OA22X1 U23376 ( .IN1(n23041), .IN2(n20627), .IN3(n21433), .IN4(n20639), .Q(
        n20414) );
  OA22X1 U23377 ( .IN1(n21436), .IN2(n20642), .IN3(n23044), .IN4(n20630), .Q(
        n20413) );
  INVX0 U23378 ( .INP(m0s8_data_i[13]), .ZN(n21442) );
  OA22X1 U23379 ( .IN1(n21443), .IN2(n20636), .IN3(n21442), .IN4(n20628), .Q(
        n20412) );
  NAND4X0 U23380 ( .IN1(n20415), .IN2(n20414), .IN3(n20413), .IN4(n20412), 
        .QN(n20416) );
  NOR2X0 U23381 ( .IN1(n20417), .IN2(n20416), .QN(n20419) );
  NAND2X0 U23382 ( .IN1(n29369), .IN2(n23053), .QN(n20418) );
  NAND2X0 U23383 ( .IN1(n20419), .IN2(n20418), .QN(m7_data_o[13]) );
  OA22X1 U23384 ( .IN1(n23062), .IN2(n20628), .IN3(n20849), .IN4(n20640), .Q(
        n20423) );
  OA22X1 U23385 ( .IN1(n23061), .IN2(n20639), .IN3(n23064), .IN4(n20637), .Q(
        n20422) );
  OA22X1 U23386 ( .IN1(n23070), .IN2(n20614), .IN3(n23068), .IN4(n20627), .Q(
        n20421) );
  NAND2X0 U23387 ( .IN1(m0s9_data_i[14]), .IN2(n29375), .QN(n20420) );
  NAND4X0 U23388 ( .IN1(n20423), .IN2(n20422), .IN3(n20421), .IN4(n20420), 
        .QN(n20429) );
  OA22X1 U23389 ( .IN1(n23060), .IN2(n20641), .IN3(n21452), .IN4(n20631), .Q(
        n20427) );
  INVX0 U23390 ( .INP(m0s3_data_i[14]), .ZN(n21459) );
  OA22X1 U23391 ( .IN1(n23066), .IN2(n20553), .IN3(n21459), .IN4(n20638), .Q(
        n20426) );
  OA22X1 U23392 ( .IN1(n21461), .IN2(n20630), .IN3(n21457), .IN4(n20636), .Q(
        n20425) );
  OA22X1 U23393 ( .IN1(n21460), .IN2(n20642), .IN3(n21458), .IN4(n20643), .Q(
        n20424) );
  NAND4X0 U23394 ( .IN1(n20427), .IN2(n20426), .IN3(n20425), .IN4(n20424), 
        .QN(n20428) );
  NOR2X0 U23395 ( .IN1(n20429), .IN2(n20428), .QN(n20431) );
  NAND2X0 U23396 ( .IN1(n29369), .IN2(n23078), .QN(n20430) );
  NAND2X0 U23397 ( .IN1(n20431), .IN2(n20430), .QN(m7_data_o[14]) );
  OA22X1 U23398 ( .IN1(n23094), .IN2(n20636), .IN3(n21478), .IN4(n20627), .Q(
        n20435) );
  OA22X1 U23399 ( .IN1(n21481), .IN2(n20614), .IN3(n21471), .IN4(n20629), .Q(
        n20434) );
  OA22X1 U23400 ( .IN1(n21479), .IN2(n20642), .IN3(n20862), .IN4(n20640), .Q(
        n20433) );
  NAND2X0 U23401 ( .IN1(m0s5_data_i[15]), .IN2(n29379), .QN(n20432) );
  NAND4X0 U23402 ( .IN1(n20435), .IN2(n20434), .IN3(n20433), .IN4(n20432), 
        .QN(n20441) );
  OA22X1 U23403 ( .IN1(n23086), .IN2(n20639), .IN3(n23084), .IN4(n20630), .Q(
        n20439) );
  OA22X1 U23404 ( .IN1(n23092), .IN2(n20628), .IN3(n23088), .IN4(n20643), .Q(
        n20438) );
  INVX0 U23405 ( .INP(m0s2_data_i[15]), .ZN(n21470) );
  OA22X1 U23406 ( .IN1(n23090), .IN2(n20638), .IN3(n21470), .IN4(n20641), .Q(
        n20437) );
  OA22X1 U23407 ( .IN1(n21477), .IN2(n20553), .IN3(n21480), .IN4(n20637), .Q(
        n20436) );
  NAND4X0 U23408 ( .IN1(n20439), .IN2(n20438), .IN3(n20437), .IN4(n20436), 
        .QN(n20440) );
  NOR2X0 U23409 ( .IN1(n20441), .IN2(n20440), .QN(n20443) );
  NAND2X0 U23410 ( .IN1(n29369), .IN2(n23103), .QN(n20442) );
  NAND2X0 U23411 ( .IN1(n20443), .IN2(n20442), .QN(m7_data_o[15]) );
  OA22X1 U23412 ( .IN1(n20641), .IN2(n21490), .IN3(n20629), .IN4(n21493), .Q(
        n20447) );
  OA22X1 U23413 ( .IN1(n20639), .IN2(n21503), .IN3(n20642), .IN4(n21502), .Q(
        n20446) );
  OA22X1 U23414 ( .IN1(n20637), .IN2(n21494), .IN3(n20638), .IN4(n21491), .Q(
        n20445) );
  NAND2X0 U23415 ( .IN1(n29385), .IN2(m0s0_data_i[16]), .QN(n20444) );
  NAND4X0 U23416 ( .IN1(n20447), .IN2(n20446), .IN3(n20445), .IN4(n20444), 
        .QN(n20453) );
  OA22X1 U23417 ( .IN1(n20631), .IN2(n22009), .IN3(n20630), .IN4(n21501), .Q(
        n20451) );
  OA22X1 U23418 ( .IN1(n20643), .IN2(n22012), .IN3(n20628), .IN4(n21499), .Q(
        n20450) );
  OA22X1 U23419 ( .IN1(n20640), .IN2(n22010), .IN3(n20614), .IN4(n21492), .Q(
        n20449) );
  OA22X1 U23420 ( .IN1(n20636), .IN2(n21500), .IN3(n20627), .IN4(n22011), .Q(
        n20448) );
  NAND4X0 U23421 ( .IN1(n20451), .IN2(n20450), .IN3(n20449), .IN4(n20448), 
        .QN(n20452) );
  NOR2X0 U23422 ( .IN1(n20453), .IN2(n20452), .QN(n20456) );
  NOR2X0 U23423 ( .IN1(n23501), .IN2(n20454), .QN(n20650) );
  NAND2X0 U23424 ( .IN1(s15_data_i[16]), .IN2(n20650), .QN(n20455) );
  NAND2X0 U23425 ( .IN1(n20456), .IN2(n20455), .QN(m7_data_o[16]) );
  OA22X1 U23426 ( .IN1(n20640), .IN2(n22836), .IN3(n20642), .IN4(n21521), .Q(
        n20460) );
  OA22X1 U23427 ( .IN1(n20629), .IN2(n22835), .IN3(n20614), .IN4(n21519), .Q(
        n20459) );
  OA22X1 U23428 ( .IN1(n20637), .IN2(n22833), .IN3(n20627), .IN4(n22832), .Q(
        n20458) );
  NAND2X0 U23429 ( .IN1(n29381), .IN2(m0s3_data_i[17]), .QN(n20457) );
  NAND4X0 U23430 ( .IN1(n20460), .IN2(n20459), .IN3(n20458), .IN4(n20457), 
        .QN(n20466) );
  OA22X1 U23431 ( .IN1(n20641), .IN2(n21512), .IN3(n20636), .IN4(n22831), .Q(
        n20464) );
  OA22X1 U23432 ( .IN1(n20630), .IN2(n22834), .IN3(n20628), .IN4(n22397), .Q(
        n20463) );
  OA22X1 U23433 ( .IN1(n20553), .IN2(n21520), .IN3(n20643), .IN4(n22837), .Q(
        n20462) );
  OA22X1 U23434 ( .IN1(n20639), .IN2(n21518), .IN3(n20631), .IN4(n21513), .Q(
        n20461) );
  NAND4X0 U23435 ( .IN1(n20464), .IN2(n20463), .IN3(n20462), .IN4(n20461), 
        .QN(n20465) );
  NOR2X0 U23436 ( .IN1(n20466), .IN2(n20465), .QN(n20468) );
  NAND2X0 U23437 ( .IN1(s15_data_i[17]), .IN2(n20650), .QN(n20467) );
  NAND2X0 U23438 ( .IN1(n20468), .IN2(n20467), .QN(m7_data_o[17]) );
  OA22X1 U23439 ( .IN1(n20636), .IN2(n22411), .IN3(n20631), .IN4(n22414), .Q(
        n20472) );
  OA22X1 U23440 ( .IN1(n20628), .IN2(n21531), .IN3(n20642), .IN4(n22412), .Q(
        n20471) );
  OA22X1 U23441 ( .IN1(n20638), .IN2(n22413), .IN3(n20614), .IN4(n20901), .Q(
        n20470) );
  NAND2X0 U23442 ( .IN1(n29382), .IN2(m0s2_data_i[18]), .QN(n20469) );
  NAND4X0 U23443 ( .IN1(n20472), .IN2(n20471), .IN3(n20470), .IN4(n20469), 
        .QN(n20478) );
  OA22X1 U23444 ( .IN1(n20640), .IN2(n21539), .IN3(n20630), .IN4(n21540), .Q(
        n20476) );
  OA22X1 U23445 ( .IN1(n20627), .IN2(n21537), .IN3(n20643), .IN4(n22410), .Q(
        n20475) );
  OA22X1 U23446 ( .IN1(n20553), .IN2(n22415), .IN3(n20629), .IN4(n21530), .Q(
        n20474) );
  OA22X1 U23447 ( .IN1(n20639), .IN2(n22037), .IN3(n20637), .IN4(n21536), .Q(
        n20473) );
  NAND4X0 U23448 ( .IN1(n20476), .IN2(n20475), .IN3(n20474), .IN4(n20473), 
        .QN(n20477) );
  NOR2X0 U23449 ( .IN1(n20478), .IN2(n20477), .QN(n20480) );
  NAND2X0 U23450 ( .IN1(s15_data_i[18]), .IN2(n20650), .QN(n20479) );
  NAND2X0 U23451 ( .IN1(n20480), .IN2(n20479), .QN(m7_data_o[18]) );
  OA22X1 U23452 ( .IN1(n20641), .IN2(n21558), .IN3(n20631), .IN4(n22050), .Q(
        n20484) );
  OA22X1 U23453 ( .IN1(n20640), .IN2(n22430), .IN3(n20627), .IN4(n21549), .Q(
        n20483) );
  OA22X1 U23454 ( .IN1(n20636), .IN2(n22435), .IN3(n20629), .IN4(n22429), .Q(
        n20482) );
  NAND2X0 U23455 ( .IN1(n29374), .IN2(m0s10_data_i[19]), .QN(n20481) );
  NAND4X0 U23456 ( .IN1(n20484), .IN2(n20483), .IN3(n20482), .IN4(n20481), 
        .QN(n20490) );
  OA22X1 U23457 ( .IN1(n20637), .IN2(n21556), .IN3(n20553), .IN4(n22433), .Q(
        n20488) );
  OA22X1 U23458 ( .IN1(n20638), .IN2(n22431), .IN3(n20628), .IN4(n21550), .Q(
        n20487) );
  OA22X1 U23459 ( .IN1(n20639), .IN2(n21557), .IN3(n20642), .IN4(n21551), .Q(
        n20486) );
  OA22X1 U23460 ( .IN1(n20614), .IN2(n22428), .IN3(n20643), .IN4(n22434), .Q(
        n20485) );
  NAND4X0 U23461 ( .IN1(n20488), .IN2(n20487), .IN3(n20486), .IN4(n20485), 
        .QN(n20489) );
  NOR2X0 U23462 ( .IN1(n20490), .IN2(n20489), .QN(n20492) );
  NAND2X0 U23463 ( .IN1(s15_data_i[19]), .IN2(n20650), .QN(n20491) );
  NAND2X0 U23464 ( .IN1(n20492), .IN2(n20491), .QN(m7_data_o[19]) );
  OA22X1 U23465 ( .IN1(n20641), .IN2(n22452), .IN3(n20630), .IN4(n21574), .Q(
        n20496) );
  OA22X1 U23466 ( .IN1(n20638), .IN2(n21568), .IN3(n20628), .IN4(n21573), .Q(
        n20495) );
  OA22X1 U23467 ( .IN1(n20627), .IN2(n22450), .IN3(n20629), .IN4(n22447), .Q(
        n20494) );
  NAND2X0 U23468 ( .IN1(n29380), .IN2(m0s4_data_i[20]), .QN(n20493) );
  NAND4X0 U23469 ( .IN1(n20496), .IN2(n20495), .IN3(n20494), .IN4(n20493), 
        .QN(n20502) );
  OA22X1 U23470 ( .IN1(n20631), .IN2(n22448), .IN3(n20553), .IN4(n22451), .Q(
        n20500) );
  OA22X1 U23471 ( .IN1(n20639), .IN2(n21575), .IN3(n20614), .IN4(n22453), .Q(
        n20499) );
  OA22X1 U23472 ( .IN1(n20640), .IN2(n21567), .IN3(n20636), .IN4(n21576), .Q(
        n20498) );
  OA22X1 U23473 ( .IN1(n20643), .IN2(n22449), .IN3(n20642), .IN4(n22454), .Q(
        n20497) );
  NAND4X0 U23474 ( .IN1(n20500), .IN2(n20499), .IN3(n20498), .IN4(n20497), 
        .QN(n20501) );
  NOR2X0 U23475 ( .IN1(n20502), .IN2(n20501), .QN(n20504) );
  NAND2X0 U23476 ( .IN1(s15_data_i[20]), .IN2(n20650), .QN(n20503) );
  NAND2X0 U23477 ( .IN1(n20504), .IN2(n20503), .QN(m7_data_o[20]) );
  OA22X1 U23478 ( .IN1(n20636), .IN2(n22857), .IN3(n20630), .IN4(n22849), .Q(
        n20508) );
  OA22X1 U23479 ( .IN1(n20553), .IN2(n22853), .IN3(n20642), .IN4(n22855), .Q(
        n20507) );
  OA22X1 U23480 ( .IN1(n20640), .IN2(n21587), .IN3(n20629), .IN4(n21594), .Q(
        n20506) );
  NAND2X0 U23481 ( .IN1(n29376), .IN2(m0s8_data_i[21]), .QN(n20505) );
  NAND4X0 U23482 ( .IN1(n20508), .IN2(n20507), .IN3(n20506), .IN4(n20505), 
        .QN(n20514) );
  OA22X1 U23483 ( .IN1(n20638), .IN2(n21593), .IN3(n20614), .IN4(n21586), .Q(
        n20512) );
  OA22X1 U23484 ( .IN1(n20641), .IN2(n22856), .IN3(n20631), .IN4(n22851), .Q(
        n20511) );
  OA22X1 U23485 ( .IN1(n20639), .IN2(n22466), .IN3(n20643), .IN4(n22852), .Q(
        n20510) );
  OA22X1 U23486 ( .IN1(n20637), .IN2(n22850), .IN3(n20627), .IN4(n20942), .Q(
        n20509) );
  NAND4X0 U23487 ( .IN1(n20512), .IN2(n20511), .IN3(n20510), .IN4(n20509), 
        .QN(n20513) );
  NOR2X0 U23488 ( .IN1(n20514), .IN2(n20513), .QN(n20516) );
  NAND2X0 U23489 ( .IN1(s15_data_i[21]), .IN2(n20650), .QN(n20515) );
  NAND2X0 U23490 ( .IN1(n20516), .IN2(n20515), .QN(m7_data_o[21]) );
  OA22X1 U23491 ( .IN1(n20639), .IN2(n21612), .IN3(n20642), .IN4(n22872), .Q(
        n20520) );
  OA22X1 U23492 ( .IN1(n20641), .IN2(n22870), .IN3(n20628), .IN4(n22873), .Q(
        n20519) );
  OA22X1 U23493 ( .IN1(n20640), .IN2(n21611), .IN3(n20629), .IN4(n21610), .Q(
        n20518) );
  NAND2X0 U23494 ( .IN1(n29377), .IN2(m0s7_data_i[22]), .QN(n20517) );
  NAND4X0 U23495 ( .IN1(n20520), .IN2(n20519), .IN3(n20518), .IN4(n20517), 
        .QN(n20526) );
  OA22X1 U23496 ( .IN1(n20631), .IN2(n21609), .IN3(n20643), .IN4(n22875), .Q(
        n20524) );
  OA22X1 U23497 ( .IN1(n20638), .IN2(n22871), .IN3(n20627), .IN4(n20951), .Q(
        n20523) );
  OA22X1 U23498 ( .IN1(n20553), .IN2(n21604), .IN3(n20614), .IN4(n21603), .Q(
        n20522) );
  OA22X1 U23499 ( .IN1(n20637), .IN2(n22876), .IN3(n20630), .IN4(n22869), .Q(
        n20521) );
  NAND4X0 U23500 ( .IN1(n20524), .IN2(n20523), .IN3(n20522), .IN4(n20521), 
        .QN(n20525) );
  NOR2X0 U23501 ( .IN1(n20526), .IN2(n20525), .QN(n20528) );
  NAND2X0 U23502 ( .IN1(s15_data_i[22]), .IN2(n20650), .QN(n20527) );
  NAND2X0 U23503 ( .IN1(n20528), .IN2(n20527), .QN(m7_data_o[22]) );
  OA22X1 U23504 ( .IN1(n20630), .IN2(n22494), .IN3(n20629), .IN4(n21633), .Q(
        n20532) );
  OA22X1 U23505 ( .IN1(n20638), .IN2(n21631), .IN3(n20643), .IN4(n21622), .Q(
        n20531) );
  OA22X1 U23506 ( .IN1(n20639), .IN2(n22491), .IN3(n20628), .IN4(n22492), .Q(
        n20530) );
  NAND2X0 U23507 ( .IN1(n29382), .IN2(m0s2_data_i[23]), .QN(n20529) );
  NAND4X0 U23508 ( .IN1(n20532), .IN2(n20531), .IN3(n20530), .IN4(n20529), 
        .QN(n20538) );
  OA22X1 U23509 ( .IN1(n20637), .IN2(n20968), .IN3(n20614), .IN4(n21621), .Q(
        n20536) );
  OA22X1 U23510 ( .IN1(n20640), .IN2(n21632), .IN3(n20642), .IN4(n21625), .Q(
        n20535) );
  OA22X1 U23511 ( .IN1(n20627), .IN2(n21630), .IN3(n20631), .IN4(n21624), .Q(
        n20534) );
  OA22X1 U23512 ( .IN1(n20636), .IN2(n22495), .IN3(n20553), .IN4(n21634), .Q(
        n20533) );
  NAND4X0 U23513 ( .IN1(n20536), .IN2(n20535), .IN3(n20534), .IN4(n20533), 
        .QN(n20537) );
  NOR2X0 U23514 ( .IN1(n20538), .IN2(n20537), .QN(n20540) );
  NAND2X0 U23515 ( .IN1(s15_data_i[23]), .IN2(n20650), .QN(n20539) );
  NAND2X0 U23516 ( .IN1(n20540), .IN2(n20539), .QN(m7_data_o[23]) );
  OA22X1 U23517 ( .IN1(n20553), .IN2(n21649), .IN3(n20614), .IN4(n22893), .Q(
        n20544) );
  OA22X1 U23518 ( .IN1(n20636), .IN2(n22891), .IN3(n20629), .IN4(n21650), .Q(
        n20543) );
  OA22X1 U23519 ( .IN1(n20637), .IN2(n21644), .IN3(n20631), .IN4(n22895), .Q(
        n20542) );
  NAND2X0 U23520 ( .IN1(n29373), .IN2(m0s11_data_i[24]), .QN(n20541) );
  NAND4X0 U23521 ( .IN1(n20544), .IN2(n20543), .IN3(n20542), .IN4(n20541), 
        .QN(n20550) );
  OA22X1 U23522 ( .IN1(n20641), .IN2(n22890), .IN3(n20628), .IN4(n21653), .Q(
        n20548) );
  OA22X1 U23523 ( .IN1(n20639), .IN2(n22896), .IN3(n20642), .IN4(n22889), .Q(
        n20547) );
  OA22X1 U23524 ( .IN1(n20638), .IN2(n21643), .IN3(n20643), .IN4(n21652), .Q(
        n20546) );
  OA22X1 U23525 ( .IN1(n20640), .IN2(n22888), .IN3(n20630), .IN4(n22892), .Q(
        n20545) );
  NAND4X0 U23526 ( .IN1(n20548), .IN2(n20547), .IN3(n20546), .IN4(n20545), 
        .QN(n20549) );
  NOR2X0 U23527 ( .IN1(n20550), .IN2(n20549), .QN(n20552) );
  NAND2X0 U23528 ( .IN1(s15_data_i[24]), .IN2(n20650), .QN(n20551) );
  NAND2X0 U23529 ( .IN1(n20552), .IN2(n20551), .QN(m7_data_o[24]) );
  OA22X1 U23530 ( .IN1(n20640), .IN2(n20993), .IN3(n20638), .IN4(n22521), .Q(
        n20557) );
  OA22X1 U23531 ( .IN1(n20553), .IN2(n21664), .IN3(n20643), .IN4(n22522), .Q(
        n20556) );
  OA22X1 U23532 ( .IN1(n20641), .IN2(n21663), .IN3(n20636), .IN4(n21672), .Q(
        n20555) );
  NAND2X0 U23533 ( .IN1(n29370), .IN2(m0s14_data_i[25]), .QN(n20554) );
  NAND4X0 U23534 ( .IN1(n20557), .IN2(n20556), .IN3(n20555), .IN4(n20554), 
        .QN(n20563) );
  OA22X1 U23535 ( .IN1(n20637), .IN2(n21665), .IN3(n20629), .IN4(n22520), .Q(
        n20561) );
  OA22X1 U23536 ( .IN1(n20628), .IN2(n21671), .IN3(n20642), .IN4(n22119), .Q(
        n20560) );
  OA22X1 U23537 ( .IN1(n20639), .IN2(n21662), .IN3(n20627), .IN4(n21670), .Q(
        n20559) );
  OA22X1 U23538 ( .IN1(n20631), .IN2(n22525), .IN3(n20630), .IN4(n22523), .Q(
        n20558) );
  NAND4X0 U23539 ( .IN1(n20561), .IN2(n20560), .IN3(n20559), .IN4(n20558), 
        .QN(n20562) );
  NOR2X0 U23540 ( .IN1(n20563), .IN2(n20562), .QN(n20565) );
  NAND2X0 U23541 ( .IN1(s15_data_i[25]), .IN2(n20650), .QN(n20564) );
  NAND2X0 U23542 ( .IN1(n20565), .IN2(n20564), .QN(m7_data_o[25]) );
  OA22X1 U23543 ( .IN1(n20639), .IN2(n21695), .IN3(n20642), .IN4(n22539), .Q(
        n20569) );
  OA22X1 U23544 ( .IN1(n20636), .IN2(n21683), .IN3(n20643), .IN4(n21686), .Q(
        n20568) );
  OA22X1 U23545 ( .IN1(n20641), .IN2(n21682), .IN3(n20553), .IN4(n21692), .Q(
        n20567) );
  NAND2X0 U23546 ( .IN1(n29371), .IN2(m0s13_data_i[26]), .QN(n20566) );
  NAND4X0 U23547 ( .IN1(n20569), .IN2(n20568), .IN3(n20567), .IN4(n20566), 
        .QN(n20575) );
  OA22X1 U23548 ( .IN1(n20614), .IN2(n21681), .IN3(n20628), .IN4(n22538), .Q(
        n20573) );
  OA22X1 U23549 ( .IN1(n20638), .IN2(n21694), .IN3(n20629), .IN4(n21693), .Q(
        n20572) );
  OA22X1 U23550 ( .IN1(n20637), .IN2(n21685), .IN3(n20627), .IN4(n22541), .Q(
        n20571) );
  OA22X1 U23551 ( .IN1(n20631), .IN2(n21684), .IN3(n20630), .IN4(n22540), .Q(
        n20570) );
  NAND4X0 U23552 ( .IN1(n20573), .IN2(n20572), .IN3(n20571), .IN4(n20570), 
        .QN(n20574) );
  NOR2X0 U23553 ( .IN1(n20575), .IN2(n20574), .QN(n20577) );
  NAND2X0 U23554 ( .IN1(s15_data_i[26]), .IN2(n20650), .QN(n20576) );
  NAND2X0 U23555 ( .IN1(n20577), .IN2(n20576), .QN(m7_data_o[26]) );
  OA22X1 U23556 ( .IN1(n20641), .IN2(n22916), .IN3(n20637), .IN4(n21711), .Q(
        n20581) );
  OA22X1 U23557 ( .IN1(n20636), .IN2(n22908), .IN3(n20642), .IN4(n21715), .Q(
        n20580) );
  OA22X1 U23558 ( .IN1(n20640), .IN2(n22918), .IN3(n20638), .IN4(n22912), .Q(
        n20579) );
  NAND2X0 U23559 ( .IN1(n29379), .IN2(m0s5_data_i[27]), .QN(n20578) );
  NAND4X0 U23560 ( .IN1(n20581), .IN2(n20580), .IN3(n20579), .IN4(n20578), 
        .QN(n20587) );
  OA22X1 U23561 ( .IN1(n20614), .IN2(n21710), .IN3(n20643), .IN4(n22915), .Q(
        n20585) );
  OA22X1 U23562 ( .IN1(n20639), .IN2(n22910), .IN3(n20628), .IN4(n22913), .Q(
        n20584) );
  OA22X1 U23563 ( .IN1(n20630), .IN2(n22911), .IN3(n20629), .IN4(n21714), .Q(
        n20583) );
  OA22X1 U23564 ( .IN1(n20627), .IN2(n21713), .IN3(n20553), .IN4(n21018), .Q(
        n20582) );
  NAND4X0 U23565 ( .IN1(n20585), .IN2(n20584), .IN3(n20583), .IN4(n20582), 
        .QN(n20586) );
  NOR2X0 U23566 ( .IN1(n20587), .IN2(n20586), .QN(n20589) );
  NAND2X0 U23567 ( .IN1(s15_data_i[27]), .IN2(n20650), .QN(n20588) );
  NAND2X0 U23568 ( .IN1(n20589), .IN2(n20588), .QN(m7_data_o[27]) );
  OA22X1 U23569 ( .IN1(n20614), .IN2(n21725), .IN3(n20628), .IN4(n21739), .Q(
        n20593) );
  OA22X1 U23570 ( .IN1(n20630), .IN2(n21729), .IN3(n20643), .IN4(n22935), .Q(
        n20592) );
  OA22X1 U23571 ( .IN1(n20636), .IN2(n21737), .IN3(n20638), .IN4(n21743), .Q(
        n20591) );
  NAND2X0 U23572 ( .IN1(n29383), .IN2(m0s1_data_i[28]), .QN(n20590) );
  NAND4X0 U23573 ( .IN1(n20593), .IN2(n20592), .IN3(n20591), .IN4(n20590), 
        .QN(n20599) );
  OA22X1 U23574 ( .IN1(n20641), .IN2(n21741), .IN3(n20631), .IN4(n22936), .Q(
        n20597) );
  OA22X1 U23575 ( .IN1(n20640), .IN2(n22932), .IN3(n20629), .IN4(n22934), .Q(
        n20596) );
  OA22X1 U23576 ( .IN1(n20637), .IN2(n22938), .IN3(n20553), .IN4(n22568), .Q(
        n20595) );
  OA22X1 U23577 ( .IN1(n20627), .IN2(n22930), .IN3(n20642), .IN4(n22940), .Q(
        n20594) );
  NAND4X0 U23578 ( .IN1(n20597), .IN2(n20596), .IN3(n20595), .IN4(n20594), 
        .QN(n20598) );
  NOR2X0 U23579 ( .IN1(n20599), .IN2(n20598), .QN(n20601) );
  NAND2X0 U23580 ( .IN1(s15_data_i[28]), .IN2(n20650), .QN(n20600) );
  NAND2X0 U23581 ( .IN1(n20601), .IN2(n20600), .QN(m7_data_o[28]) );
  OA22X1 U23582 ( .IN1(n20629), .IN2(n22955), .IN3(n20628), .IN4(n21048), .Q(
        n20605) );
  OA22X1 U23583 ( .IN1(n20638), .IN2(n22953), .IN3(n20630), .IN4(n22961), .Q(
        n20604) );
  OA22X1 U23584 ( .IN1(n20614), .IN2(n21050), .IN3(n20643), .IN4(n22957), .Q(
        n20603) );
  NAND2X0 U23585 ( .IN1(n29373), .IN2(m0s11_data_i[29]), .QN(n20602) );
  NAND4X0 U23586 ( .IN1(n20605), .IN2(n20604), .IN3(n20603), .IN4(n20602), 
        .QN(n20611) );
  OA22X1 U23587 ( .IN1(n20640), .IN2(n21041), .IN3(n20553), .IN4(n21043), .Q(
        n20609) );
  OA22X1 U23588 ( .IN1(n20641), .IN2(n21049), .IN3(n20631), .IN4(n21040), .Q(
        n20608) );
  OA22X1 U23589 ( .IN1(n20639), .IN2(n22959), .IN3(n20642), .IN4(n22963), .Q(
        n20607) );
  OA22X1 U23590 ( .IN1(n20637), .IN2(n21051), .IN3(n20636), .IN4(n22583), .Q(
        n20606) );
  NAND4X0 U23591 ( .IN1(n20609), .IN2(n20608), .IN3(n20607), .IN4(n20606), 
        .QN(n20610) );
  NOR2X0 U23592 ( .IN1(n20611), .IN2(n20610), .QN(n20613) );
  NAND2X0 U23593 ( .IN1(s15_data_i[29]), .IN2(n20650), .QN(n20612) );
  NAND2X0 U23594 ( .IN1(n20613), .IN2(n20612), .QN(m7_data_o[29]) );
  OA22X1 U23595 ( .IN1(n20640), .IN2(n22602), .IN3(n20614), .IN4(n22597), .Q(
        n20618) );
  OA22X1 U23596 ( .IN1(n20631), .IN2(n21072), .IN3(n20630), .IN4(n22598), .Q(
        n20617) );
  OA22X1 U23597 ( .IN1(n20641), .IN2(n22603), .IN3(n20628), .IN4(n21061), .Q(
        n20616) );
  NAND2X0 U23598 ( .IN1(n29381), .IN2(m0s3_data_i[30]), .QN(n20615) );
  NAND4X0 U23599 ( .IN1(n20618), .IN2(n20617), .IN3(n20616), .IN4(n20615), 
        .QN(n20624) );
  OA22X1 U23600 ( .IN1(n20636), .IN2(n21060), .IN3(n20629), .IN4(n21067), .Q(
        n20622) );
  OA22X1 U23601 ( .IN1(n20627), .IN2(n21062), .IN3(n20642), .IN4(n21071), .Q(
        n20621) );
  OA22X1 U23602 ( .IN1(n20637), .IN2(n21069), .IN3(n20643), .IN4(n22600), .Q(
        n20620) );
  OA22X1 U23603 ( .IN1(n20639), .IN2(n22601), .IN3(n20553), .IN4(n22177), .Q(
        n20619) );
  NAND4X0 U23604 ( .IN1(n20622), .IN2(n20621), .IN3(n20620), .IN4(n20619), 
        .QN(n20623) );
  NOR2X0 U23605 ( .IN1(n20624), .IN2(n20623), .QN(n20626) );
  NAND2X0 U23606 ( .IN1(s15_data_i[30]), .IN2(n20650), .QN(n20625) );
  NAND2X0 U23607 ( .IN1(n20626), .IN2(n20625), .QN(m7_data_o[30]) );
  OA22X1 U23608 ( .IN1(n20627), .IN2(n21086), .IN3(n20553), .IN4(n21107), .Q(
        n20635) );
  OA22X1 U23609 ( .IN1(n20629), .IN2(n21102), .IN3(n20628), .IN4(n21083), .Q(
        n20634) );
  OA22X1 U23610 ( .IN1(n20631), .IN2(n22616), .IN3(n20630), .IN4(n21088), .Q(
        n20633) );
  NAND2X0 U23611 ( .IN1(n29370), .IN2(m0s14_data_i[31]), .QN(n20632) );
  NAND4X0 U23612 ( .IN1(n20635), .IN2(n20634), .IN3(n20633), .IN4(n20632), 
        .QN(n20649) );
  OA22X1 U23613 ( .IN1(n20637), .IN2(n21105), .IN3(n20636), .IN4(n21090), .Q(
        n20647) );
  OA22X1 U23614 ( .IN1(n20639), .IN2(n21099), .IN3(n20638), .IN4(n22617), .Q(
        n20646) );
  OA22X1 U23615 ( .IN1(n20641), .IN2(n22619), .IN3(n20640), .IN4(n22618), .Q(
        n20645) );
  OA22X1 U23616 ( .IN1(n20643), .IN2(n21097), .IN3(n20642), .IN4(n21081), .Q(
        n20644) );
  NAND4X0 U23617 ( .IN1(n20647), .IN2(n20646), .IN3(n20645), .IN4(n20644), 
        .QN(n20648) );
  NOR2X0 U23618 ( .IN1(n20649), .IN2(n20648), .QN(n20652) );
  NAND2X0 U23619 ( .IN1(s15_data_i[31]), .IN2(n20650), .QN(n20651) );
  NAND2X0 U23620 ( .IN1(n20652), .IN2(n20651), .QN(m7_data_o[31]) );
  INVX0 U23621 ( .INP(m6s0_addr[31]), .ZN(n28956) );
  NOR2X0 U23622 ( .IN1(m6s0_addr[30]), .IN2(n28956), .QN(n20663) );
  NOR2X0 U23623 ( .IN1(m6s0_addr[29]), .IN2(m6s0_addr[28]), .QN(n20662) );
  NAND2X0 U23624 ( .IN1(n20663), .IN2(n20662), .QN(n21084) );
  INVX0 U23625 ( .INP(n21084), .ZN(n29357) );
  AND3X1 U23626 ( .IN1(n23245), .IN2(n23122), .IN3(n23121), .Q(n29109) );
  NAND2X0 U23627 ( .IN1(n29357), .IN2(n29109), .QN(n25675) );
  NOR2X0 U23628 ( .IN1(m6s0_addr[31]), .IN2(m6s0_addr[30]), .QN(n20659) );
  INVX0 U23629 ( .INP(m6s0_addr[29]), .ZN(n28922) );
  NOR2X0 U23630 ( .IN1(m6s0_addr[28]), .IN2(n28922), .QN(n20657) );
  AND2X1 U23631 ( .IN1(n20659), .IN2(n20657), .Q(n29363) );
  NAND3X0 U23632 ( .IN1(n23210), .IN2(n23113), .IN3(n23112), .QN(n27772) );
  NAND2X0 U23633 ( .IN1(n29363), .IN2(n29001), .QN(n27499) );
  OA22X1 U23634 ( .IN1(n23246), .IN2(n25675), .IN3(n23214), .IN4(n27499), .Q(
        n20656) );
  INVX0 U23635 ( .INP(m6s0_addr[30]), .ZN(n28937) );
  NOR2X0 U23636 ( .IN1(n28956), .IN2(n28937), .QN(n20658) );
  AND2X1 U23637 ( .IN1(n20658), .IN2(n20662), .Q(n29353) );
  NAND3X0 U23638 ( .IN1(n23151), .IN2(n23152), .IN3(n23150), .QN(n24738) );
  NAND2X0 U23639 ( .IN1(n29353), .IN2(n29183), .QN(n24453) );
  AND2X1 U23640 ( .IN1(n20662), .IN2(n20659), .Q(n29366) );
  NAND3X0 U23641 ( .IN1(n23155), .IN2(n23156), .IN3(n23154), .QN(n28847) );
  NAND2X0 U23642 ( .IN1(n29366), .IN2(n28966), .QN(n28114) );
  OA22X1 U23643 ( .IN1(n21141), .IN2(n24453), .IN3(n23252), .IN4(n28114), .Q(
        n20655) );
  INVX0 U23644 ( .INP(m6s0_addr[28]), .ZN(n28907) );
  NOR2X0 U23645 ( .IN1(m6s0_addr[29]), .IN2(n28907), .QN(n20660) );
  NAND2X0 U23646 ( .IN1(n20663), .IN2(n20660), .QN(n21103) );
  INVX0 U23647 ( .INP(n21103), .ZN(n29356) );
  AND3X1 U23648 ( .IN1(n23249), .IN2(n23116), .IN3(n23115), .Q(n29138) );
  NAND2X0 U23649 ( .IN1(n29356), .IN2(n29138), .QN(n25374) );
  AND2X1 U23650 ( .IN1(n20663), .IN2(n20657), .Q(n29355) );
  NAND3X0 U23651 ( .IN1(n23159), .IN2(n23160), .IN3(n23158), .QN(n25355) );
  NAND2X0 U23652 ( .IN1(n29355), .IN2(n29145), .QN(n25068) );
  OA22X1 U23653 ( .IN1(n23253), .IN2(n25374), .IN3(n23219), .IN4(n25068), .Q(
        n20654) );
  NOR2X0 U23654 ( .IN1(m6s0_addr[31]), .IN2(n28937), .QN(n20661) );
  NAND2X0 U23655 ( .IN1(n20660), .IN2(n20661), .QN(n21101) );
  INVX0 U23656 ( .INP(n21101), .ZN(n29360) );
  AND3X1 U23657 ( .IN1(n23133), .IN2(n23134), .IN3(n23132), .Q(n29057) );
  NAND2X0 U23658 ( .IN1(n29360), .IN2(n29057), .QN(n26591) );
  OR2X1 U23659 ( .IN1(n21144), .IN2(n26591), .Q(n20653) );
  NAND4X0 U23660 ( .IN1(n20656), .IN2(n20655), .IN3(n20654), .IN4(n20653), 
        .QN(n20670) );
  AND2X1 U23661 ( .IN1(n20661), .IN2(n20657), .Q(n29359) );
  NAND3X0 U23662 ( .IN1(n23138), .IN2(n23137), .IN3(n23136), .QN(n26541) );
  NAND2X0 U23663 ( .IN1(n29359), .IN2(n29074), .QN(n26284) );
  AND2X1 U23664 ( .IN1(n20658), .IN2(n20657), .Q(n29351) );
  NAND3X0 U23665 ( .IN1(n23125), .IN2(n23126), .IN3(n23124), .QN(n24096) );
  NAND2X0 U23666 ( .IN1(n29351), .IN2(n29220), .QN(n23851) );
  OA22X1 U23667 ( .IN1(n21126), .IN2(n26284), .IN3(n21123), .IN4(n23851), .Q(
        n20668) );
  NOR2X0 U23668 ( .IN1(n28922), .IN2(n28907), .QN(n20664) );
  AND2X1 U23669 ( .IN1(n20664), .IN2(n20659), .Q(n29362) );
  NAND3X0 U23670 ( .IN1(n23166), .IN2(n23165), .IN3(n23164), .QN(n27492) );
  NAND2X0 U23671 ( .IN1(n29362), .IN2(n29029), .QN(n27193) );
  NAND2X0 U23672 ( .IN1(n20664), .IN2(n20661), .QN(n21091) );
  INVX0 U23673 ( .INP(n21091), .ZN(n29358) );
  AND3X1 U23674 ( .IN1(n23144), .IN2(n23145), .IN3(n23143), .Q(n29100) );
  NAND2X0 U23675 ( .IN1(n29358), .IN2(n29100), .QN(n25980) );
  OA22X1 U23676 ( .IN1(n21120), .IN2(n27193), .IN3(n23220), .IN4(n25980), .Q(
        n20667) );
  NAND2X0 U23677 ( .IN1(n20658), .IN2(n20660), .QN(n21068) );
  INVX0 U23678 ( .INP(n21068), .ZN(n29352) );
  AND3X1 U23679 ( .IN1(n23130), .IN2(n23129), .IN3(n23128), .Q(n29208) );
  NAND2X0 U23680 ( .IN1(n29352), .IN2(n29208), .QN(n24150) );
  AND2X1 U23681 ( .IN1(n20660), .IN2(n20659), .Q(n29364) );
  NAND3X0 U23682 ( .IN1(n23142), .IN2(n23141), .IN3(n23140), .QN(n28078) );
  NAND2X0 U23683 ( .IN1(n29364), .IN2(n28983), .QN(n27810) );
  OA22X1 U23684 ( .IN1(n23213), .IN2(n24150), .IN3(n21138), .IN4(n27810), .Q(
        n20666) );
  AND2X1 U23685 ( .IN1(n20662), .IN2(n20661), .Q(n29361) );
  NAND3X0 U23686 ( .IN1(n23243), .IN2(n23119), .IN3(n23118), .QN(n27183) );
  NAND2X0 U23687 ( .IN1(n29361), .IN2(n29039), .QN(n26896) );
  NAND2X0 U23688 ( .IN1(n20664), .IN2(n20663), .QN(n21087) );
  INVX0 U23689 ( .INP(n21087), .ZN(n29354) );
  AND3X1 U23690 ( .IN1(n23148), .IN2(n23147), .IN3(n23146), .Q(n29171) );
  NAND2X0 U23691 ( .IN1(n29354), .IN2(n29171), .QN(n24758) );
  OA22X1 U23692 ( .IN1(n23247), .IN2(n26896), .IN3(n21137), .IN4(n24758), .Q(
        n20665) );
  NAND4X0 U23693 ( .IN1(n20668), .IN2(n20667), .IN3(n20666), .IN4(n20665), 
        .QN(n20669) );
  NOR2X0 U23694 ( .IN1(n20670), .IN2(n20669), .QN(n20672) );
  NAND2X0 U23695 ( .IN1(n23389), .IN2(n23261), .QN(n20671) );
  NAND2X0 U23696 ( .IN1(n20672), .IN2(n20671), .QN(m6_ack_o) );
  INVX0 U23697 ( .INP(n29363), .ZN(n21085) );
  OA22X1 U23698 ( .IN1(n22205), .IN2(n21085), .IN3(n21162), .IN4(n21091), .Q(
        n20676) );
  INVX0 U23699 ( .INP(n29355), .ZN(n21089) );
  OA22X1 U23700 ( .IN1(n22207), .IN2(n21089), .IN3(n21159), .IN4(n21103), .Q(
        n20675) );
  INVX0 U23701 ( .INP(n29359), .ZN(n21082) );
  OA22X1 U23702 ( .IN1(n21153), .IN2(n21082), .IN3(n21154), .IN4(n21027), .Q(
        n20674) );
  NAND2X0 U23703 ( .IN1(m0s12_data_i[0]), .IN2(n29353), .QN(n20673) );
  NAND4X0 U23704 ( .IN1(n20676), .IN2(n20675), .IN3(n20674), .IN4(n20673), 
        .QN(n20682) );
  INVX0 U23705 ( .INP(n29366), .ZN(n21108) );
  OA22X1 U23706 ( .IN1(n22204), .IN2(n21108), .IN3(n21160), .IN4(n21101), .Q(
        n20680) );
  OA22X1 U23707 ( .IN1(n22208), .IN2(n21087), .IN3(n21823), .IN4(n21068), .Q(
        n20679) );
  INVX0 U23708 ( .INP(n29364), .ZN(n21100) );
  INVX0 U23709 ( .INP(n29361), .ZN(n21106) );
  OA22X1 U23710 ( .IN1(n21161), .IN2(n21100), .IN3(n22203), .IN4(n21106), .Q(
        n20678) );
  INVX0 U23711 ( .INP(n29362), .ZN(n21104) );
  OA22X1 U23712 ( .IN1(n22206), .IN2(n21104), .IN3(n21163), .IN4(n21084), .Q(
        n20677) );
  NAND4X0 U23713 ( .IN1(n20680), .IN2(n20679), .IN3(n20678), .IN4(n20677), 
        .QN(n20681) );
  NOR2X0 U23714 ( .IN1(n20682), .IN2(n20681), .QN(n20684) );
  INVX0 U23715 ( .INP(n20886), .ZN(n29350) );
  NAND2X0 U23716 ( .IN1(n29350), .IN2(n22218), .QN(n20683) );
  NAND2X0 U23717 ( .IN1(n20684), .IN2(n20683), .QN(m6_data_o[0]) );
  INVX0 U23718 ( .INP(n29353), .ZN(n21098) );
  INVX0 U23719 ( .INP(n29351), .ZN(n21027) );
  OA22X1 U23720 ( .IN1(n21185), .IN2(n21098), .IN3(n22224), .IN4(n21027), .Q(
        n20688) );
  OA22X1 U23721 ( .IN1(n21176), .IN2(n21104), .IN3(n21174), .IN4(n21084), .Q(
        n20687) );
  OA22X1 U23722 ( .IN1(n21184), .IN2(n21068), .IN3(n21175), .IN4(n21082), .Q(
        n20686) );
  NAND2X0 U23723 ( .IN1(m0s4_data_i[1]), .IN2(n29361), .QN(n20685) );
  NAND4X0 U23724 ( .IN1(n20688), .IN2(n20687), .IN3(n20686), .IN4(n20685), 
        .QN(n20695) );
  OA22X1 U23725 ( .IN1(n21182), .IN2(n21100), .IN3(n21186), .IN4(n21089), .Q(
        n20693) );
  OA22X1 U23726 ( .IN1(n21177), .IN2(n21101), .IN3(n22226), .IN4(n21091), .Q(
        n20692) );
  OA22X1 U23727 ( .IN1(n21183), .IN2(n21103), .IN3(n22223), .IN4(n21108), .Q(
        n20691) );
  OA22X1 U23728 ( .IN1(n22225), .IN2(n21085), .IN3(n20689), .IN4(n21087), .Q(
        n20690) );
  NAND4X0 U23729 ( .IN1(n20693), .IN2(n20692), .IN3(n20691), .IN4(n20690), 
        .QN(n20694) );
  NOR2X0 U23730 ( .IN1(n20695), .IN2(n20694), .QN(n20697) );
  NAND2X0 U23731 ( .IN1(n29350), .IN2(n22235), .QN(n20696) );
  NAND2X0 U23732 ( .IN1(n20697), .IN2(n20696), .QN(m6_data_o[1]) );
  OA22X1 U23733 ( .IN1(n21197), .IN2(n21106), .IN3(n21206), .IN4(n21089), .Q(
        n20701) );
  OA22X1 U23734 ( .IN1(n21208), .IN2(n21082), .IN3(n21211), .IN4(n21101), .Q(
        n20700) );
  OA22X1 U23735 ( .IN1(n21210), .IN2(n21103), .IN3(n21196), .IN4(n21084), .Q(
        n20699) );
  NAND2X0 U23736 ( .IN1(m0s12_data_i[2]), .IN2(n29353), .QN(n20698) );
  NAND4X0 U23737 ( .IN1(n20701), .IN2(n20700), .IN3(n20699), .IN4(n20698), 
        .QN(n20708) );
  OA22X1 U23738 ( .IN1(n21209), .IN2(n21091), .IN3(n20702), .IN4(n21087), .Q(
        n20706) );
  OA22X1 U23739 ( .IN1(n21195), .IN2(n21027), .IN3(n21207), .IN4(n21085), .Q(
        n20705) );
  OA22X1 U23740 ( .IN1(n21200), .IN2(n21104), .IN3(n21212), .IN4(n21068), .Q(
        n20704) );
  OA22X1 U23741 ( .IN1(n21205), .IN2(n21108), .IN3(n21199), .IN4(n21100), .Q(
        n20703) );
  NAND4X0 U23742 ( .IN1(n20706), .IN2(n20705), .IN3(n20704), .IN4(n20703), 
        .QN(n20707) );
  NOR2X0 U23743 ( .IN1(n20708), .IN2(n20707), .QN(n20710) );
  NAND2X0 U23744 ( .IN1(n29350), .IN2(n22247), .QN(n20709) );
  NAND2X0 U23745 ( .IN1(n20710), .IN2(n20709), .QN(m6_data_o[2]) );
  OA22X1 U23746 ( .IN1(n21222), .IN2(n21091), .IN3(n22637), .IN4(n21101), .Q(
        n20714) );
  OA22X1 U23747 ( .IN1(n21225), .IN2(n21085), .IN3(n22636), .IN4(n21068), .Q(
        n20713) );
  OA22X1 U23748 ( .IN1(n21224), .IN2(n21082), .IN3(n21232), .IN4(n21089), .Q(
        n20712) );
  NAND2X0 U23749 ( .IN1(m0s14_data_i[3]), .IN2(n29351), .QN(n20711) );
  NAND4X0 U23750 ( .IN1(n20714), .IN2(n20713), .IN3(n20712), .IN4(n20711), 
        .QN(n20720) );
  OA22X1 U23751 ( .IN1(n21221), .IN2(n21104), .IN3(n21233), .IN4(n21084), .Q(
        n20718) );
  OA22X1 U23752 ( .IN1(n21234), .IN2(n21087), .IN3(n22634), .IN4(n21106), .Q(
        n20717) );
  OA22X1 U23753 ( .IN1(n22635), .IN2(n21098), .IN3(n21223), .IN4(n21103), .Q(
        n20716) );
  OA22X1 U23754 ( .IN1(n21226), .IN2(n21100), .IN3(n21235), .IN4(n21108), .Q(
        n20715) );
  NAND4X0 U23755 ( .IN1(n20718), .IN2(n20717), .IN3(n20716), .IN4(n20715), 
        .QN(n20719) );
  NOR2X0 U23756 ( .IN1(n20720), .IN2(n20719), .QN(n20722) );
  NAND2X0 U23757 ( .IN1(n29350), .IN2(n22646), .QN(n20721) );
  NAND2X0 U23758 ( .IN1(n20722), .IN2(n20721), .QN(m6_data_o[3]) );
  OA22X1 U23759 ( .IN1(n22652), .IN2(n21085), .IN3(n21245), .IN4(n21089), .Q(
        n20726) );
  OA22X1 U23760 ( .IN1(n21248), .IN2(n21082), .IN3(n21257), .IN4(n21091), .Q(
        n20725) );
  OA22X1 U23761 ( .IN1(n21256), .IN2(n21084), .IN3(n21244), .IN4(n21027), .Q(
        n20724) );
  NAND2X0 U23762 ( .IN1(m0s11_data_i[4]), .IN2(n29354), .QN(n20723) );
  NAND4X0 U23763 ( .IN1(n20726), .IN2(n20725), .IN3(n20724), .IN4(n20723), 
        .QN(n20733) );
  OA22X1 U23764 ( .IN1(n20727), .IN2(n21104), .IN3(n22654), .IN4(n21098), .Q(
        n20731) );
  OA22X1 U23765 ( .IN1(n21246), .IN2(n21100), .IN3(n22653), .IN4(n21068), .Q(
        n20730) );
  OA22X1 U23766 ( .IN1(n21253), .IN2(n21101), .IN3(n21254), .IN4(n21108), .Q(
        n20729) );
  OA22X1 U23767 ( .IN1(n22651), .IN2(n21106), .IN3(n21247), .IN4(n21103), .Q(
        n20728) );
  NAND4X0 U23768 ( .IN1(n20731), .IN2(n20730), .IN3(n20729), .IN4(n20728), 
        .QN(n20732) );
  NOR2X0 U23769 ( .IN1(n20733), .IN2(n20732), .QN(n20735) );
  NAND2X0 U23770 ( .IN1(n29350), .IN2(n22663), .QN(n20734) );
  NAND2X0 U23771 ( .IN1(n20735), .IN2(n20734), .QN(m6_data_o[4]) );
  OA22X1 U23772 ( .IN1(n20736), .IN2(n21101), .IN3(n22670), .IN4(n21091), .Q(
        n20740) );
  OA22X1 U23773 ( .IN1(n22668), .IN2(n21104), .IN3(n22671), .IN4(n21068), .Q(
        n20739) );
  OA22X1 U23774 ( .IN1(n22669), .IN2(n21085), .IN3(n21276), .IN4(n21084), .Q(
        n20738) );
  NAND2X0 U23775 ( .IN1(m0s12_data_i[5]), .IN2(n29353), .QN(n20737) );
  NAND4X0 U23776 ( .IN1(n20740), .IN2(n20739), .IN3(n20738), .IN4(n20737), 
        .QN(n20746) );
  OA22X1 U23777 ( .IN1(n21279), .IN2(n21082), .IN3(n21269), .IN4(n21106), .Q(
        n20744) );
  OA22X1 U23778 ( .IN1(n21278), .IN2(n21089), .IN3(n21267), .IN4(n21103), .Q(
        n20743) );
  OA22X1 U23779 ( .IN1(n21277), .IN2(n21108), .IN3(n21268), .IN4(n21087), .Q(
        n20742) );
  OA22X1 U23780 ( .IN1(n21275), .IN2(n21027), .IN3(n21274), .IN4(n21100), .Q(
        n20741) );
  NAND4X0 U23781 ( .IN1(n20744), .IN2(n20743), .IN3(n20742), .IN4(n20741), 
        .QN(n20745) );
  NOR2X0 U23782 ( .IN1(n20746), .IN2(n20745), .QN(n20748) );
  NAND2X0 U23783 ( .IN1(n29350), .IN2(n22680), .QN(n20747) );
  NAND2X0 U23784 ( .IN1(n20748), .IN2(n20747), .QN(m6_data_o[5]) );
  OA22X1 U23785 ( .IN1(n21289), .IN2(n21091), .IN3(n21297), .IN4(n21085), .Q(
        n20752) );
  OA22X1 U23786 ( .IN1(n22685), .IN2(n21104), .IN3(n21301), .IN4(n21100), .Q(
        n20751) );
  OA22X1 U23787 ( .IN1(n22686), .IN2(n21089), .IN3(n21300), .IN4(n21103), .Q(
        n20750) );
  NAND2X0 U23788 ( .IN1(m0s8_data_i[6]), .IN2(n29357), .QN(n20749) );
  NAND4X0 U23789 ( .IN1(n20752), .IN2(n20751), .IN3(n20750), .IN4(n20749), 
        .QN(n20759) );
  OA22X1 U23790 ( .IN1(n21292), .IN2(n21101), .IN3(n21298), .IN4(n21082), .Q(
        n20757) );
  OA22X1 U23791 ( .IN1(n21291), .IN2(n21098), .IN3(n21290), .IN4(n21106), .Q(
        n20756) );
  OA22X1 U23792 ( .IN1(n21288), .IN2(n21027), .IN3(n20753), .IN4(n21087), .Q(
        n20755) );
  OA22X1 U23793 ( .IN1(n22687), .IN2(n21068), .IN3(n21299), .IN4(n21108), .Q(
        n20754) );
  NAND4X0 U23794 ( .IN1(n20757), .IN2(n20756), .IN3(n20755), .IN4(n20754), 
        .QN(n20758) );
  NOR2X0 U23795 ( .IN1(n20759), .IN2(n20758), .QN(n20761) );
  NAND2X0 U23796 ( .IN1(n29350), .IN2(n22697), .QN(n20760) );
  NAND2X0 U23797 ( .IN1(n20761), .IN2(n20760), .QN(m6_data_o[6]) );
  OA22X1 U23798 ( .IN1(n21322), .IN2(n21103), .IN3(n21314), .IN4(n21089), .Q(
        n20765) );
  OA22X1 U23799 ( .IN1(n22705), .IN2(n21106), .IN3(n21320), .IN4(n21104), .Q(
        n20764) );
  OA22X1 U23800 ( .IN1(n21311), .IN2(n21100), .IN3(n21323), .IN4(n21027), .Q(
        n20763) );
  NAND2X0 U23801 ( .IN1(m0s8_data_i[7]), .IN2(n29357), .QN(n20762) );
  NAND4X0 U23802 ( .IN1(n20765), .IN2(n20764), .IN3(n20763), .IN4(n20762), 
        .QN(n20772) );
  OA22X1 U23803 ( .IN1(n21321), .IN2(n21082), .IN3(n21313), .IN4(n21068), .Q(
        n20770) );
  OA22X1 U23804 ( .IN1(n21312), .IN2(n21101), .IN3(n22702), .IN4(n21085), .Q(
        n20769) );
  OA22X1 U23805 ( .IN1(n22704), .IN2(n21098), .IN3(n21310), .IN4(n21087), .Q(
        n20768) );
  OA22X1 U23806 ( .IN1(n22703), .IN2(n21108), .IN3(n20766), .IN4(n21091), .Q(
        n20767) );
  NAND4X0 U23807 ( .IN1(n20770), .IN2(n20769), .IN3(n20768), .IN4(n20767), 
        .QN(n20771) );
  NOR2X0 U23808 ( .IN1(n20772), .IN2(n20771), .QN(n20774) );
  NAND2X0 U23809 ( .IN1(n29350), .IN2(n22714), .QN(n20773) );
  NAND2X0 U23810 ( .IN1(n20774), .IN2(n20773), .QN(m6_data_o[7]) );
  OA22X1 U23811 ( .IN1(n21345), .IN2(n21082), .IN3(n22721), .IN4(n21108), .Q(
        n20778) );
  OA22X1 U23812 ( .IN1(n21333), .IN2(n21087), .IN3(n21346), .IN4(n21068), .Q(
        n20777) );
  OA22X1 U23813 ( .IN1(n21344), .IN2(n21098), .IN3(n21336), .IN4(n21085), .Q(
        n20776) );
  NAND2X0 U23814 ( .IN1(m0s3_data_i[8]), .IN2(n29362), .QN(n20775) );
  NAND4X0 U23815 ( .IN1(n20778), .IN2(n20777), .IN3(n20776), .IN4(n20775), 
        .QN(n20784) );
  OA22X1 U23816 ( .IN1(n21337), .IN2(n21089), .IN3(n22719), .IN4(n21084), .Q(
        n20782) );
  OA22X1 U23817 ( .IN1(n21342), .IN2(n21101), .IN3(n22722), .IN4(n21100), .Q(
        n20781) );
  OA22X1 U23818 ( .IN1(n22720), .IN2(n21091), .IN3(n21332), .IN4(n21103), .Q(
        n20780) );
  OA22X1 U23819 ( .IN1(n21335), .IN2(n21106), .IN3(n21343), .IN4(n21027), .Q(
        n20779) );
  NAND4X0 U23820 ( .IN1(n20782), .IN2(n20781), .IN3(n20780), .IN4(n20779), 
        .QN(n20783) );
  NOR2X0 U23821 ( .IN1(n20784), .IN2(n20783), .QN(n20786) );
  NAND2X0 U23822 ( .IN1(n29350), .IN2(n22731), .QN(n20785) );
  NAND2X0 U23823 ( .IN1(n20786), .IN2(n20785), .QN(m6_data_o[8]) );
  OA22X1 U23824 ( .IN1(n21356), .IN2(n21082), .IN3(n22979), .IN4(n21098), .Q(
        n20791) );
  OA22X1 U23825 ( .IN1(n22980), .IN2(n21106), .IN3(n22736), .IN4(n21091), .Q(
        n20790) );
  OA22X1 U23826 ( .IN1(n21357), .IN2(n21085), .IN3(n20787), .IN4(n21100), .Q(
        n20789) );
  NAND2X0 U23827 ( .IN1(m0s14_data_i[9]), .IN2(n29351), .QN(n20788) );
  NAND4X0 U23828 ( .IN1(n20791), .IN2(n20790), .IN3(n20789), .IN4(n20788), 
        .QN(n20797) );
  OA22X1 U23829 ( .IN1(n22984), .IN2(n21103), .IN3(n21363), .IN4(n21068), .Q(
        n20795) );
  OA22X1 U23830 ( .IN1(n21364), .IN2(n21089), .IN3(n21362), .IN4(n21108), .Q(
        n20794) );
  OA22X1 U23831 ( .IN1(n22981), .IN2(n21104), .IN3(n21355), .IN4(n21087), .Q(
        n20793) );
  OA22X1 U23832 ( .IN1(n22978), .IN2(n21084), .IN3(n22983), .IN4(n21101), .Q(
        n20792) );
  NAND4X0 U23833 ( .IN1(n20795), .IN2(n20794), .IN3(n20793), .IN4(n20792), 
        .QN(n20796) );
  NOR2X0 U23834 ( .IN1(n20797), .IN2(n20796), .QN(n20799) );
  NAND2X0 U23835 ( .IN1(n29350), .IN2(n22993), .QN(n20798) );
  NAND2X0 U23836 ( .IN1(n20799), .IN2(n20798), .QN(m6_data_o[9]) );
  OA22X1 U23837 ( .IN1(n21374), .IN2(n21082), .IN3(n21384), .IN4(n21100), .Q(
        n20803) );
  OA22X1 U23838 ( .IN1(n22750), .IN2(n21091), .IN3(n22752), .IN4(n21104), .Q(
        n20802) );
  OA22X1 U23839 ( .IN1(n21383), .IN2(n21068), .IN3(n22749), .IN4(n21085), .Q(
        n20801) );
  NAND2X0 U23840 ( .IN1(m0s4_data_i[10]), .IN2(n29361), .QN(n20800) );
  NAND4X0 U23841 ( .IN1(n20803), .IN2(n20802), .IN3(n20801), .IN4(n20800), 
        .QN(n20809) );
  OA22X1 U23842 ( .IN1(n21385), .IN2(n21103), .IN3(n21377), .IN4(n21084), .Q(
        n20807) );
  OA22X1 U23843 ( .IN1(n21382), .IN2(n21087), .IN3(n22751), .IN4(n21089), .Q(
        n20806) );
  OA22X1 U23844 ( .IN1(n22329), .IN2(n21027), .IN3(n21375), .IN4(n21108), .Q(
        n20805) );
  OA22X1 U23845 ( .IN1(n22754), .IN2(n21098), .IN3(n21376), .IN4(n21101), .Q(
        n20804) );
  NAND4X0 U23846 ( .IN1(n20807), .IN2(n20806), .IN3(n20805), .IN4(n20804), 
        .QN(n20808) );
  NOR2X0 U23847 ( .IN1(n20809), .IN2(n20808), .QN(n20811) );
  NAND2X0 U23848 ( .IN1(n29350), .IN2(n22763), .QN(n20810) );
  NAND2X0 U23849 ( .IN1(n20811), .IN2(n20810), .QN(m6_data_o[10]) );
  OA22X1 U23850 ( .IN1(n23004), .IN2(n21082), .IN3(n21394), .IN4(n21101), .Q(
        n20815) );
  OA22X1 U23851 ( .IN1(n22999), .IN2(n21027), .IN3(n21396), .IN4(n21103), .Q(
        n20814) );
  OA22X1 U23852 ( .IN1(n23001), .IN2(n21087), .IN3(n21395), .IN4(n21089), .Q(
        n20813) );
  NAND2X0 U23853 ( .IN1(m0s12_data_i[11]), .IN2(n29353), .QN(n20812) );
  NAND4X0 U23854 ( .IN1(n20815), .IN2(n20814), .IN3(n20813), .IN4(n20812), 
        .QN(n20821) );
  OA22X1 U23855 ( .IN1(n21406), .IN2(n21068), .IN3(n23002), .IN4(n21104), .Q(
        n20819) );
  OA22X1 U23856 ( .IN1(n21404), .IN2(n21100), .IN3(n23000), .IN4(n21084), .Q(
        n20818) );
  OA22X1 U23857 ( .IN1(n21399), .IN2(n21085), .IN3(n21398), .IN4(n21108), .Q(
        n20817) );
  OA22X1 U23858 ( .IN1(n21405), .IN2(n21091), .IN3(n22998), .IN4(n21106), .Q(
        n20816) );
  NAND4X0 U23859 ( .IN1(n20819), .IN2(n20818), .IN3(n20817), .IN4(n20816), 
        .QN(n20820) );
  NOR2X0 U23860 ( .IN1(n20821), .IN2(n20820), .QN(n20823) );
  NAND2X0 U23861 ( .IN1(n29350), .IN2(n23013), .QN(n20822) );
  NAND2X0 U23862 ( .IN1(n20823), .IN2(n20822), .QN(m6_data_o[11]) );
  OA22X1 U23863 ( .IN1(n23023), .IN2(n21104), .IN3(n21415), .IN4(n21101), .Q(
        n20828) );
  OA22X1 U23864 ( .IN1(n20824), .IN2(n21082), .IN3(n23020), .IN4(n21100), .Q(
        n20827) );
  OA22X1 U23865 ( .IN1(n23024), .IN2(n21027), .IN3(n21421), .IN4(n21106), .Q(
        n20826) );
  NAND2X0 U23866 ( .IN1(m0s10_data_i[12]), .IN2(n29355), .QN(n20825) );
  NAND4X0 U23867 ( .IN1(n20828), .IN2(n20827), .IN3(n20826), .IN4(n20825), 
        .QN(n20834) );
  OA22X1 U23868 ( .IN1(n21416), .IN2(n21084), .IN3(n23022), .IN4(n21103), .Q(
        n20832) );
  OA22X1 U23869 ( .IN1(n23018), .IN2(n21087), .IN3(n22780), .IN4(n21068), .Q(
        n20831) );
  OA22X1 U23870 ( .IN1(n23026), .IN2(n21085), .IN3(n21422), .IN4(n21091), .Q(
        n20830) );
  OA22X1 U23871 ( .IN1(n23019), .IN2(n21108), .IN3(n23025), .IN4(n21098), .Q(
        n20829) );
  NAND4X0 U23872 ( .IN1(n20832), .IN2(n20831), .IN3(n20830), .IN4(n20829), 
        .QN(n20833) );
  NOR2X0 U23873 ( .IN1(n20834), .IN2(n20833), .QN(n20836) );
  NAND2X0 U23874 ( .IN1(n29350), .IN2(n23034), .QN(n20835) );
  NAND2X0 U23875 ( .IN1(n20836), .IN2(n20835), .QN(m6_data_o[12]) );
  OA22X1 U23876 ( .IN1(n21441), .IN2(n21106), .IN3(n23040), .IN4(n21085), .Q(
        n20840) );
  OA22X1 U23877 ( .IN1(n21442), .IN2(n21084), .IN3(n21433), .IN4(n21100), .Q(
        n20839) );
  OA22X1 U23878 ( .IN1(n23044), .IN2(n21089), .IN3(n21435), .IN4(n21098), .Q(
        n20838) );
  NAND2X0 U23879 ( .IN1(m0s13_data_i[13]), .IN2(n29352), .QN(n20837) );
  NAND4X0 U23880 ( .IN1(n20840), .IN2(n20839), .IN3(n20838), .IN4(n20837), 
        .QN(n20846) );
  OA22X1 U23881 ( .IN1(n23042), .IN2(n21108), .IN3(n22793), .IN4(n21104), .Q(
        n20844) );
  OA22X1 U23882 ( .IN1(n21443), .IN2(n21091), .IN3(n23043), .IN4(n21103), .Q(
        n20843) );
  OA22X1 U23883 ( .IN1(n21436), .IN2(n21082), .IN3(n21432), .IN4(n21101), .Q(
        n20842) );
  OA22X1 U23884 ( .IN1(n23041), .IN2(n21087), .IN3(n23039), .IN4(n21027), .Q(
        n20841) );
  NAND4X0 U23885 ( .IN1(n20844), .IN2(n20843), .IN3(n20842), .IN4(n20841), 
        .QN(n20845) );
  NOR2X0 U23886 ( .IN1(n20846), .IN2(n20845), .QN(n20848) );
  NAND2X0 U23887 ( .IN1(n29350), .IN2(n23053), .QN(n20847) );
  NAND2X0 U23888 ( .IN1(n20848), .IN2(n20847), .QN(m6_data_o[13]) );
  OA22X1 U23889 ( .IN1(n23062), .IN2(n21084), .IN3(n23061), .IN4(n21100), .Q(
        n20853) );
  OA22X1 U23890 ( .IN1(n21460), .IN2(n21082), .IN3(n20849), .IN4(n21068), .Q(
        n20852) );
  OA22X1 U23891 ( .IN1(n23060), .IN2(n21085), .IN3(n21457), .IN4(n21091), .Q(
        n20851) );
  NAND2X0 U23892 ( .IN1(m0s9_data_i[14]), .IN2(n29356), .QN(n20850) );
  NAND4X0 U23893 ( .IN1(n20853), .IN2(n20852), .IN3(n20851), .IN4(n20850), 
        .QN(n20859) );
  OA22X1 U23894 ( .IN1(n21459), .IN2(n21104), .IN3(n21452), .IN4(n21101), .Q(
        n20857) );
  OA22X1 U23895 ( .IN1(n23070), .IN2(n21027), .IN3(n21458), .IN4(n21098), .Q(
        n20856) );
  OA22X1 U23896 ( .IN1(n21461), .IN2(n21089), .IN3(n23068), .IN4(n21087), .Q(
        n20855) );
  OA22X1 U23897 ( .IN1(n23066), .IN2(n21108), .IN3(n23064), .IN4(n21106), .Q(
        n20854) );
  NAND4X0 U23898 ( .IN1(n20857), .IN2(n20856), .IN3(n20855), .IN4(n20854), 
        .QN(n20858) );
  NOR2X0 U23899 ( .IN1(n20859), .IN2(n20858), .QN(n20861) );
  NAND2X0 U23900 ( .IN1(n29350), .IN2(n23078), .QN(n20860) );
  NAND2X0 U23901 ( .IN1(n20861), .IN2(n20860), .QN(m6_data_o[14]) );
  OA22X1 U23902 ( .IN1(n23090), .IN2(n21104), .IN3(n21477), .IN4(n21108), .Q(
        n20866) );
  OA22X1 U23903 ( .IN1(n23084), .IN2(n21089), .IN3(n20862), .IN4(n21068), .Q(
        n20865) );
  OA22X1 U23904 ( .IN1(n21481), .IN2(n21027), .IN3(n23088), .IN4(n21098), .Q(
        n20864) );
  NAND2X0 U23905 ( .IN1(m0s8_data_i[15]), .IN2(n29357), .QN(n20863) );
  NAND4X0 U23906 ( .IN1(n20866), .IN2(n20865), .IN3(n20864), .IN4(n20863), 
        .QN(n20872) );
  OA22X1 U23907 ( .IN1(n23094), .IN2(n21091), .IN3(n21471), .IN4(n21103), .Q(
        n20870) );
  OA22X1 U23908 ( .IN1(n23086), .IN2(n21100), .IN3(n21472), .IN4(n21101), .Q(
        n20869) );
  OA22X1 U23909 ( .IN1(n21470), .IN2(n21085), .IN3(n21479), .IN4(n21082), .Q(
        n20868) );
  OA22X1 U23910 ( .IN1(n21478), .IN2(n21087), .IN3(n21480), .IN4(n21106), .Q(
        n20867) );
  NAND4X0 U23911 ( .IN1(n20870), .IN2(n20869), .IN3(n20868), .IN4(n20867), 
        .QN(n20871) );
  NOR2X0 U23912 ( .IN1(n20872), .IN2(n20871), .QN(n20874) );
  NAND2X0 U23913 ( .IN1(n29350), .IN2(n23103), .QN(n20873) );
  NAND2X0 U23914 ( .IN1(n20874), .IN2(n20873), .QN(m6_data_o[15]) );
  OA22X1 U23915 ( .IN1(n21084), .IN2(n21499), .IN3(n21098), .IN4(n22012), .Q(
        n20878) );
  OA22X1 U23916 ( .IN1(n21068), .IN2(n22010), .IN3(n21089), .IN4(n21501), .Q(
        n20877) );
  OA22X1 U23917 ( .IN1(n21103), .IN2(n21493), .IN3(n21082), .IN4(n21502), .Q(
        n20876) );
  NAND2X0 U23918 ( .IN1(n29360), .IN2(m0s5_data_i[16]), .QN(n20875) );
  NAND4X0 U23919 ( .IN1(n20878), .IN2(n20877), .IN3(n20876), .IN4(n20875), 
        .QN(n20885) );
  OA22X1 U23920 ( .IN1(n21100), .IN2(n21503), .IN3(n21027), .IN4(n21492), .Q(
        n20883) );
  OA22X1 U23921 ( .IN1(n21087), .IN2(n22011), .IN3(n21106), .IN4(n21494), .Q(
        n20882) );
  OA22X1 U23922 ( .IN1(n21108), .IN2(n20879), .IN3(n21091), .IN4(n21500), .Q(
        n20881) );
  OA22X1 U23923 ( .IN1(n21104), .IN2(n21491), .IN3(n21085), .IN4(n21490), .Q(
        n20880) );
  NAND4X0 U23924 ( .IN1(n20883), .IN2(n20882), .IN3(n20881), .IN4(n20880), 
        .QN(n20884) );
  NOR2X0 U23925 ( .IN1(n20885), .IN2(n20884), .QN(n20888) );
  NOR2X0 U23926 ( .IN1(n23501), .IN2(n20886), .QN(n21115) );
  NAND2X0 U23927 ( .IN1(s15_data_i[16]), .IN2(n21115), .QN(n20887) );
  NAND2X0 U23928 ( .IN1(n20888), .IN2(n20887), .QN(m6_data_o[16]) );
  OA22X1 U23929 ( .IN1(n21106), .IN2(n22833), .IN3(n21103), .IN4(n22835), .Q(
        n20892) );
  OA22X1 U23930 ( .IN1(n21087), .IN2(n22832), .IN3(n21101), .IN4(n21513), .Q(
        n20891) );
  OA22X1 U23931 ( .IN1(n21104), .IN2(n22830), .IN3(n21089), .IN4(n22834), .Q(
        n20890) );
  NAND2X0 U23932 ( .IN1(n29359), .IN2(m0s6_data_i[17]), .QN(n20889) );
  NAND4X0 U23933 ( .IN1(n20892), .IN2(n20891), .IN3(n20890), .IN4(n20889), 
        .QN(n20898) );
  OA22X1 U23934 ( .IN1(n21100), .IN2(n21518), .IN3(n21091), .IN4(n22831), .Q(
        n20896) );
  OA22X1 U23935 ( .IN1(n21098), .IN2(n22837), .IN3(n21085), .IN4(n21512), .Q(
        n20895) );
  OA22X1 U23936 ( .IN1(n21068), .IN2(n22836), .IN3(n21108), .IN4(n21520), .Q(
        n20894) );
  OA22X1 U23937 ( .IN1(n21084), .IN2(n22397), .IN3(n21027), .IN4(n21519), .Q(
        n20893) );
  NAND4X0 U23938 ( .IN1(n20896), .IN2(n20895), .IN3(n20894), .IN4(n20893), 
        .QN(n20897) );
  NOR2X0 U23939 ( .IN1(n20898), .IN2(n20897), .QN(n20900) );
  NAND2X0 U23940 ( .IN1(s15_data_i[17]), .IN2(n21115), .QN(n20899) );
  NAND2X0 U23941 ( .IN1(n20900), .IN2(n20899), .QN(m6_data_o[17]) );
  OA22X1 U23942 ( .IN1(n21101), .IN2(n22414), .IN3(n21089), .IN4(n21540), .Q(
        n20905) );
  OA22X1 U23943 ( .IN1(n21091), .IN2(n22411), .IN3(n21027), .IN4(n20901), .Q(
        n20904) );
  OA22X1 U23944 ( .IN1(n21108), .IN2(n22415), .IN3(n21082), .IN4(n22412), .Q(
        n20903) );
  NAND2X0 U23945 ( .IN1(n29354), .IN2(m0s11_data_i[18]), .QN(n20902) );
  NAND4X0 U23946 ( .IN1(n20905), .IN2(n20904), .IN3(n20903), .IN4(n20902), 
        .QN(n20911) );
  OA22X1 U23947 ( .IN1(n21068), .IN2(n21539), .IN3(n21103), .IN4(n21530), .Q(
        n20909) );
  OA22X1 U23948 ( .IN1(n21104), .IN2(n22413), .IN3(n21100), .IN4(n22037), .Q(
        n20908) );
  OA22X1 U23949 ( .IN1(n21084), .IN2(n21531), .IN3(n21085), .IN4(n21538), .Q(
        n20907) );
  OA22X1 U23950 ( .IN1(n21106), .IN2(n21536), .IN3(n21098), .IN4(n22410), .Q(
        n20906) );
  NAND4X0 U23951 ( .IN1(n20909), .IN2(n20908), .IN3(n20907), .IN4(n20906), 
        .QN(n20910) );
  NOR2X0 U23952 ( .IN1(n20911), .IN2(n20910), .QN(n20913) );
  NAND2X0 U23953 ( .IN1(s15_data_i[18]), .IN2(n21115), .QN(n20912) );
  NAND2X0 U23954 ( .IN1(n20913), .IN2(n20912), .QN(m6_data_o[18]) );
  OA22X1 U23955 ( .IN1(n21084), .IN2(n21550), .IN3(n21089), .IN4(n22432), .Q(
        n20917) );
  OA22X1 U23956 ( .IN1(n21087), .IN2(n21549), .IN3(n21068), .IN4(n22430), .Q(
        n20916) );
  OA22X1 U23957 ( .IN1(n21100), .IN2(n21557), .IN3(n21091), .IN4(n22435), .Q(
        n20915) );
  NAND2X0 U23958 ( .IN1(n29353), .IN2(m0s12_data_i[19]), .QN(n20914) );
  NAND4X0 U23959 ( .IN1(n20917), .IN2(n20916), .IN3(n20915), .IN4(n20914), 
        .QN(n20923) );
  OA22X1 U23960 ( .IN1(n21108), .IN2(n22433), .IN3(n21106), .IN4(n21556), .Q(
        n20921) );
  OA22X1 U23961 ( .IN1(n21101), .IN2(n22050), .IN3(n21082), .IN4(n21551), .Q(
        n20920) );
  OA22X1 U23962 ( .IN1(n21104), .IN2(n22431), .IN3(n21027), .IN4(n22428), .Q(
        n20919) );
  OA22X1 U23963 ( .IN1(n21085), .IN2(n21558), .IN3(n21103), .IN4(n22429), .Q(
        n20918) );
  NAND4X0 U23964 ( .IN1(n20921), .IN2(n20920), .IN3(n20919), .IN4(n20918), 
        .QN(n20922) );
  NOR2X0 U23965 ( .IN1(n20923), .IN2(n20922), .QN(n20925) );
  NAND2X0 U23966 ( .IN1(s15_data_i[19]), .IN2(n21115), .QN(n20924) );
  NAND2X0 U23967 ( .IN1(n20925), .IN2(n20924), .QN(m6_data_o[19]) );
  OA22X1 U23968 ( .IN1(n21085), .IN2(n22452), .IN3(n21103), .IN4(n22447), .Q(
        n20929) );
  OA22X1 U23969 ( .IN1(n21104), .IN2(n21568), .IN3(n21100), .IN4(n21575), .Q(
        n20928) );
  OA22X1 U23970 ( .IN1(n21091), .IN2(n21576), .IN3(n21089), .IN4(n21574), .Q(
        n20927) );
  NAND2X0 U23971 ( .IN1(n29366), .IN2(m0s0_data_i[20]), .QN(n20926) );
  NAND4X0 U23972 ( .IN1(n20929), .IN2(n20928), .IN3(n20927), .IN4(n20926), 
        .QN(n20935) );
  OA22X1 U23973 ( .IN1(n21101), .IN2(n22448), .IN3(n21098), .IN4(n22449), .Q(
        n20933) );
  OA22X1 U23974 ( .IN1(n21084), .IN2(n21573), .IN3(n21082), .IN4(n22454), .Q(
        n20932) );
  OA22X1 U23975 ( .IN1(n21087), .IN2(n22450), .IN3(n21027), .IN4(n22453), .Q(
        n20931) );
  OA22X1 U23976 ( .IN1(n21068), .IN2(n21567), .IN3(n21106), .IN4(n21577), .Q(
        n20930) );
  NAND4X0 U23977 ( .IN1(n20933), .IN2(n20932), .IN3(n20931), .IN4(n20930), 
        .QN(n20934) );
  NOR2X0 U23978 ( .IN1(n20935), .IN2(n20934), .QN(n20937) );
  NAND2X0 U23979 ( .IN1(s15_data_i[20]), .IN2(n21115), .QN(n20936) );
  NAND2X0 U23980 ( .IN1(n20937), .IN2(n20936), .QN(m6_data_o[20]) );
  OA22X1 U23981 ( .IN1(n21108), .IN2(n22853), .IN3(n21100), .IN4(n22466), .Q(
        n20941) );
  OA22X1 U23982 ( .IN1(n21085), .IN2(n22856), .IN3(n21103), .IN4(n21594), .Q(
        n20940) );
  OA22X1 U23983 ( .IN1(n21084), .IN2(n21592), .IN3(n21106), .IN4(n22850), .Q(
        n20939) );
  NAND2X0 U23984 ( .IN1(n29355), .IN2(m0s10_data_i[21]), .QN(n20938) );
  NAND4X0 U23985 ( .IN1(n20941), .IN2(n20940), .IN3(n20939), .IN4(n20938), 
        .QN(n20948) );
  OA22X1 U23986 ( .IN1(n21101), .IN2(n22851), .IN3(n21104), .IN4(n21593), .Q(
        n20946) );
  OA22X1 U23987 ( .IN1(n21087), .IN2(n20942), .IN3(n21068), .IN4(n21587), .Q(
        n20945) );
  OA22X1 U23988 ( .IN1(n21091), .IN2(n22857), .IN3(n21027), .IN4(n21586), .Q(
        n20944) );
  OA22X1 U23989 ( .IN1(n21098), .IN2(n22852), .IN3(n21082), .IN4(n22855), .Q(
        n20943) );
  NAND4X0 U23990 ( .IN1(n20946), .IN2(n20945), .IN3(n20944), .IN4(n20943), 
        .QN(n20947) );
  NOR2X0 U23991 ( .IN1(n20948), .IN2(n20947), .QN(n20950) );
  NAND2X0 U23992 ( .IN1(s15_data_i[21]), .IN2(n21115), .QN(n20949) );
  NAND2X0 U23993 ( .IN1(n20950), .IN2(n20949), .QN(m6_data_o[21]) );
  OA22X1 U23994 ( .IN1(n21087), .IN2(n20951), .IN3(n21085), .IN4(n22870), .Q(
        n20955) );
  OA22X1 U23995 ( .IN1(n21068), .IN2(n21611), .IN3(n21104), .IN4(n22871), .Q(
        n20954) );
  OA22X1 U23996 ( .IN1(n21098), .IN2(n22875), .IN3(n21089), .IN4(n22869), .Q(
        n20953) );
  NAND2X0 U23997 ( .IN1(n29358), .IN2(m0s7_data_i[22]), .QN(n20952) );
  NAND4X0 U23998 ( .IN1(n20955), .IN2(n20954), .IN3(n20953), .IN4(n20952), 
        .QN(n20961) );
  OA22X1 U23999 ( .IN1(n21103), .IN2(n21610), .IN3(n21082), .IN4(n22872), .Q(
        n20959) );
  OA22X1 U24000 ( .IN1(n21101), .IN2(n21609), .IN3(n21100), .IN4(n21612), .Q(
        n20958) );
  OA22X1 U24001 ( .IN1(n21084), .IN2(n22873), .IN3(n21106), .IN4(n22876), .Q(
        n20957) );
  OA22X1 U24002 ( .IN1(n21108), .IN2(n21604), .IN3(n21027), .IN4(n21603), .Q(
        n20956) );
  NAND4X0 U24003 ( .IN1(n20959), .IN2(n20958), .IN3(n20957), .IN4(n20956), 
        .QN(n20960) );
  NOR2X0 U24004 ( .IN1(n20961), .IN2(n20960), .QN(n20963) );
  NAND2X0 U24005 ( .IN1(s15_data_i[22]), .IN2(n21115), .QN(n20962) );
  NAND2X0 U24006 ( .IN1(n20963), .IN2(n20962), .QN(m6_data_o[22]) );
  OA22X1 U24007 ( .IN1(n21108), .IN2(n21634), .IN3(n21082), .IN4(n21625), .Q(
        n20967) );
  OA22X1 U24008 ( .IN1(n21087), .IN2(n21630), .IN3(n21104), .IN4(n21631), .Q(
        n20966) );
  OA22X1 U24009 ( .IN1(n21084), .IN2(n22492), .IN3(n21085), .IN4(n21623), .Q(
        n20965) );
  NAND2X0 U24010 ( .IN1(n29360), .IN2(m0s5_data_i[23]), .QN(n20964) );
  NAND4X0 U24011 ( .IN1(n20967), .IN2(n20966), .IN3(n20965), .IN4(n20964), 
        .QN(n20974) );
  OA22X1 U24012 ( .IN1(n21100), .IN2(n22491), .IN3(n21089), .IN4(n22494), .Q(
        n20972) );
  OA22X1 U24013 ( .IN1(n21068), .IN2(n21632), .IN3(n21098), .IN4(n21622), .Q(
        n20971) );
  OA22X1 U24014 ( .IN1(n21091), .IN2(n22495), .IN3(n21027), .IN4(n21621), .Q(
        n20970) );
  OA22X1 U24015 ( .IN1(n21106), .IN2(n20968), .IN3(n21103), .IN4(n21633), .Q(
        n20969) );
  NAND4X0 U24016 ( .IN1(n20972), .IN2(n20971), .IN3(n20970), .IN4(n20969), 
        .QN(n20973) );
  NOR2X0 U24017 ( .IN1(n20974), .IN2(n20973), .QN(n20976) );
  NAND2X0 U24018 ( .IN1(s15_data_i[23]), .IN2(n21115), .QN(n20975) );
  NAND2X0 U24019 ( .IN1(n20976), .IN2(n20975), .QN(m6_data_o[23]) );
  OA22X1 U24020 ( .IN1(n21108), .IN2(n21649), .IN3(n21100), .IN4(n22896), .Q(
        n20980) );
  OA22X1 U24021 ( .IN1(n21068), .IN2(n22888), .IN3(n21082), .IN4(n22889), .Q(
        n20979) );
  OA22X1 U24022 ( .IN1(n21085), .IN2(n22890), .IN3(n21089), .IN4(n22892), .Q(
        n20978) );
  NAND2X0 U24023 ( .IN1(n29360), .IN2(m0s5_data_i[24]), .QN(n20977) );
  NAND4X0 U24024 ( .IN1(n20980), .IN2(n20979), .IN3(n20978), .IN4(n20977), 
        .QN(n20986) );
  OA22X1 U24025 ( .IN1(n21084), .IN2(n21653), .IN3(n21103), .IN4(n21650), .Q(
        n20984) );
  OA22X1 U24026 ( .IN1(n21087), .IN2(n21651), .IN3(n21091), .IN4(n22891), .Q(
        n20983) );
  OA22X1 U24027 ( .IN1(n21104), .IN2(n21643), .IN3(n21106), .IN4(n21644), .Q(
        n20982) );
  OA22X1 U24028 ( .IN1(n21098), .IN2(n21652), .IN3(n21027), .IN4(n22893), .Q(
        n20981) );
  NAND4X0 U24029 ( .IN1(n20984), .IN2(n20983), .IN3(n20982), .IN4(n20981), 
        .QN(n20985) );
  NOR2X0 U24030 ( .IN1(n20986), .IN2(n20985), .QN(n20988) );
  NAND2X0 U24031 ( .IN1(s15_data_i[24]), .IN2(n21115), .QN(n20987) );
  NAND2X0 U24032 ( .IN1(n20988), .IN2(n20987), .QN(m6_data_o[24]) );
  OA22X1 U24033 ( .IN1(n21101), .IN2(n22525), .IN3(n21082), .IN4(n22119), .Q(
        n20992) );
  OA22X1 U24034 ( .IN1(n21084), .IN2(n21671), .IN3(n21027), .IN4(n22524), .Q(
        n20991) );
  OA22X1 U24035 ( .IN1(n21106), .IN2(n21665), .IN3(n21098), .IN4(n22522), .Q(
        n20990) );
  NAND2X0 U24036 ( .IN1(n29362), .IN2(m0s3_data_i[25]), .QN(n20989) );
  NAND4X0 U24037 ( .IN1(n20992), .IN2(n20991), .IN3(n20990), .IN4(n20989), 
        .QN(n20999) );
  OA22X1 U24038 ( .IN1(n21068), .IN2(n20993), .IN3(n21103), .IN4(n22520), .Q(
        n20997) );
  OA22X1 U24039 ( .IN1(n21087), .IN2(n21670), .IN3(n21091), .IN4(n21672), .Q(
        n20996) );
  OA22X1 U24040 ( .IN1(n21108), .IN2(n21664), .IN3(n21100), .IN4(n21662), .Q(
        n20995) );
  OA22X1 U24041 ( .IN1(n21085), .IN2(n21663), .IN3(n21089), .IN4(n22523), .Q(
        n20994) );
  NAND4X0 U24042 ( .IN1(n20997), .IN2(n20996), .IN3(n20995), .IN4(n20994), 
        .QN(n20998) );
  NOR2X0 U24043 ( .IN1(n20999), .IN2(n20998), .QN(n21001) );
  NAND2X0 U24044 ( .IN1(s15_data_i[25]), .IN2(n21115), .QN(n21000) );
  NAND2X0 U24045 ( .IN1(n21001), .IN2(n21000), .QN(m6_data_o[25]) );
  OA22X1 U24046 ( .IN1(n21087), .IN2(n22541), .IN3(n21106), .IN4(n21685), .Q(
        n21005) );
  OA22X1 U24047 ( .IN1(n21084), .IN2(n22538), .IN3(n21085), .IN4(n21682), .Q(
        n21004) );
  OA22X1 U24048 ( .IN1(n21098), .IN2(n21686), .IN3(n21082), .IN4(n22539), .Q(
        n21003) );
  NAND2X0 U24049 ( .IN1(n29352), .IN2(m0s13_data_i[26]), .QN(n21002) );
  NAND4X0 U24050 ( .IN1(n21005), .IN2(n21004), .IN3(n21003), .IN4(n21002), 
        .QN(n21011) );
  OA22X1 U24051 ( .IN1(n21100), .IN2(n21695), .IN3(n21103), .IN4(n21693), .Q(
        n21009) );
  OA22X1 U24052 ( .IN1(n21089), .IN2(n22540), .IN3(n21027), .IN4(n21681), .Q(
        n21008) );
  OA22X1 U24053 ( .IN1(n21108), .IN2(n21692), .IN3(n21101), .IN4(n21684), .Q(
        n21007) );
  OA22X1 U24054 ( .IN1(n21104), .IN2(n21694), .IN3(n21091), .IN4(n21683), .Q(
        n21006) );
  NAND4X0 U24055 ( .IN1(n21009), .IN2(n21008), .IN3(n21007), .IN4(n21006), 
        .QN(n21010) );
  NOR2X0 U24056 ( .IN1(n21011), .IN2(n21010), .QN(n21013) );
  NAND2X0 U24057 ( .IN1(s15_data_i[26]), .IN2(n21115), .QN(n21012) );
  NAND2X0 U24058 ( .IN1(n21013), .IN2(n21012), .QN(m6_data_o[26]) );
  OA22X1 U24059 ( .IN1(n21101), .IN2(n21705), .IN3(n21103), .IN4(n21714), .Q(
        n21017) );
  OA22X1 U24060 ( .IN1(n21106), .IN2(n21711), .IN3(n21091), .IN4(n22908), .Q(
        n21016) );
  OA22X1 U24061 ( .IN1(n21068), .IN2(n22918), .IN3(n21082), .IN4(n21715), .Q(
        n21015) );
  NAND2X0 U24062 ( .IN1(n29353), .IN2(m0s12_data_i[27]), .QN(n21014) );
  NAND4X0 U24063 ( .IN1(n21017), .IN2(n21016), .IN3(n21015), .IN4(n21014), 
        .QN(n21024) );
  OA22X1 U24064 ( .IN1(n21100), .IN2(n22910), .IN3(n21027), .IN4(n21710), .Q(
        n21022) );
  OA22X1 U24065 ( .IN1(n21108), .IN2(n21018), .IN3(n21089), .IN4(n22911), .Q(
        n21021) );
  OA22X1 U24066 ( .IN1(n21084), .IN2(n22913), .IN3(n21085), .IN4(n22916), .Q(
        n21020) );
  OA22X1 U24067 ( .IN1(n21087), .IN2(n21713), .IN3(n21104), .IN4(n22912), .Q(
        n21019) );
  NAND4X0 U24068 ( .IN1(n21022), .IN2(n21021), .IN3(n21020), .IN4(n21019), 
        .QN(n21023) );
  NOR2X0 U24069 ( .IN1(n21024), .IN2(n21023), .QN(n21026) );
  NAND2X0 U24070 ( .IN1(s15_data_i[27]), .IN2(n21115), .QN(n21025) );
  NAND2X0 U24071 ( .IN1(n21026), .IN2(n21025), .QN(m6_data_o[27]) );
  OA22X1 U24072 ( .IN1(n21098), .IN2(n22935), .IN3(n21085), .IN4(n21741), .Q(
        n21031) );
  OA22X1 U24073 ( .IN1(n21100), .IN2(n22941), .IN3(n21103), .IN4(n22934), .Q(
        n21030) );
  OA22X1 U24074 ( .IN1(n21027), .IN2(n21725), .IN3(n21082), .IN4(n22940), .Q(
        n21029) );
  NAND2X0 U24075 ( .IN1(n29354), .IN2(m0s11_data_i[28]), .QN(n21028) );
  NAND4X0 U24076 ( .IN1(n21031), .IN2(n21030), .IN3(n21029), .IN4(n21028), 
        .QN(n21037) );
  OA22X1 U24077 ( .IN1(n21108), .IN2(n22568), .IN3(n21091), .IN4(n21737), .Q(
        n21035) );
  OA22X1 U24078 ( .IN1(n21101), .IN2(n22936), .IN3(n21084), .IN4(n21739), .Q(
        n21034) );
  OA22X1 U24079 ( .IN1(n21106), .IN2(n22938), .IN3(n21089), .IN4(n21729), .Q(
        n21033) );
  OA22X1 U24080 ( .IN1(n21068), .IN2(n22932), .IN3(n21104), .IN4(n21743), .Q(
        n21032) );
  NAND4X0 U24081 ( .IN1(n21035), .IN2(n21034), .IN3(n21033), .IN4(n21032), 
        .QN(n21036) );
  NOR2X0 U24082 ( .IN1(n21037), .IN2(n21036), .QN(n21039) );
  NAND2X0 U24083 ( .IN1(s15_data_i[28]), .IN2(n21115), .QN(n21038) );
  NAND2X0 U24084 ( .IN1(n21039), .IN2(n21038), .QN(m6_data_o[28]) );
  OA22X1 U24085 ( .IN1(n21068), .IN2(n21041), .IN3(n21101), .IN4(n21040), .Q(
        n21047) );
  OA22X1 U24086 ( .IN1(n21087), .IN2(n21042), .IN3(n21103), .IN4(n22955), .Q(
        n21046) );
  OA22X1 U24087 ( .IN1(n21108), .IN2(n21043), .IN3(n21091), .IN4(n22583), .Q(
        n21045) );
  NAND2X0 U24088 ( .IN1(n29355), .IN2(m0s10_data_i[29]), .QN(n21044) );
  NAND4X0 U24089 ( .IN1(n21047), .IN2(n21046), .IN3(n21045), .IN4(n21044), 
        .QN(n21057) );
  OA22X1 U24090 ( .IN1(n21104), .IN2(n22953), .IN3(n21098), .IN4(n22957), .Q(
        n21055) );
  OA22X1 U24091 ( .IN1(n21084), .IN2(n21048), .IN3(n21082), .IN4(n22963), .Q(
        n21054) );
  OA22X1 U24092 ( .IN1(n21100), .IN2(n22959), .IN3(n21085), .IN4(n21049), .Q(
        n21053) );
  OA22X1 U24093 ( .IN1(n21106), .IN2(n21051), .IN3(n21027), .IN4(n21050), .Q(
        n21052) );
  NAND4X0 U24094 ( .IN1(n21055), .IN2(n21054), .IN3(n21053), .IN4(n21052), 
        .QN(n21056) );
  NOR2X0 U24095 ( .IN1(n21057), .IN2(n21056), .QN(n21059) );
  NAND2X0 U24096 ( .IN1(s15_data_i[29]), .IN2(n21115), .QN(n21058) );
  NAND2X0 U24097 ( .IN1(n21059), .IN2(n21058), .QN(m6_data_o[29]) );
  OA22X1 U24098 ( .IN1(n21084), .IN2(n21061), .IN3(n21091), .IN4(n21060), .Q(
        n21066) );
  OA22X1 U24099 ( .IN1(n21100), .IN2(n22601), .IN3(n21085), .IN4(n22603), .Q(
        n21065) );
  OA22X1 U24100 ( .IN1(n21087), .IN2(n21062), .IN3(n21108), .IN4(n22177), .Q(
        n21064) );
  NAND2X0 U24101 ( .IN1(n29351), .IN2(m0s14_data_i[30]), .QN(n21063) );
  NAND4X0 U24102 ( .IN1(n21066), .IN2(n21065), .IN3(n21064), .IN4(n21063), 
        .QN(n21078) );
  OA22X1 U24103 ( .IN1(n21068), .IN2(n22602), .IN3(n21103), .IN4(n21067), .Q(
        n21076) );
  OA22X1 U24104 ( .IN1(n21106), .IN2(n21069), .IN3(n21089), .IN4(n22598), .Q(
        n21075) );
  OA22X1 U24105 ( .IN1(n21104), .IN2(n21070), .IN3(n21098), .IN4(n22600), .Q(
        n21074) );
  OA22X1 U24106 ( .IN1(n21101), .IN2(n21072), .IN3(n21082), .IN4(n21071), .Q(
        n21073) );
  NAND4X0 U24107 ( .IN1(n21076), .IN2(n21075), .IN3(n21074), .IN4(n21073), 
        .QN(n21077) );
  NOR2X0 U24108 ( .IN1(n21078), .IN2(n21077), .QN(n21080) );
  NAND2X0 U24109 ( .IN1(s15_data_i[30]), .IN2(n21115), .QN(n21079) );
  NAND2X0 U24110 ( .IN1(n21080), .IN2(n21079), .QN(m6_data_o[30]) );
  OA22X1 U24111 ( .IN1(n21084), .IN2(n21083), .IN3(n21082), .IN4(n21081), .Q(
        n21095) );
  OA22X1 U24112 ( .IN1(n21087), .IN2(n21086), .IN3(n21085), .IN4(n22619), .Q(
        n21094) );
  OA22X1 U24113 ( .IN1(n21091), .IN2(n21090), .IN3(n21089), .IN4(n21088), .Q(
        n21093) );
  NAND2X0 U24114 ( .IN1(n29352), .IN2(m0s13_data_i[31]), .QN(n21092) );
  NAND4X0 U24115 ( .IN1(n21095), .IN2(n21094), .IN3(n21093), .IN4(n21092), 
        .QN(n21114) );
  OA22X1 U24116 ( .IN1(n21098), .IN2(n21097), .IN3(n21027), .IN4(n21096), .Q(
        n21112) );
  OA22X1 U24117 ( .IN1(n21101), .IN2(n22616), .IN3(n21100), .IN4(n21099), .Q(
        n21111) );
  OA22X1 U24118 ( .IN1(n21104), .IN2(n22617), .IN3(n21103), .IN4(n21102), .Q(
        n21110) );
  OA22X1 U24119 ( .IN1(n21108), .IN2(n21107), .IN3(n21106), .IN4(n21105), .Q(
        n21109) );
  NAND4X0 U24120 ( .IN1(n21112), .IN2(n21111), .IN3(n21110), .IN4(n21109), 
        .QN(n21113) );
  NOR2X0 U24121 ( .IN1(n21114), .IN2(n21113), .QN(n21117) );
  NAND2X0 U24122 ( .IN1(s15_data_i[31]), .IN2(n21115), .QN(n21116) );
  NAND2X0 U24123 ( .IN1(n21117), .IN2(n21116), .QN(m6_data_o[31]) );
  NOR3X0 U24124 ( .IN1(n23166), .IN2(n21118), .IN3(n23164), .QN(n29019) );
  NAND2X0 U24125 ( .IN1(n29343), .IN2(n29019), .QN(n27200) );
  INVX0 U24126 ( .INP(n21738), .ZN(n29339) );
  NOR3X0 U24127 ( .IN1(n23145), .IN2(n21119), .IN3(n23143), .QN(n29094) );
  NAND2X0 U24128 ( .IN1(n29339), .IN2(n29094), .QN(n25976) );
  OA22X1 U24129 ( .IN1(n21120), .IN2(n27200), .IN3(n23220), .IN4(n25976), .Q(
        n21132) );
  NAND2X0 U24130 ( .IN1(n23123), .IN2(n21121), .QN(n25967) );
  NAND2X0 U24131 ( .IN1(n29338), .IN2(n29118), .QN(n25677) );
  INVX0 U24132 ( .INP(n21726), .ZN(n29332) );
  NOR3X0 U24133 ( .IN1(n23126), .IN2(n23124), .IN3(n21122), .QN(n29226) );
  NAND2X0 U24134 ( .IN1(n29332), .IN2(n29226), .QN(n23843) );
  OA22X1 U24135 ( .IN1(n23246), .IN2(n25677), .IN3(n21123), .IN4(n23843), .Q(
        n21131) );
  NOR3X0 U24136 ( .IN1(n23243), .IN2(n21124), .IN3(n23118), .QN(n29045) );
  NAND2X0 U24137 ( .IN1(n29342), .IN2(n29045), .QN(n26889) );
  NOR3X0 U24138 ( .IN1(n23138), .IN2(n21125), .IN3(n23136), .QN(n29084) );
  NAND2X0 U24139 ( .IN1(n29340), .IN2(n29084), .QN(n26285) );
  OA22X1 U24140 ( .IN1(n23247), .IN2(n26889), .IN3(n21126), .IN4(n26285), .Q(
        n21130) );
  NOR2X0 U24141 ( .IN1(n21127), .IN2(n23129), .QN(n21128) );
  NAND2X0 U24142 ( .IN1(n23212), .IN2(n21128), .QN(n24418) );
  NAND2X0 U24143 ( .IN1(n29333), .IN2(n29199), .QN(n24148) );
  OR2X1 U24144 ( .IN1(n23213), .IN2(n24148), .Q(n21129) );
  NAND4X0 U24145 ( .IN1(n21132), .IN2(n21131), .IN3(n21130), .IN4(n21129), 
        .QN(n21150) );
  NOR3X0 U24146 ( .IN1(n23210), .IN2(n21133), .IN3(n23113), .QN(n29010) );
  NAND2X0 U24147 ( .IN1(n29344), .IN2(n29010), .QN(n27502) );
  NOR3X0 U24148 ( .IN1(n23160), .IN2(n21134), .IN3(n23158), .QN(n29156) );
  NAND2X0 U24149 ( .IN1(n29336), .IN2(n29156), .QN(n25069) );
  OA22X1 U24150 ( .IN1(n23214), .IN2(n27502), .IN3(n23219), .IN4(n25069), .Q(
        n21148) );
  NOR3X0 U24151 ( .IN1(n23142), .IN2(n23140), .IN3(n21135), .QN(n28991) );
  NAND2X0 U24152 ( .IN1(n29345), .IN2(n28991), .QN(n27803) );
  NOR3X0 U24153 ( .IN1(n23148), .IN2(n23147), .IN3(n21136), .QN(n29173) );
  NAND2X0 U24154 ( .IN1(n29335), .IN2(n29173), .QN(n24764) );
  OA22X1 U24155 ( .IN1(n21138), .IN2(n27803), .IN3(n21137), .IN4(n24764), .Q(
        n21147) );
  NOR3X0 U24156 ( .IN1(n23152), .IN2(n23151), .IN3(n21139), .QN(n29189) );
  NAND2X0 U24157 ( .IN1(n29334), .IN2(n29189), .QN(n24457) );
  NOR3X0 U24158 ( .IN1(n23156), .IN2(n23154), .IN3(n21140), .QN(n28965) );
  NAND2X0 U24159 ( .IN1(n29347), .IN2(n28965), .QN(n28108) );
  OA22X1 U24160 ( .IN1(n21141), .IN2(n24457), .IN3(n23252), .IN4(n28108), .Q(
        n21146) );
  NOR3X0 U24161 ( .IN1(n23249), .IN2(n21142), .IN3(n23116), .QN(n29136) );
  NAND2X0 U24162 ( .IN1(n29337), .IN2(n29136), .QN(n25370) );
  NOR3X0 U24163 ( .IN1(n23134), .IN2(n21143), .IN3(n23132), .QN(n29056) );
  NAND2X0 U24164 ( .IN1(n29341), .IN2(n29056), .QN(n26586) );
  OA22X1 U24165 ( .IN1(n23253), .IN2(n25370), .IN3(n21144), .IN4(n26586), .Q(
        n21145) );
  NAND4X0 U24166 ( .IN1(n21148), .IN2(n21147), .IN3(n21146), .IN4(n21145), 
        .QN(n21149) );
  NOR2X0 U24167 ( .IN1(n21150), .IN2(n21149), .QN(n21152) );
  NAND2X0 U24168 ( .IN1(n23364), .IN2(n23261), .QN(n21151) );
  NAND2X0 U24169 ( .IN1(n21152), .IN2(n21151), .QN(m5_ack_o) );
  OA22X1 U24170 ( .IN1(n21823), .IN2(n21704), .IN3(n22205), .IN4(n21742), .Q(
        n21158) );
  OA22X1 U24171 ( .IN1(n21153), .IN2(n21745), .IN3(n22203), .IN4(n21712), .Q(
        n21157) );
  OA22X1 U24172 ( .IN1(n21154), .IN2(n21726), .IN3(n22204), .IN4(n21724), .Q(
        n21156) );
  NAND2X0 U24173 ( .IN1(m0s12_data_i[0]), .IN2(n29334), .QN(n21155) );
  NAND4X0 U24174 ( .IN1(n21158), .IN2(n21157), .IN3(n21156), .IN4(n21155), 
        .QN(n21169) );
  OA22X1 U24175 ( .IN1(n22207), .IN2(n21730), .IN3(n21159), .IN4(n21746), .Q(
        n21167) );
  OA22X1 U24176 ( .IN1(n21161), .IN2(n21727), .IN3(n21160), .IN4(n21736), .Q(
        n21166) );
  OA22X1 U24177 ( .IN1(n22206), .IN2(n21744), .IN3(n21162), .IN4(n21738), .Q(
        n21165) );
  OA22X1 U24178 ( .IN1(n22208), .IN2(n21728), .IN3(n21163), .IN4(n21740), .Q(
        n21164) );
  NAND4X0 U24179 ( .IN1(n21167), .IN2(n21166), .IN3(n21165), .IN4(n21164), 
        .QN(n21168) );
  NOR2X0 U24180 ( .IN1(n21169), .IN2(n21168), .QN(n21172) );
  INVX0 U24181 ( .INP(n21170), .ZN(n29331) );
  NAND2X0 U24182 ( .IN1(n29331), .IN2(n22218), .QN(n21171) );
  NAND2X0 U24183 ( .IN1(n21172), .IN2(n21171), .QN(m5_data_o[0]) );
  OA22X1 U24184 ( .IN1(n22224), .IN2(n21726), .IN3(n21173), .IN4(n21712), .Q(
        n21181) );
  OA22X1 U24185 ( .IN1(n21175), .IN2(n21745), .IN3(n21174), .IN4(n21740), .Q(
        n21180) );
  OA22X1 U24186 ( .IN1(n21177), .IN2(n21736), .IN3(n21176), .IN4(n21744), .Q(
        n21179) );
  NAND2X0 U24187 ( .IN1(m0s11_data_i[1]), .IN2(n29335), .QN(n21178) );
  NAND4X0 U24188 ( .IN1(n21181), .IN2(n21180), .IN3(n21179), .IN4(n21178), 
        .QN(n21192) );
  OA22X1 U24189 ( .IN1(n22226), .IN2(n21738), .IN3(n21182), .IN4(n21727), .Q(
        n21190) );
  OA22X1 U24190 ( .IN1(n21183), .IN2(n21746), .IN3(n22223), .IN4(n21724), .Q(
        n21189) );
  OA22X1 U24191 ( .IN1(n21185), .IN2(n21735), .IN3(n21184), .IN4(n21704), .Q(
        n21188) );
  OA22X1 U24192 ( .IN1(n22225), .IN2(n21742), .IN3(n21186), .IN4(n21730), .Q(
        n21187) );
  NAND4X0 U24193 ( .IN1(n21190), .IN2(n21189), .IN3(n21188), .IN4(n21187), 
        .QN(n21191) );
  NOR2X0 U24194 ( .IN1(n21192), .IN2(n21191), .QN(n21194) );
  NAND2X0 U24195 ( .IN1(n29331), .IN2(n22235), .QN(n21193) );
  NAND2X0 U24196 ( .IN1(n21194), .IN2(n21193), .QN(m5_data_o[1]) );
  OA22X1 U24197 ( .IN1(n21196), .IN2(n21740), .IN3(n21195), .IN4(n21726), .Q(
        n21204) );
  OA22X1 U24198 ( .IN1(n21198), .IN2(n21735), .IN3(n21197), .IN4(n21712), .Q(
        n21203) );
  OA22X1 U24199 ( .IN1(n21200), .IN2(n21744), .IN3(n21199), .IN4(n21727), .Q(
        n21202) );
  NAND2X0 U24200 ( .IN1(m0s11_data_i[2]), .IN2(n29335), .QN(n21201) );
  NAND4X0 U24201 ( .IN1(n21204), .IN2(n21203), .IN3(n21202), .IN4(n21201), 
        .QN(n21218) );
  OA22X1 U24202 ( .IN1(n21206), .IN2(n21730), .IN3(n21205), .IN4(n21724), .Q(
        n21216) );
  OA22X1 U24203 ( .IN1(n21208), .IN2(n21745), .IN3(n21207), .IN4(n21742), .Q(
        n21215) );
  OA22X1 U24204 ( .IN1(n21210), .IN2(n21746), .IN3(n21209), .IN4(n21738), .Q(
        n21214) );
  OA22X1 U24205 ( .IN1(n21212), .IN2(n21704), .IN3(n21211), .IN4(n21736), .Q(
        n21213) );
  NAND4X0 U24206 ( .IN1(n21216), .IN2(n21215), .IN3(n21214), .IN4(n21213), 
        .QN(n21217) );
  NOR2X0 U24207 ( .IN1(n21218), .IN2(n21217), .QN(n21220) );
  NAND2X0 U24208 ( .IN1(n29331), .IN2(n22247), .QN(n21219) );
  NAND2X0 U24209 ( .IN1(n21220), .IN2(n21219), .QN(m5_data_o[2]) );
  OA22X1 U24210 ( .IN1(n21222), .IN2(n21738), .IN3(n21221), .IN4(n21744), .Q(
        n21230) );
  OA22X1 U24211 ( .IN1(n21224), .IN2(n21745), .IN3(n21223), .IN4(n21746), .Q(
        n21229) );
  OA22X1 U24212 ( .IN1(n21226), .IN2(n21727), .IN3(n21225), .IN4(n21742), .Q(
        n21228) );
  NAND2X0 U24213 ( .IN1(m0s13_data_i[3]), .IN2(n29333), .QN(n21227) );
  NAND4X0 U24214 ( .IN1(n21230), .IN2(n21229), .IN3(n21228), .IN4(n21227), 
        .QN(n21241) );
  OA22X1 U24215 ( .IN1(n22634), .IN2(n21712), .IN3(n21231), .IN4(n21726), .Q(
        n21239) );
  OA22X1 U24216 ( .IN1(n21233), .IN2(n21740), .IN3(n21232), .IN4(n21730), .Q(
        n21238) );
  OA22X1 U24217 ( .IN1(n21234), .IN2(n21728), .IN3(n22637), .IN4(n21736), .Q(
        n21237) );
  OA22X1 U24218 ( .IN1(n22635), .IN2(n21735), .IN3(n21235), .IN4(n21724), .Q(
        n21236) );
  NAND4X0 U24219 ( .IN1(n21239), .IN2(n21238), .IN3(n21237), .IN4(n21236), 
        .QN(n21240) );
  NOR2X0 U24220 ( .IN1(n21241), .IN2(n21240), .QN(n21243) );
  NAND2X0 U24221 ( .IN1(n29331), .IN2(n22646), .QN(n21242) );
  NAND2X0 U24222 ( .IN1(n21243), .IN2(n21242), .QN(m5_data_o[3]) );
  OA22X1 U24223 ( .IN1(n22653), .IN2(n21704), .IN3(n21244), .IN4(n21726), .Q(
        n21252) );
  OA22X1 U24224 ( .IN1(n21246), .IN2(n21727), .IN3(n21245), .IN4(n21730), .Q(
        n21251) );
  OA22X1 U24225 ( .IN1(n21248), .IN2(n21745), .IN3(n21247), .IN4(n21746), .Q(
        n21250) );
  NAND2X0 U24226 ( .IN1(m0s3_data_i[4]), .IN2(n29343), .QN(n21249) );
  NAND4X0 U24227 ( .IN1(n21252), .IN2(n21251), .IN3(n21250), .IN4(n21249), 
        .QN(n21263) );
  OA22X1 U24228 ( .IN1(n21253), .IN2(n21736), .IN3(n22652), .IN4(n21742), .Q(
        n21261) );
  OA22X1 U24229 ( .IN1(n21255), .IN2(n21728), .IN3(n21254), .IN4(n21724), .Q(
        n21260) );
  OA22X1 U24230 ( .IN1(n22651), .IN2(n21712), .IN3(n21256), .IN4(n21740), .Q(
        n21259) );
  OA22X1 U24231 ( .IN1(n22654), .IN2(n21735), .IN3(n21257), .IN4(n21738), .Q(
        n21258) );
  NAND4X0 U24232 ( .IN1(n21261), .IN2(n21260), .IN3(n21259), .IN4(n21258), 
        .QN(n21262) );
  NOR2X0 U24233 ( .IN1(n21263), .IN2(n21262), .QN(n21265) );
  NAND2X0 U24234 ( .IN1(n29331), .IN2(n22663), .QN(n21264) );
  NAND2X0 U24235 ( .IN1(n21265), .IN2(n21264), .QN(m5_data_o[4]) );
  OA22X1 U24236 ( .IN1(n22671), .IN2(n21704), .IN3(n21266), .IN4(n21735), .Q(
        n21273) );
  OA22X1 U24237 ( .IN1(n22668), .IN2(n21744), .IN3(n21267), .IN4(n21746), .Q(
        n21272) );
  OA22X1 U24238 ( .IN1(n21269), .IN2(n21712), .IN3(n21268), .IN4(n21728), .Q(
        n21271) );
  NAND2X0 U24239 ( .IN1(m0s5_data_i[5]), .IN2(n29341), .QN(n21270) );
  NAND4X0 U24240 ( .IN1(n21273), .IN2(n21272), .IN3(n21271), .IN4(n21270), 
        .QN(n21285) );
  OA22X1 U24241 ( .IN1(n22669), .IN2(n21742), .IN3(n21274), .IN4(n21727), .Q(
        n21283) );
  OA22X1 U24242 ( .IN1(n21275), .IN2(n21726), .IN3(n22670), .IN4(n21738), .Q(
        n21282) );
  OA22X1 U24243 ( .IN1(n21277), .IN2(n21724), .IN3(n21276), .IN4(n21740), .Q(
        n21281) );
  OA22X1 U24244 ( .IN1(n21279), .IN2(n21745), .IN3(n21278), .IN4(n21730), .Q(
        n21280) );
  NAND4X0 U24245 ( .IN1(n21283), .IN2(n21282), .IN3(n21281), .IN4(n21280), 
        .QN(n21284) );
  NOR2X0 U24246 ( .IN1(n21285), .IN2(n21284), .QN(n21287) );
  NAND2X0 U24247 ( .IN1(n29331), .IN2(n22680), .QN(n21286) );
  NAND2X0 U24248 ( .IN1(n21287), .IN2(n21286), .QN(m5_data_o[5]) );
  OA22X1 U24249 ( .IN1(n21289), .IN2(n21738), .IN3(n21288), .IN4(n21726), .Q(
        n21296) );
  OA22X1 U24250 ( .IN1(n21291), .IN2(n21735), .IN3(n21290), .IN4(n21712), .Q(
        n21295) );
  OA22X1 U24251 ( .IN1(n21292), .IN2(n21736), .IN3(n22688), .IN4(n21740), .Q(
        n21294) );
  NAND2X0 U24252 ( .IN1(m0s11_data_i[6]), .IN2(n29335), .QN(n21293) );
  NAND4X0 U24253 ( .IN1(n21296), .IN2(n21295), .IN3(n21294), .IN4(n21293), 
        .QN(n21307) );
  OA22X1 U24254 ( .IN1(n21297), .IN2(n21742), .IN3(n22687), .IN4(n21704), .Q(
        n21305) );
  OA22X1 U24255 ( .IN1(n22686), .IN2(n21730), .IN3(n21298), .IN4(n21745), .Q(
        n21304) );
  OA22X1 U24256 ( .IN1(n21300), .IN2(n21746), .IN3(n21299), .IN4(n21724), .Q(
        n21303) );
  OA22X1 U24257 ( .IN1(n22685), .IN2(n21744), .IN3(n21301), .IN4(n21727), .Q(
        n21302) );
  NAND4X0 U24258 ( .IN1(n21305), .IN2(n21304), .IN3(n21303), .IN4(n21302), 
        .QN(n21306) );
  NOR2X0 U24259 ( .IN1(n21307), .IN2(n21306), .QN(n21309) );
  NAND2X0 U24260 ( .IN1(n29331), .IN2(n22697), .QN(n21308) );
  NAND2X0 U24261 ( .IN1(n21309), .IN2(n21308), .QN(m5_data_o[6]) );
  OA22X1 U24262 ( .IN1(n21311), .IN2(n21727), .IN3(n21310), .IN4(n21728), .Q(
        n21318) );
  OA22X1 U24263 ( .IN1(n21312), .IN2(n21736), .IN3(n22702), .IN4(n21742), .Q(
        n21317) );
  OA22X1 U24264 ( .IN1(n21314), .IN2(n21730), .IN3(n21313), .IN4(n21704), .Q(
        n21316) );
  NAND2X0 U24265 ( .IN1(m0s7_data_i[7]), .IN2(n29339), .QN(n21315) );
  NAND4X0 U24266 ( .IN1(n21318), .IN2(n21317), .IN3(n21316), .IN4(n21315), 
        .QN(n21329) );
  OA22X1 U24267 ( .IN1(n22704), .IN2(n21735), .IN3(n21319), .IN4(n21740), .Q(
        n21327) );
  OA22X1 U24268 ( .IN1(n21321), .IN2(n21745), .IN3(n21320), .IN4(n21744), .Q(
        n21326) );
  OA22X1 U24269 ( .IN1(n21322), .IN2(n21746), .IN3(n22703), .IN4(n21724), .Q(
        n21325) );
  OA22X1 U24270 ( .IN1(n22705), .IN2(n21712), .IN3(n21323), .IN4(n21726), .Q(
        n21324) );
  NAND4X0 U24271 ( .IN1(n21327), .IN2(n21326), .IN3(n21325), .IN4(n21324), 
        .QN(n21328) );
  NOR2X0 U24272 ( .IN1(n21329), .IN2(n21328), .QN(n21331) );
  NAND2X0 U24273 ( .IN1(n29331), .IN2(n22714), .QN(n21330) );
  NAND2X0 U24274 ( .IN1(n21331), .IN2(n21330), .QN(m5_data_o[7]) );
  OA22X1 U24275 ( .IN1(n21333), .IN2(n21728), .IN3(n21332), .IN4(n21746), .Q(
        n21341) );
  OA22X1 U24276 ( .IN1(n21335), .IN2(n21712), .IN3(n21334), .IN4(n21744), .Q(
        n21340) );
  OA22X1 U24277 ( .IN1(n21337), .IN2(n21730), .IN3(n21336), .IN4(n21742), .Q(
        n21339) );
  NAND2X0 U24278 ( .IN1(m0s8_data_i[8]), .IN2(n29338), .QN(n21338) );
  NAND4X0 U24279 ( .IN1(n21341), .IN2(n21340), .IN3(n21339), .IN4(n21338), 
        .QN(n21352) );
  OA22X1 U24280 ( .IN1(n21342), .IN2(n21736), .IN3(n22720), .IN4(n21738), .Q(
        n21350) );
  OA22X1 U24281 ( .IN1(n21344), .IN2(n21735), .IN3(n21343), .IN4(n21726), .Q(
        n21349) );
  OA22X1 U24282 ( .IN1(n22722), .IN2(n21727), .IN3(n21345), .IN4(n21745), .Q(
        n21348) );
  OA22X1 U24283 ( .IN1(n22721), .IN2(n21724), .IN3(n21346), .IN4(n21704), .Q(
        n21347) );
  NAND4X0 U24284 ( .IN1(n21350), .IN2(n21349), .IN3(n21348), .IN4(n21347), 
        .QN(n21351) );
  NOR2X0 U24285 ( .IN1(n21352), .IN2(n21351), .QN(n21354) );
  NAND2X0 U24286 ( .IN1(n29331), .IN2(n22731), .QN(n21353) );
  NAND2X0 U24287 ( .IN1(n21354), .IN2(n21353), .QN(m5_data_o[8]) );
  OA22X1 U24288 ( .IN1(n21355), .IN2(n21728), .IN3(n22980), .IN4(n21712), .Q(
        n21361) );
  OA22X1 U24289 ( .IN1(n22984), .IN2(n21746), .IN3(n21356), .IN4(n21745), .Q(
        n21360) );
  OA22X1 U24290 ( .IN1(n21357), .IN2(n21742), .IN3(n22979), .IN4(n21735), .Q(
        n21359) );
  NAND2X0 U24291 ( .IN1(m0s1_data_i[9]), .IN2(n29345), .QN(n21358) );
  NAND4X0 U24292 ( .IN1(n21361), .IN2(n21360), .IN3(n21359), .IN4(n21358), 
        .QN(n21371) );
  OA22X1 U24293 ( .IN1(n21363), .IN2(n21704), .IN3(n21362), .IN4(n21724), .Q(
        n21369) );
  OA22X1 U24294 ( .IN1(n21364), .IN2(n21730), .IN3(n22983), .IN4(n21736), .Q(
        n21368) );
  OA22X1 U24295 ( .IN1(n22978), .IN2(n21740), .IN3(n21365), .IN4(n21726), .Q(
        n21367) );
  OA22X1 U24296 ( .IN1(n22981), .IN2(n21744), .IN3(n22736), .IN4(n21738), .Q(
        n21366) );
  NAND4X0 U24297 ( .IN1(n21369), .IN2(n21368), .IN3(n21367), .IN4(n21366), 
        .QN(n21370) );
  NOR2X0 U24298 ( .IN1(n21371), .IN2(n21370), .QN(n21373) );
  NAND2X0 U24299 ( .IN1(n29331), .IN2(n22993), .QN(n21372) );
  NAND2X0 U24300 ( .IN1(n21373), .IN2(n21372), .QN(m5_data_o[9]) );
  OA22X1 U24301 ( .IN1(n21374), .IN2(n21745), .IN3(n22753), .IN4(n21712), .Q(
        n21381) );
  OA22X1 U24302 ( .IN1(n22752), .IN2(n21744), .IN3(n21375), .IN4(n21724), .Q(
        n21380) );
  OA22X1 U24303 ( .IN1(n21377), .IN2(n21740), .IN3(n21376), .IN4(n21736), .Q(
        n21379) );
  NAND2X0 U24304 ( .IN1(m0s7_data_i[10]), .IN2(n29339), .QN(n21378) );
  NAND4X0 U24305 ( .IN1(n21381), .IN2(n21380), .IN3(n21379), .IN4(n21378), 
        .QN(n21391) );
  OA22X1 U24306 ( .IN1(n21383), .IN2(n21704), .IN3(n21382), .IN4(n21728), .Q(
        n21389) );
  OA22X1 U24307 ( .IN1(n22754), .IN2(n21735), .IN3(n22751), .IN4(n21730), .Q(
        n21388) );
  OA22X1 U24308 ( .IN1(n21385), .IN2(n21746), .IN3(n21384), .IN4(n21727), .Q(
        n21387) );
  OA22X1 U24309 ( .IN1(n22329), .IN2(n21726), .IN3(n22749), .IN4(n21742), .Q(
        n21386) );
  NAND4X0 U24310 ( .IN1(n21389), .IN2(n21388), .IN3(n21387), .IN4(n21386), 
        .QN(n21390) );
  NOR2X0 U24311 ( .IN1(n21391), .IN2(n21390), .QN(n21393) );
  NAND2X0 U24312 ( .IN1(n29331), .IN2(n22763), .QN(n21392) );
  NAND2X0 U24313 ( .IN1(n21393), .IN2(n21392), .QN(m5_data_o[10]) );
  OA22X1 U24314 ( .IN1(n21395), .IN2(n21730), .IN3(n21394), .IN4(n21736), .Q(
        n21403) );
  OA22X1 U24315 ( .IN1(n21397), .IN2(n21735), .IN3(n21396), .IN4(n21746), .Q(
        n21402) );
  OA22X1 U24316 ( .IN1(n21399), .IN2(n21742), .IN3(n21398), .IN4(n21724), .Q(
        n21401) );
  NAND2X0 U24317 ( .IN1(m0s8_data_i[11]), .IN2(n29338), .QN(n21400) );
  NAND4X0 U24318 ( .IN1(n21403), .IN2(n21402), .IN3(n21401), .IN4(n21400), 
        .QN(n21412) );
  OA22X1 U24319 ( .IN1(n23004), .IN2(n21745), .IN3(n21404), .IN4(n21727), .Q(
        n21410) );
  OA22X1 U24320 ( .IN1(n21405), .IN2(n21738), .IN3(n22998), .IN4(n21712), .Q(
        n21409) );
  OA22X1 U24321 ( .IN1(n21406), .IN2(n21704), .IN3(n23001), .IN4(n21728), .Q(
        n21408) );
  OA22X1 U24322 ( .IN1(n22999), .IN2(n21726), .IN3(n23002), .IN4(n21744), .Q(
        n21407) );
  NAND4X0 U24323 ( .IN1(n21410), .IN2(n21409), .IN3(n21408), .IN4(n21407), 
        .QN(n21411) );
  NOR2X0 U24324 ( .IN1(n21412), .IN2(n21411), .QN(n21414) );
  NAND2X0 U24325 ( .IN1(n29331), .IN2(n23013), .QN(n21413) );
  NAND2X0 U24326 ( .IN1(n21414), .IN2(n21413), .QN(m5_data_o[11]) );
  OA22X1 U24327 ( .IN1(n21416), .IN2(n21740), .IN3(n21415), .IN4(n21736), .Q(
        n21420) );
  OA22X1 U24328 ( .IN1(n23025), .IN2(n21735), .IN3(n23023), .IN4(n21744), .Q(
        n21419) );
  OA22X1 U24329 ( .IN1(n23026), .IN2(n21742), .IN3(n23020), .IN4(n21727), .Q(
        n21418) );
  NAND2X0 U24330 ( .IN1(m0s6_data_i[12]), .IN2(n29340), .QN(n21417) );
  NAND4X0 U24331 ( .IN1(n21420), .IN2(n21419), .IN3(n21418), .IN4(n21417), 
        .QN(n21429) );
  OA22X1 U24332 ( .IN1(n21421), .IN2(n21712), .IN3(n22780), .IN4(n21704), .Q(
        n21427) );
  OA22X1 U24333 ( .IN1(n21423), .IN2(n21730), .IN3(n21422), .IN4(n21738), .Q(
        n21426) );
  OA22X1 U24334 ( .IN1(n23019), .IN2(n21724), .IN3(n23018), .IN4(n21728), .Q(
        n21425) );
  OA22X1 U24335 ( .IN1(n23024), .IN2(n21726), .IN3(n23022), .IN4(n21746), .Q(
        n21424) );
  NAND4X0 U24336 ( .IN1(n21427), .IN2(n21426), .IN3(n21425), .IN4(n21424), 
        .QN(n21428) );
  NOR2X0 U24337 ( .IN1(n21429), .IN2(n21428), .QN(n21431) );
  NAND2X0 U24338 ( .IN1(n29331), .IN2(n23034), .QN(n21430) );
  NAND2X0 U24339 ( .IN1(n21431), .IN2(n21430), .QN(m5_data_o[12]) );
  OA22X1 U24340 ( .IN1(n23042), .IN2(n21724), .IN3(n21432), .IN4(n21736), .Q(
        n21440) );
  OA22X1 U24341 ( .IN1(n21434), .IN2(n21704), .IN3(n21433), .IN4(n21727), .Q(
        n21439) );
  OA22X1 U24342 ( .IN1(n21436), .IN2(n21745), .IN3(n21435), .IN4(n21735), .Q(
        n21438) );
  NAND2X0 U24343 ( .IN1(m0s10_data_i[13]), .IN2(n29336), .QN(n21437) );
  NAND4X0 U24344 ( .IN1(n21440), .IN2(n21439), .IN3(n21438), .IN4(n21437), 
        .QN(n21449) );
  OA22X1 U24345 ( .IN1(n23041), .IN2(n21728), .IN3(n21441), .IN4(n21712), .Q(
        n21447) );
  OA22X1 U24346 ( .IN1(n21443), .IN2(n21738), .IN3(n21442), .IN4(n21740), .Q(
        n21446) );
  OA22X1 U24347 ( .IN1(n23040), .IN2(n21742), .IN3(n23039), .IN4(n21726), .Q(
        n21445) );
  OA22X1 U24348 ( .IN1(n22793), .IN2(n21744), .IN3(n23043), .IN4(n21746), .Q(
        n21444) );
  NAND4X0 U24349 ( .IN1(n21447), .IN2(n21446), .IN3(n21445), .IN4(n21444), 
        .QN(n21448) );
  NOR2X0 U24350 ( .IN1(n21449), .IN2(n21448), .QN(n21451) );
  NAND2X0 U24351 ( .IN1(n29331), .IN2(n23053), .QN(n21450) );
  NAND2X0 U24352 ( .IN1(n21451), .IN2(n21450), .QN(m5_data_o[13]) );
  OA22X1 U24353 ( .IN1(n23061), .IN2(n21727), .IN3(n21452), .IN4(n21736), .Q(
        n21456) );
  OA22X1 U24354 ( .IN1(n23070), .IN2(n21726), .IN3(n23064), .IN4(n21712), .Q(
        n21455) );
  OA22X1 U24355 ( .IN1(n23062), .IN2(n21740), .IN3(n23058), .IN4(n21746), .Q(
        n21454) );
  NAND2X0 U24356 ( .IN1(m0s13_data_i[14]), .IN2(n29333), .QN(n21453) );
  NAND4X0 U24357 ( .IN1(n21456), .IN2(n21455), .IN3(n21454), .IN4(n21453), 
        .QN(n21467) );
  OA22X1 U24358 ( .IN1(n21457), .IN2(n21738), .IN3(n23068), .IN4(n21728), .Q(
        n21465) );
  OA22X1 U24359 ( .IN1(n23060), .IN2(n21742), .IN3(n21458), .IN4(n21735), .Q(
        n21464) );
  OA22X1 U24360 ( .IN1(n21460), .IN2(n21745), .IN3(n21459), .IN4(n21744), .Q(
        n21463) );
  OA22X1 U24361 ( .IN1(n23066), .IN2(n21724), .IN3(n21461), .IN4(n21730), .Q(
        n21462) );
  NAND4X0 U24362 ( .IN1(n21465), .IN2(n21464), .IN3(n21463), .IN4(n21462), 
        .QN(n21466) );
  NOR2X0 U24363 ( .IN1(n21467), .IN2(n21466), .QN(n21469) );
  NAND2X0 U24364 ( .IN1(n29331), .IN2(n23078), .QN(n21468) );
  NAND2X0 U24365 ( .IN1(n21469), .IN2(n21468), .QN(m5_data_o[14]) );
  OA22X1 U24366 ( .IN1(n21470), .IN2(n21742), .IN3(n23094), .IN4(n21738), .Q(
        n21476) );
  OA22X1 U24367 ( .IN1(n21471), .IN2(n21746), .IN3(n23084), .IN4(n21730), .Q(
        n21475) );
  OA22X1 U24368 ( .IN1(n23090), .IN2(n21744), .IN3(n21472), .IN4(n21736), .Q(
        n21474) );
  NAND2X0 U24369 ( .IN1(m0s13_data_i[15]), .IN2(n29333), .QN(n21473) );
  NAND4X0 U24370 ( .IN1(n21476), .IN2(n21475), .IN3(n21474), .IN4(n21473), 
        .QN(n21487) );
  OA22X1 U24371 ( .IN1(n23086), .IN2(n21727), .IN3(n21477), .IN4(n21724), .Q(
        n21485) );
  OA22X1 U24372 ( .IN1(n21478), .IN2(n21728), .IN3(n23088), .IN4(n21735), .Q(
        n21484) );
  OA22X1 U24373 ( .IN1(n21479), .IN2(n21745), .IN3(n23092), .IN4(n21740), .Q(
        n21483) );
  OA22X1 U24374 ( .IN1(n21481), .IN2(n21726), .IN3(n21480), .IN4(n21712), .Q(
        n21482) );
  NAND4X0 U24375 ( .IN1(n21485), .IN2(n21484), .IN3(n21483), .IN4(n21482), 
        .QN(n21486) );
  NOR2X0 U24376 ( .IN1(n21487), .IN2(n21486), .QN(n21489) );
  NAND2X0 U24377 ( .IN1(n29331), .IN2(n23103), .QN(n21488) );
  NAND2X0 U24378 ( .IN1(n21489), .IN2(n21488), .QN(m5_data_o[15]) );
  OA22X1 U24379 ( .IN1(n21744), .IN2(n21491), .IN3(n21742), .IN4(n21490), .Q(
        n21498) );
  OA22X1 U24380 ( .IN1(n21746), .IN2(n21493), .IN3(n21726), .IN4(n21492), .Q(
        n21497) );
  OA22X1 U24381 ( .IN1(n21704), .IN2(n22010), .IN3(n21712), .IN4(n21494), .Q(
        n21496) );
  NAND2X0 U24382 ( .IN1(n29347), .IN2(m0s0_data_i[16]), .QN(n21495) );
  NAND4X0 U24383 ( .IN1(n21498), .IN2(n21497), .IN3(n21496), .IN4(n21495), 
        .QN(n21509) );
  OA22X1 U24384 ( .IN1(n21740), .IN2(n21499), .IN3(n21735), .IN4(n22012), .Q(
        n21507) );
  OA22X1 U24385 ( .IN1(n21730), .IN2(n21501), .IN3(n21738), .IN4(n21500), .Q(
        n21506) );
  OA22X1 U24386 ( .IN1(n21727), .IN2(n21503), .IN3(n21745), .IN4(n21502), .Q(
        n21505) );
  OA22X1 U24387 ( .IN1(n21736), .IN2(n22009), .IN3(n21728), .IN4(n22011), .Q(
        n21504) );
  NAND4X0 U24388 ( .IN1(n21507), .IN2(n21506), .IN3(n21505), .IN4(n21504), 
        .QN(n21508) );
  NOR2X0 U24389 ( .IN1(n21509), .IN2(n21508), .QN(n21511) );
  NAND2X0 U24390 ( .IN1(s15_data_i[16]), .IN2(n21753), .QN(n21510) );
  NAND2X0 U24391 ( .IN1(n21511), .IN2(n21510), .QN(m5_data_o[16]) );
  OA22X1 U24392 ( .IN1(n21740), .IN2(n22397), .IN3(n21738), .IN4(n22831), .Q(
        n21517) );
  OA22X1 U24393 ( .IN1(n21730), .IN2(n22834), .IN3(n21728), .IN4(n22832), .Q(
        n21516) );
  OA22X1 U24394 ( .IN1(n21736), .IN2(n21513), .IN3(n21742), .IN4(n21512), .Q(
        n21515) );
  NAND2X0 U24395 ( .IN1(n29343), .IN2(m0s3_data_i[17]), .QN(n21514) );
  NAND4X0 U24396 ( .IN1(n21517), .IN2(n21516), .IN3(n21515), .IN4(n21514), 
        .QN(n21527) );
  OA22X1 U24397 ( .IN1(n21727), .IN2(n21518), .IN3(n21735), .IN4(n22837), .Q(
        n21525) );
  OA22X1 U24398 ( .IN1(n21746), .IN2(n22835), .IN3(n21726), .IN4(n21519), .Q(
        n21524) );
  OA22X1 U24399 ( .IN1(n21704), .IN2(n22836), .IN3(n21712), .IN4(n22833), .Q(
        n21523) );
  OA22X1 U24400 ( .IN1(n21745), .IN2(n21521), .IN3(n21724), .IN4(n21520), .Q(
        n21522) );
  NAND4X0 U24401 ( .IN1(n21525), .IN2(n21524), .IN3(n21523), .IN4(n21522), 
        .QN(n21526) );
  NOR2X0 U24402 ( .IN1(n21527), .IN2(n21526), .QN(n21529) );
  NAND2X0 U24403 ( .IN1(s15_data_i[17]), .IN2(n21753), .QN(n21528) );
  NAND2X0 U24404 ( .IN1(n21529), .IN2(n21528), .QN(m5_data_o[17]) );
  OA22X1 U24405 ( .IN1(n21736), .IN2(n22414), .IN3(n21746), .IN4(n21530), .Q(
        n21535) );
  OA22X1 U24406 ( .IN1(n21740), .IN2(n21531), .IN3(n21738), .IN4(n22411), .Q(
        n21534) );
  OA22X1 U24407 ( .IN1(n21744), .IN2(n22413), .IN3(n21724), .IN4(n22415), .Q(
        n21533) );
  NAND2X0 U24408 ( .IN1(n29332), .IN2(m0s14_data_i[18]), .QN(n21532) );
  NAND4X0 U24409 ( .IN1(n21535), .IN2(n21534), .IN3(n21533), .IN4(n21532), 
        .QN(n21546) );
  OA22X1 U24410 ( .IN1(n21728), .IN2(n21537), .IN3(n21712), .IN4(n21536), .Q(
        n21544) );
  OA22X1 U24411 ( .IN1(n21742), .IN2(n21538), .IN3(n21745), .IN4(n22412), .Q(
        n21543) );
  OA22X1 U24412 ( .IN1(n21735), .IN2(n22410), .IN3(n21704), .IN4(n21539), .Q(
        n21542) );
  OA22X1 U24413 ( .IN1(n21727), .IN2(n22037), .IN3(n21730), .IN4(n21540), .Q(
        n21541) );
  NAND4X0 U24414 ( .IN1(n21544), .IN2(n21543), .IN3(n21542), .IN4(n21541), 
        .QN(n21545) );
  NOR2X0 U24415 ( .IN1(n21546), .IN2(n21545), .QN(n21548) );
  NAND2X0 U24416 ( .IN1(s15_data_i[18]), .IN2(n21753), .QN(n21547) );
  NAND2X0 U24417 ( .IN1(n21548), .IN2(n21547), .QN(m5_data_o[18]) );
  OA22X1 U24418 ( .IN1(n21728), .IN2(n21549), .IN3(n21744), .IN4(n22431), .Q(
        n21555) );
  OA22X1 U24419 ( .IN1(n21740), .IN2(n21550), .IN3(n21735), .IN4(n22434), .Q(
        n21554) );
  OA22X1 U24420 ( .IN1(n21736), .IN2(n22050), .IN3(n21745), .IN4(n21551), .Q(
        n21553) );
  NAND2X0 U24421 ( .IN1(n29347), .IN2(m0s0_data_i[19]), .QN(n21552) );
  NAND4X0 U24422 ( .IN1(n21555), .IN2(n21554), .IN3(n21553), .IN4(n21552), 
        .QN(n21564) );
  OA22X1 U24423 ( .IN1(n21712), .IN2(n21556), .IN3(n21726), .IN4(n22428), .Q(
        n21562) );
  OA22X1 U24424 ( .IN1(n21727), .IN2(n21557), .IN3(n21746), .IN4(n22429), .Q(
        n21561) );
  OA22X1 U24425 ( .IN1(n21738), .IN2(n22435), .IN3(n21742), .IN4(n21558), .Q(
        n21560) );
  OA22X1 U24426 ( .IN1(n21730), .IN2(n22432), .IN3(n21704), .IN4(n22430), .Q(
        n21559) );
  NAND4X0 U24427 ( .IN1(n21562), .IN2(n21561), .IN3(n21560), .IN4(n21559), 
        .QN(n21563) );
  NOR2X0 U24428 ( .IN1(n21564), .IN2(n21563), .QN(n21566) );
  NAND2X0 U24429 ( .IN1(s15_data_i[19]), .IN2(n21753), .QN(n21565) );
  NAND2X0 U24430 ( .IN1(n21566), .IN2(n21565), .QN(m5_data_o[19]) );
  OA22X1 U24431 ( .IN1(n21742), .IN2(n22452), .IN3(n21726), .IN4(n22453), .Q(
        n21572) );
  OA22X1 U24432 ( .IN1(n21744), .IN2(n21568), .IN3(n21704), .IN4(n21567), .Q(
        n21571) );
  OA22X1 U24433 ( .IN1(n21745), .IN2(n22454), .IN3(n21724), .IN4(n22451), .Q(
        n21570) );
  NAND2X0 U24434 ( .IN1(n29337), .IN2(m0s9_data_i[20]), .QN(n21569) );
  NAND4X0 U24435 ( .IN1(n21572), .IN2(n21571), .IN3(n21570), .IN4(n21569), 
        .QN(n21583) );
  OA22X1 U24436 ( .IN1(n21736), .IN2(n22448), .IN3(n21740), .IN4(n21573), .Q(
        n21581) );
  OA22X1 U24437 ( .IN1(n21727), .IN2(n21575), .IN3(n21730), .IN4(n21574), .Q(
        n21580) );
  OA22X1 U24438 ( .IN1(n21728), .IN2(n22450), .IN3(n21738), .IN4(n21576), .Q(
        n21579) );
  OA22X1 U24439 ( .IN1(n21735), .IN2(n22449), .IN3(n21712), .IN4(n21577), .Q(
        n21578) );
  NAND4X0 U24440 ( .IN1(n21581), .IN2(n21580), .IN3(n21579), .IN4(n21578), 
        .QN(n21582) );
  NOR2X0 U24441 ( .IN1(n21583), .IN2(n21582), .QN(n21585) );
  NAND2X0 U24442 ( .IN1(s15_data_i[20]), .IN2(n21753), .QN(n21584) );
  NAND2X0 U24443 ( .IN1(n21585), .IN2(n21584), .QN(m5_data_o[20]) );
  OA22X1 U24444 ( .IN1(n21735), .IN2(n22852), .IN3(n21724), .IN4(n22853), .Q(
        n21591) );
  OA22X1 U24445 ( .IN1(n21730), .IN2(n22849), .IN3(n21726), .IN4(n21586), .Q(
        n21590) );
  OA22X1 U24446 ( .IN1(n21736), .IN2(n22851), .IN3(n21704), .IN4(n21587), .Q(
        n21589) );
  NAND2X0 U24447 ( .IN1(n29335), .IN2(m0s11_data_i[21]), .QN(n21588) );
  NAND4X0 U24448 ( .IN1(n21591), .IN2(n21590), .IN3(n21589), .IN4(n21588), 
        .QN(n21600) );
  OA22X1 U24449 ( .IN1(n21740), .IN2(n21592), .IN3(n21742), .IN4(n22856), .Q(
        n21598) );
  OA22X1 U24450 ( .IN1(n21727), .IN2(n22466), .IN3(n21712), .IN4(n22850), .Q(
        n21597) );
  OA22X1 U24451 ( .IN1(n21746), .IN2(n21594), .IN3(n21744), .IN4(n21593), .Q(
        n21596) );
  OA22X1 U24452 ( .IN1(n21738), .IN2(n22857), .IN3(n21745), .IN4(n22855), .Q(
        n21595) );
  NAND4X0 U24453 ( .IN1(n21598), .IN2(n21597), .IN3(n21596), .IN4(n21595), 
        .QN(n21599) );
  NOR2X0 U24454 ( .IN1(n21600), .IN2(n21599), .QN(n21602) );
  NAND2X0 U24455 ( .IN1(s15_data_i[21]), .IN2(n21753), .QN(n21601) );
  NAND2X0 U24456 ( .IN1(n21602), .IN2(n21601), .QN(m5_data_o[21]) );
  OA22X1 U24457 ( .IN1(n21730), .IN2(n22869), .IN3(n21735), .IN4(n22875), .Q(
        n21608) );
  OA22X1 U24458 ( .IN1(n21740), .IN2(n22873), .IN3(n21726), .IN4(n21603), .Q(
        n21607) );
  OA22X1 U24459 ( .IN1(n21742), .IN2(n22870), .IN3(n21724), .IN4(n21604), .Q(
        n21606) );
  NAND2X0 U24460 ( .IN1(n29335), .IN2(m0s11_data_i[22]), .QN(n21605) );
  NAND4X0 U24461 ( .IN1(n21608), .IN2(n21607), .IN3(n21606), .IN4(n21605), 
        .QN(n21618) );
  OA22X1 U24462 ( .IN1(n21736), .IN2(n21609), .IN3(n21745), .IN4(n22872), .Q(
        n21616) );
  OA22X1 U24463 ( .IN1(n21746), .IN2(n21610), .IN3(n21738), .IN4(n22874), .Q(
        n21615) );
  OA22X1 U24464 ( .IN1(n21744), .IN2(n22871), .IN3(n21704), .IN4(n21611), .Q(
        n21614) );
  OA22X1 U24465 ( .IN1(n21727), .IN2(n21612), .IN3(n21712), .IN4(n22876), .Q(
        n21613) );
  NAND4X0 U24466 ( .IN1(n21616), .IN2(n21615), .IN3(n21614), .IN4(n21613), 
        .QN(n21617) );
  NOR2X0 U24467 ( .IN1(n21618), .IN2(n21617), .QN(n21620) );
  NAND2X0 U24468 ( .IN1(s15_data_i[22]), .IN2(n21753), .QN(n21619) );
  NAND2X0 U24469 ( .IN1(n21620), .IN2(n21619), .QN(m5_data_o[22]) );
  OA22X1 U24470 ( .IN1(n21735), .IN2(n21622), .IN3(n21726), .IN4(n21621), .Q(
        n21629) );
  OA22X1 U24471 ( .IN1(n21736), .IN2(n21624), .IN3(n21742), .IN4(n21623), .Q(
        n21628) );
  OA22X1 U24472 ( .IN1(n21727), .IN2(n22491), .IN3(n21745), .IN4(n21625), .Q(
        n21627) );
  NAND2X0 U24473 ( .IN1(n29342), .IN2(m0s4_data_i[23]), .QN(n21626) );
  NAND4X0 U24474 ( .IN1(n21629), .IN2(n21628), .IN3(n21627), .IN4(n21626), 
        .QN(n21640) );
  OA22X1 U24475 ( .IN1(n21728), .IN2(n21630), .IN3(n21738), .IN4(n22495), .Q(
        n21638) );
  OA22X1 U24476 ( .IN1(n21730), .IN2(n22494), .IN3(n21744), .IN4(n21631), .Q(
        n21637) );
  OA22X1 U24477 ( .IN1(n21746), .IN2(n21633), .IN3(n21704), .IN4(n21632), .Q(
        n21636) );
  OA22X1 U24478 ( .IN1(n21740), .IN2(n22492), .IN3(n21724), .IN4(n21634), .Q(
        n21635) );
  NAND4X0 U24479 ( .IN1(n21638), .IN2(n21637), .IN3(n21636), .IN4(n21635), 
        .QN(n21639) );
  NOR2X0 U24480 ( .IN1(n21640), .IN2(n21639), .QN(n21642) );
  NAND2X0 U24481 ( .IN1(s15_data_i[23]), .IN2(n21753), .QN(n21641) );
  NAND2X0 U24482 ( .IN1(n21642), .IN2(n21641), .QN(m5_data_o[23]) );
  OA22X1 U24483 ( .IN1(n21744), .IN2(n21643), .IN3(n21704), .IN4(n22888), .Q(
        n21648) );
  OA22X1 U24484 ( .IN1(n21730), .IN2(n22892), .IN3(n21712), .IN4(n21644), .Q(
        n21647) );
  OA22X1 U24485 ( .IN1(n21736), .IN2(n22895), .IN3(n21726), .IN4(n22893), .Q(
        n21646) );
  NAND2X0 U24486 ( .IN1(n29340), .IN2(m0s6_data_i[24]), .QN(n21645) );
  NAND4X0 U24487 ( .IN1(n21648), .IN2(n21647), .IN3(n21646), .IN4(n21645), 
        .QN(n21659) );
  OA22X1 U24488 ( .IN1(n21746), .IN2(n21650), .IN3(n21724), .IN4(n21649), .Q(
        n21657) );
  OA22X1 U24489 ( .IN1(n21727), .IN2(n22896), .IN3(n21728), .IN4(n21651), .Q(
        n21656) );
  OA22X1 U24490 ( .IN1(n21735), .IN2(n21652), .IN3(n21742), .IN4(n22890), .Q(
        n21655) );
  OA22X1 U24491 ( .IN1(n21740), .IN2(n21653), .IN3(n21738), .IN4(n22891), .Q(
        n21654) );
  NAND4X0 U24492 ( .IN1(n21657), .IN2(n21656), .IN3(n21655), .IN4(n21654), 
        .QN(n21658) );
  NOR2X0 U24493 ( .IN1(n21659), .IN2(n21658), .QN(n21661) );
  NAND2X0 U24494 ( .IN1(s15_data_i[24]), .IN2(n21753), .QN(n21660) );
  NAND2X0 U24495 ( .IN1(n21661), .IN2(n21660), .QN(m5_data_o[24]) );
  OA22X1 U24496 ( .IN1(n21727), .IN2(n21662), .IN3(n21726), .IN4(n22524), .Q(
        n21669) );
  OA22X1 U24497 ( .IN1(n21736), .IN2(n22525), .IN3(n21742), .IN4(n21663), .Q(
        n21668) );
  OA22X1 U24498 ( .IN1(n21712), .IN2(n21665), .IN3(n21724), .IN4(n21664), .Q(
        n21667) );
  NAND2X0 U24499 ( .IN1(n29333), .IN2(m0s13_data_i[25]), .QN(n21666) );
  NAND4X0 U24500 ( .IN1(n21669), .IN2(n21668), .IN3(n21667), .IN4(n21666), 
        .QN(n21678) );
  OA22X1 U24501 ( .IN1(n21728), .IN2(n21670), .IN3(n21745), .IN4(n22119), .Q(
        n21676) );
  OA22X1 U24502 ( .IN1(n21746), .IN2(n22520), .IN3(n21744), .IN4(n22521), .Q(
        n21675) );
  OA22X1 U24503 ( .IN1(n21740), .IN2(n21671), .IN3(n21735), .IN4(n22522), .Q(
        n21674) );
  OA22X1 U24504 ( .IN1(n21730), .IN2(n22523), .IN3(n21738), .IN4(n21672), .Q(
        n21673) );
  NAND4X0 U24505 ( .IN1(n21676), .IN2(n21675), .IN3(n21674), .IN4(n21673), 
        .QN(n21677) );
  NOR2X0 U24506 ( .IN1(n21678), .IN2(n21677), .QN(n21680) );
  NAND2X0 U24507 ( .IN1(s15_data_i[25]), .IN2(n21753), .QN(n21679) );
  NAND2X0 U24508 ( .IN1(n21680), .IN2(n21679), .QN(m5_data_o[25]) );
  OA22X1 U24509 ( .IN1(n21742), .IN2(n21682), .IN3(n21726), .IN4(n21681), .Q(
        n21690) );
  OA22X1 U24510 ( .IN1(n21736), .IN2(n21684), .IN3(n21738), .IN4(n21683), .Q(
        n21689) );
  OA22X1 U24511 ( .IN1(n21735), .IN2(n21686), .IN3(n21712), .IN4(n21685), .Q(
        n21688) );
  NAND2X0 U24512 ( .IN1(n29340), .IN2(m0s6_data_i[26]), .QN(n21687) );
  NAND4X0 U24513 ( .IN1(n21690), .IN2(n21689), .IN3(n21688), .IN4(n21687), 
        .QN(n21701) );
  OA22X1 U24514 ( .IN1(n21740), .IN2(n22538), .IN3(n21704), .IN4(n21691), .Q(
        n21699) );
  OA22X1 U24515 ( .IN1(n21728), .IN2(n22541), .IN3(n21724), .IN4(n21692), .Q(
        n21698) );
  OA22X1 U24516 ( .IN1(n21730), .IN2(n22540), .IN3(n21746), .IN4(n21693), .Q(
        n21697) );
  OA22X1 U24517 ( .IN1(n21727), .IN2(n21695), .IN3(n21744), .IN4(n21694), .Q(
        n21696) );
  NAND4X0 U24518 ( .IN1(n21699), .IN2(n21698), .IN3(n21697), .IN4(n21696), 
        .QN(n21700) );
  NOR2X0 U24519 ( .IN1(n21701), .IN2(n21700), .QN(n21703) );
  NAND2X0 U24520 ( .IN1(s15_data_i[26]), .IN2(n21753), .QN(n21702) );
  NAND2X0 U24521 ( .IN1(n21703), .IN2(n21702), .QN(m5_data_o[26]) );
  OA22X1 U24522 ( .IN1(n21742), .IN2(n22916), .IN3(n21704), .IN4(n22918), .Q(
        n21709) );
  OA22X1 U24523 ( .IN1(n21740), .IN2(n22913), .IN3(n21735), .IN4(n22915), .Q(
        n21708) );
  OA22X1 U24524 ( .IN1(n21736), .IN2(n21705), .IN3(n21730), .IN4(n22911), .Q(
        n21707) );
  NAND2X0 U24525 ( .IN1(n29347), .IN2(m0s0_data_i[27]), .QN(n21706) );
  NAND4X0 U24526 ( .IN1(n21709), .IN2(n21708), .IN3(n21707), .IN4(n21706), 
        .QN(n21721) );
  OA22X1 U24527 ( .IN1(n21712), .IN2(n21711), .IN3(n21726), .IN4(n21710), .Q(
        n21719) );
  OA22X1 U24528 ( .IN1(n21728), .IN2(n21713), .IN3(n21744), .IN4(n22912), .Q(
        n21718) );
  OA22X1 U24529 ( .IN1(n21727), .IN2(n22910), .IN3(n21746), .IN4(n21714), .Q(
        n21717) );
  OA22X1 U24530 ( .IN1(n21738), .IN2(n22908), .IN3(n21745), .IN4(n21715), .Q(
        n21716) );
  NAND4X0 U24531 ( .IN1(n21719), .IN2(n21718), .IN3(n21717), .IN4(n21716), 
        .QN(n21720) );
  NOR2X0 U24532 ( .IN1(n21721), .IN2(n21720), .QN(n21723) );
  NAND2X0 U24533 ( .IN1(s15_data_i[27]), .IN2(n21753), .QN(n21722) );
  NAND2X0 U24534 ( .IN1(n21723), .IN2(n21722), .QN(m5_data_o[27]) );
  OA22X1 U24535 ( .IN1(n21704), .IN2(n22932), .IN3(n21724), .IN4(n22568), .Q(
        n21734) );
  OA22X1 U24536 ( .IN1(n21727), .IN2(n22941), .IN3(n21726), .IN4(n21725), .Q(
        n21733) );
  OA22X1 U24537 ( .IN1(n21730), .IN2(n21729), .IN3(n21728), .IN4(n22930), .Q(
        n21732) );
  NAND2X0 U24538 ( .IN1(n29342), .IN2(m0s4_data_i[28]), .QN(n21731) );
  NAND4X0 U24539 ( .IN1(n21734), .IN2(n21733), .IN3(n21732), .IN4(n21731), 
        .QN(n21752) );
  OA22X1 U24540 ( .IN1(n21736), .IN2(n22936), .IN3(n21735), .IN4(n22935), .Q(
        n21750) );
  OA22X1 U24541 ( .IN1(n21740), .IN2(n21739), .IN3(n21738), .IN4(n21737), .Q(
        n21749) );
  OA22X1 U24542 ( .IN1(n21744), .IN2(n21743), .IN3(n21742), .IN4(n21741), .Q(
        n21748) );
  OA22X1 U24543 ( .IN1(n21746), .IN2(n22934), .IN3(n21745), .IN4(n22940), .Q(
        n21747) );
  NAND4X0 U24544 ( .IN1(n21750), .IN2(n21749), .IN3(n21748), .IN4(n21747), 
        .QN(n21751) );
  NOR2X0 U24545 ( .IN1(n21752), .IN2(n21751), .QN(n21755) );
  NAND2X0 U24546 ( .IN1(s15_data_i[28]), .IN2(n21753), .QN(n21754) );
  NAND2X0 U24547 ( .IN1(n21755), .IN2(n21754), .QN(m5_data_o[28]) );
  NOR2X0 U24548 ( .IN1(\s15/next ), .IN2(\s15/msel/pri_out [0]), .QN(n21761)
         );
  AND3X1 U24549 ( .IN1(n13590), .IN2(m6s15_cyc), .IN3(n34598), .Q(n34043) );
  NAND3X0 U24550 ( .IN1(n13538), .IN2(m7s15_cyc), .IN3(n34518), .QN(n34028) );
  INVX0 U24551 ( .INP(n34028), .ZN(n33987) );
  NOR2X0 U24552 ( .IN1(n34043), .IN2(n33987), .QN(n34005) );
  NAND3X0 U24553 ( .IN1(n13642), .IN2(m5s15_cyc), .IN3(n34517), .QN(n34061) );
  NAND3X0 U24554 ( .IN1(n13694), .IN2(m4s15_cyc), .IN3(n34516), .QN(n34022) );
  AND2X1 U24555 ( .IN1(n34061), .IN2(n34022), .Q(n34007) );
  NAND2X0 U24556 ( .IN1(n34005), .IN2(n34007), .QN(n33997) );
  NAND3X0 U24557 ( .IN1(n13746), .IN2(m3s15_cyc), .IN3(n34515), .QN(n34029) );
  INVX0 U24558 ( .INP(n34029), .ZN(n34012) );
  AND3X1 U24559 ( .IN1(n13798), .IN2(m2s15_cyc), .IN3(n34602), .Q(n34040) );
  NOR2X0 U24560 ( .IN1(n34012), .IN2(n34040), .QN(n34008) );
  NAND3X0 U24561 ( .IN1(n13850), .IN2(m1s15_cyc), .IN3(n34514), .QN(n34049) );
  INVX0 U24562 ( .INP(n34049), .ZN(n33994) );
  NAND3X0 U24563 ( .IN1(n13914), .IN2(m0s15_cyc), .IN3(n34482), .QN(n34051) );
  INVX0 U24564 ( .INP(n34051), .ZN(n34035) );
  NOR2X0 U24565 ( .IN1(n33994), .IN2(n34035), .QN(n34003) );
  NAND2X0 U24566 ( .IN1(n34008), .IN2(n34003), .QN(n33988) );
  NOR2X0 U24567 ( .IN1(n33997), .IN2(n33988), .QN(n34219) );
  NAND2X0 U24568 ( .IN1(n33880), .IN2(n33895), .QN(n33881) );
  NAND2X0 U24569 ( .IN1(n21757), .IN2(n21756), .QN(n33887) );
  OR2X1 U24570 ( .IN1(n33881), .IN2(n33887), .Q(n33873) );
  NAND2X0 U24571 ( .IN1(n33871), .IN2(n33870), .QN(n33878) );
  INVX0 U24572 ( .INP(n33878), .ZN(n33884) );
  NAND3X0 U24573 ( .IN1(n33884), .IN2(n33889), .IN3(n33888), .QN(n33866) );
  NAND3X0 U24574 ( .IN1(m0s15_cyc), .IN2(n34298), .IN3(n34482), .QN(n33852) );
  NAND3X0 U24575 ( .IN1(m1s15_cyc), .IN2(n34302), .IN3(n34514), .QN(n33833) );
  NAND2X0 U24576 ( .IN1(n33852), .IN2(n33833), .QN(n33779) );
  INVX0 U24577 ( .INP(n33779), .ZN(n33776) );
  NAND3X0 U24578 ( .IN1(m3s15_cyc), .IN2(n34303), .IN3(n34515), .QN(n33803) );
  NAND3X0 U24579 ( .IN1(m2s15_cyc), .IN2(n34359), .IN3(n34602), .QN(n33853) );
  NAND2X0 U24580 ( .IN1(n33803), .IN2(n33853), .QN(n33774) );
  INVX0 U24581 ( .INP(n33774), .ZN(n33773) );
  NAND3X0 U24582 ( .IN1(m4s15_cyc), .IN2(n34299), .IN3(n34516), .QN(n33822) );
  INVX0 U24583 ( .INP(n33822), .ZN(n33818) );
  NAND3X0 U24584 ( .IN1(m5s15_cyc), .IN2(n34300), .IN3(n34517), .QN(n33814) );
  INVX0 U24585 ( .INP(n33814), .ZN(n33817) );
  NOR2X0 U24586 ( .IN1(n33818), .IN2(n33817), .QN(n33793) );
  NAND3X0 U24587 ( .IN1(m6s15_cyc), .IN2(n34360), .IN3(n34598), .QN(n33827) );
  INVX0 U24588 ( .INP(n33827), .ZN(n33815) );
  NAND3X0 U24589 ( .IN1(m7s15_cyc), .IN2(n34301), .IN3(n34518), .QN(n33812) );
  INVX0 U24590 ( .INP(n33812), .ZN(n33823) );
  NOR2X0 U24591 ( .IN1(n33815), .IN2(n33823), .QN(n33792) );
  NAND2X0 U24592 ( .IN1(n33793), .IN2(n33792), .QN(n33769) );
  INVX0 U24593 ( .INP(n33769), .ZN(n21758) );
  NAND4X0 U24594 ( .IN1(n33776), .IN2(n33773), .IN3(n21758), .IN4(\s15/next ), 
        .QN(n34220) );
  AO221X1 U24595 ( .IN1(n34219), .IN2(n33873), .IN3(n34219), .IN4(n33866), 
        .IN5(n34220), .Q(n21759) );
  NAND2X0 U24596 ( .IN1(n34694), .IN2(n21759), .QN(n21760) );
  NOR2X0 U24597 ( .IN1(n21761), .IN2(n21760), .QN(n17569) );
  NOR2X0 U24598 ( .IN1(\s14/next ), .IN2(\s14/msel/pri_out [1]), .QN(n21769)
         );
  INVX0 U24599 ( .INP(n21762), .ZN(n33543) );
  AND2X1 U24600 ( .IN1(n33543), .IN2(n21763), .Q(n34211) );
  NOR2X0 U24601 ( .IN1(n21764), .IN2(n33545), .QN(n34210) );
  INVX0 U24602 ( .INP(n21765), .ZN(n33708) );
  NOR2X0 U24603 ( .IN1(n33705), .IN2(n21766), .QN(n33716) );
  AND4X1 U24604 ( .IN1(n33708), .IN2(n33707), .IN3(n33716), .IN4(\s14/next ), 
        .Q(n34217) );
  NAND3X0 U24605 ( .IN1(n34211), .IN2(n34210), .IN3(n34217), .QN(n21767) );
  NAND2X0 U24606 ( .IN1(n34679), .IN2(n21767), .QN(n21768) );
  NOR2X0 U24607 ( .IN1(n21769), .IN2(n21768), .QN(n17570) );
  NOR2X0 U24608 ( .IN1(\s10/next ), .IN2(\s10/msel/pri_out [0]), .QN(n21781)
         );
  OR2X1 U24609 ( .IN1(n21770), .IN2(n32704), .Q(n32697) );
  NAND2X0 U24610 ( .IN1(n21771), .IN2(n32702), .QN(n32709) );
  NOR2X0 U24611 ( .IN1(n32697), .IN2(n32709), .QN(n34166) );
  NAND2X0 U24612 ( .IN1(n32578), .IN2(n32577), .QN(n32582) );
  NAND2X0 U24613 ( .IN1(n32583), .IN2(n32581), .QN(n32579) );
  NOR2X0 U24614 ( .IN1(n32582), .IN2(n32579), .QN(n32570) );
  INVX0 U24615 ( .INP(n32570), .ZN(n21778) );
  NOR2X0 U24616 ( .IN1(n21772), .IN2(n32567), .QN(n32580) );
  AND2X1 U24617 ( .IN1(n32565), .IN2(n32566), .Q(n32589) );
  NAND2X0 U24618 ( .IN1(n32580), .IN2(n32589), .QN(n32563) );
  NAND3X0 U24619 ( .IN1(m5s10_cyc), .IN2(n34323), .IN3(n34504), .QN(n32509) );
  NAND2X0 U24620 ( .IN1(m4s10_cyc), .IN2(n34583), .QN(n21773) );
  NOR2X0 U24621 ( .IN1(n13697), .IN2(n21773), .QN(n32539) );
  INVX0 U24622 ( .INP(n32539), .ZN(n32512) );
  NAND2X0 U24623 ( .IN1(n32509), .IN2(n32512), .QN(n32482) );
  INVX0 U24624 ( .INP(n32482), .ZN(n32473) );
  NAND2X0 U24625 ( .IN1(m6s10_cyc), .IN2(n34568), .QN(n21774) );
  NOR2X0 U24626 ( .IN1(n13593), .IN2(n21774), .QN(n32511) );
  NAND3X0 U24627 ( .IN1(m7s10_cyc), .IN2(n34353), .IN3(n34505), .QN(n32508) );
  INVX0 U24628 ( .INP(n32508), .ZN(n32527) );
  NOR2X0 U24629 ( .IN1(n32511), .IN2(n32527), .QN(n32480) );
  NAND2X0 U24630 ( .IN1(n32473), .IN2(n32480), .QN(n32463) );
  NAND2X0 U24631 ( .IN1(m0s10_cyc), .IN2(n34582), .QN(n21775) );
  NOR2X0 U24632 ( .IN1(n13920), .IN2(n21775), .QN(n32549) );
  NAND2X0 U24633 ( .IN1(m1s10_cyc), .IN2(n34611), .QN(n21776) );
  NOR2X0 U24634 ( .IN1(n13853), .IN2(n21776), .QN(n32505) );
  NOR2X0 U24635 ( .IN1(n32549), .IN2(n32505), .QN(n32481) );
  NAND3X0 U24636 ( .IN1(m2s10_cyc), .IN2(n34322), .IN3(n34503), .QN(n32526) );
  INVX0 U24637 ( .INP(n32526), .ZN(n32550) );
  AND3X1 U24638 ( .IN1(m3s10_cyc), .IN2(n34606), .IN3(n34372), .Q(n32513) );
  NOR2X0 U24639 ( .IN1(n32550), .IN2(n32513), .QN(n32460) );
  NAND2X0 U24640 ( .IN1(n32481), .IN2(n32460), .QN(n32459) );
  NOR3X0 U24641 ( .IN1(n32463), .IN2(n32459), .IN3(n34376), .QN(n34165) );
  INVX0 U24642 ( .INP(n34165), .ZN(n21777) );
  AO221X1 U24643 ( .IN1(n34166), .IN2(n21778), .IN3(n34166), .IN4(n32563), 
        .IN5(n21777), .Q(n21779) );
  NAND2X0 U24644 ( .IN1(n34695), .IN2(n21779), .QN(n21780) );
  NOR2X0 U24645 ( .IN1(n21781), .IN2(n21780), .QN(n17579) );
  NOR2X0 U24646 ( .IN1(\s7/next ), .IN2(\s7/msel/pri_out [1]), .QN(n21786) );
  NAND3X0 U24647 ( .IN1(n13894), .IN2(m0s7_cyc), .IN3(n34497), .QN(n31895) );
  NAND3X0 U24648 ( .IN1(n13838), .IN2(m1s7_cyc), .IN3(n34533), .QN(n31898) );
  NAND2X0 U24649 ( .IN1(n31895), .IN2(n31898), .QN(n31873) );
  INVX0 U24650 ( .INP(n31873), .ZN(n34133) );
  AND3X1 U24651 ( .IN1(n13786), .IN2(m2s7_cyc), .IN3(n34600), .Q(n31906) );
  NAND3X0 U24652 ( .IN1(n13734), .IN2(m3s7_cyc), .IN3(n34498), .QN(n31890) );
  INVX0 U24653 ( .INP(n31890), .ZN(n31917) );
  NOR2X0 U24654 ( .IN1(n31906), .IN2(n31917), .QN(n34134) );
  NAND3X0 U24655 ( .IN1(n13578), .IN2(m6s7_cyc), .IN3(n34567), .QN(n31916) );
  NAND3X0 U24656 ( .IN1(n13526), .IN2(m7s7_cyc), .IN3(n34499), .QN(n31892) );
  NAND2X0 U24657 ( .IN1(n31916), .IN2(n31892), .QN(n31867) );
  INVX0 U24658 ( .INP(n31867), .ZN(n31858) );
  NAND3X0 U24659 ( .IN1(n13630), .IN2(m5s7_cyc), .IN3(n34534), .QN(n31891) );
  INVX0 U24660 ( .INP(n31891), .ZN(n31902) );
  NAND3X0 U24661 ( .IN1(n13682), .IN2(m4s7_cyc), .IN3(n34594), .QN(n31908) );
  INVX0 U24662 ( .INP(n31908), .ZN(n31893) );
  NOR2X0 U24663 ( .IN1(n31902), .IN2(n31893), .QN(n31868) );
  AND2X1 U24664 ( .IN1(n31858), .IN2(n31868), .Q(n34132) );
  INVX0 U24665 ( .INP(n31629), .ZN(n21782) );
  NAND2X0 U24666 ( .IN1(n21783), .IN2(n21782), .QN(n31637) );
  NOR4X0 U24667 ( .IN1(n31630), .IN2(n31635), .IN3(n31637), .IN4(n34377), .QN(
        n34135) );
  NAND4X0 U24668 ( .IN1(n34133), .IN2(n34134), .IN3(n34132), .IN4(n34135), 
        .QN(n21784) );
  NAND2X0 U24669 ( .IN1(n34696), .IN2(n21784), .QN(n21785) );
  NOR2X0 U24670 ( .IN1(n21786), .IN2(n21785), .QN(n17584) );
  NOR2X0 U24671 ( .IN1(\s5/next ), .IN2(\s5/msel/pri_out [1]), .QN(n21791) );
  NAND3X0 U24672 ( .IN1(n13576), .IN2(m6s5_cyc), .IN3(n34529), .QN(n31273) );
  NAND3X0 U24673 ( .IN1(n13524), .IN2(m7s5_cyc), .IN3(n34530), .QN(n31287) );
  NAND2X0 U24674 ( .IN1(n31273), .IN2(n31287), .QN(n31248) );
  NAND3X0 U24675 ( .IN1(n13628), .IN2(m5s5_cyc), .IN3(n34528), .QN(n31324) );
  NAND3X0 U24676 ( .IN1(n13680), .IN2(m4s5_cyc), .IN3(n34496), .QN(n31297) );
  NAND2X0 U24677 ( .IN1(n31324), .IN2(n31297), .QN(n31260) );
  NOR2X0 U24678 ( .IN1(n31248), .IN2(n31260), .QN(n34106) );
  NAND3X0 U24679 ( .IN1(n13890), .IN2(m0s5_cyc), .IN3(n34493), .QN(n31294) );
  NAND3X0 U24680 ( .IN1(n13836), .IN2(m1s5_cyc), .IN3(n34494), .QN(n31288) );
  NAND2X0 U24681 ( .IN1(n31294), .IN2(n31288), .QN(n31257) );
  NAND3X0 U24682 ( .IN1(n13732), .IN2(m3s5_cyc), .IN3(n34495), .QN(n31284) );
  INVX0 U24683 ( .INP(n31284), .ZN(n31251) );
  NAND3X0 U24684 ( .IN1(n13784), .IN2(m2s5_cyc), .IN3(n34370), .QN(n31318) );
  INVX0 U24685 ( .INP(n31318), .ZN(n31285) );
  NOR2X0 U24686 ( .IN1(n31251), .IN2(n31285), .QN(n31256) );
  INVX0 U24687 ( .INP(n31256), .ZN(n21787) );
  NOR2X0 U24688 ( .IN1(n31257), .IN2(n21787), .QN(n34105) );
  NAND3X0 U24689 ( .IN1(m0s5_cyc), .IN2(n34344), .IN3(n34493), .QN(n31057) );
  NAND3X0 U24690 ( .IN1(m1s5_cyc), .IN2(n34343), .IN3(n34494), .QN(n31021) );
  NAND2X0 U24691 ( .IN1(n31057), .IN2(n31021), .QN(n31001) );
  INVX0 U24692 ( .INP(n31001), .ZN(n30983) );
  NAND3X0 U24693 ( .IN1(m3s5_cyc), .IN2(n34317), .IN3(n34495), .QN(n31036) );
  INVX0 U24694 ( .INP(n31036), .ZN(n31016) );
  NAND3X0 U24695 ( .IN1(m2s5_cyc), .IN2(n34587), .IN3(n34370), .QN(n31053) );
  INVX0 U24696 ( .INP(n31053), .ZN(n30977) );
  NOR2X0 U24697 ( .IN1(n31016), .IN2(n30977), .QN(n30991) );
  NAND3X0 U24698 ( .IN1(m4s5_cyc), .IN2(n34235), .IN3(n34496), .QN(n31038) );
  NAND3X0 U24699 ( .IN1(m5s5_cyc), .IN2(n34342), .IN3(n34528), .QN(n31023) );
  NAND2X0 U24700 ( .IN1(n31038), .IN2(n31023), .QN(n30992) );
  NAND3X0 U24701 ( .IN1(m6s5_cyc), .IN2(n34341), .IN3(n34529), .QN(n31008) );
  INVX0 U24702 ( .INP(n31008), .ZN(n31046) );
  NAND3X0 U24703 ( .IN1(m7s5_cyc), .IN2(n34316), .IN3(n34530), .QN(n31019) );
  INVX0 U24704 ( .INP(n31019), .ZN(n31007) );
  NOR2X0 U24705 ( .IN1(n31046), .IN2(n31007), .QN(n30997) );
  INVX0 U24706 ( .INP(n30997), .ZN(n21788) );
  NOR2X0 U24707 ( .IN1(n30992), .IN2(n21788), .QN(n30982) );
  AND4X1 U24708 ( .IN1(n30983), .IN2(n30991), .IN3(n30982), .IN4(\s5/next ), 
        .Q(n34107) );
  NAND3X0 U24709 ( .IN1(n34106), .IN2(n34105), .IN3(n34107), .QN(n21789) );
  NAND2X0 U24710 ( .IN1(n34687), .IN2(n21789), .QN(n21790) );
  NOR2X0 U24711 ( .IN1(n21791), .IN2(n21790), .QN(n17588) );
  NOR2X0 U24712 ( .IN1(\s4/next ), .IN2(\s4/msel/pri_out [1]), .QN(n21796) );
  NAND3X0 U24713 ( .IN1(m5s4_cyc), .IN2(n34313), .IN3(n34492), .QN(n30681) );
  NAND3X0 U24714 ( .IN1(m4s4_cyc), .IN2(n34338), .IN3(n34525), .QN(n30678) );
  NAND2X0 U24715 ( .IN1(n30681), .IN2(n30678), .QN(n30641) );
  NAND3X0 U24716 ( .IN1(m6s4_cyc), .IN2(n34339), .IN3(n34526), .QN(n30679) );
  NAND3X0 U24717 ( .IN1(m7s4_cyc), .IN2(n34314), .IN3(n34527), .QN(n30690) );
  NAND2X0 U24718 ( .IN1(n30679), .IN2(n30690), .QN(n30626) );
  NOR2X0 U24719 ( .IN1(n30641), .IN2(n30626), .QN(n34101) );
  NAND3X0 U24720 ( .IN1(m0s4_cyc), .IN2(n34340), .IN3(n34490), .QN(n30667) );
  NAND3X0 U24721 ( .IN1(m1s4_cyc), .IN2(n34315), .IN3(n34491), .QN(n30705) );
  NAND2X0 U24722 ( .IN1(n30667), .IN2(n30705), .QN(n30642) );
  NAND2X0 U24723 ( .IN1(m2s4_cyc), .IN2(n34577), .QN(n21792) );
  NOR2X0 U24724 ( .IN1(n13783), .IN2(n21792), .QN(n30707) );
  INVX0 U24725 ( .INP(n30707), .ZN(n30668) );
  NAND2X0 U24726 ( .IN1(m3s4_cyc), .IN2(n34578), .QN(n21793) );
  NOR2X0 U24727 ( .IN1(n13731), .IN2(n21793), .QN(n30666) );
  INVX0 U24728 ( .INP(n30666), .ZN(n30682) );
  NAND2X0 U24729 ( .IN1(n30668), .IN2(n30682), .QN(n30647) );
  NOR2X0 U24730 ( .IN1(n30642), .IN2(n30647), .QN(n34100) );
  NAND3X0 U24731 ( .IN1(n13888), .IN2(m0s4_cyc), .IN3(n34490), .QN(n30941) );
  NAND3X0 U24732 ( .IN1(n13835), .IN2(m1s4_cyc), .IN3(n34491), .QN(n30931) );
  NAND2X0 U24733 ( .IN1(n30941), .IN2(n30931), .QN(n30909) );
  INVX0 U24734 ( .INP(n30909), .ZN(n30884) );
  NAND3X0 U24735 ( .IN1(n13731), .IN2(m3s4_cyc), .IN3(n34578), .QN(n30926) );
  INVX0 U24736 ( .INP(n30926), .ZN(n30888) );
  NAND3X0 U24737 ( .IN1(n13783), .IN2(m2s4_cyc), .IN3(n34577), .QN(n30961) );
  INVX0 U24738 ( .INP(n30961), .ZN(n30928) );
  NOR2X0 U24739 ( .IN1(n30888), .IN2(n30928), .QN(n30910) );
  NAND3X0 U24740 ( .IN1(n13575), .IN2(m6s4_cyc), .IN3(n34526), .QN(n30945) );
  INVX0 U24741 ( .INP(n30945), .ZN(n30949) );
  NAND3X0 U24742 ( .IN1(n13679), .IN2(m4s4_cyc), .IN3(n34525), .QN(n30900) );
  INVX0 U24743 ( .INP(n30900), .ZN(n30947) );
  NOR2X0 U24744 ( .IN1(n30949), .IN2(n30947), .QN(n30933) );
  NAND3X0 U24745 ( .IN1(n13523), .IN2(m7s4_cyc), .IN3(n34527), .QN(n30930) );
  NAND3X0 U24746 ( .IN1(n13627), .IN2(m5s4_cyc), .IN3(n34492), .QN(n30927) );
  AND3X1 U24747 ( .IN1(n30933), .IN2(n30930), .IN3(n30927), .Q(n30890) );
  AND4X1 U24748 ( .IN1(n30884), .IN2(n30910), .IN3(n30890), .IN4(\s4/next ), 
        .Q(n34097) );
  NAND3X0 U24749 ( .IN1(n34101), .IN2(n34100), .IN3(n34097), .QN(n21794) );
  NAND2X0 U24750 ( .IN1(n34697), .IN2(n21794), .QN(n21795) );
  NOR2X0 U24751 ( .IN1(n21796), .IN2(n21795), .QN(n17590) );
  NOR2X0 U24752 ( .IN1(\s3/next ), .IN2(\s3/msel/pri_out [0]), .QN(n21805) );
  NAND3X0 U24753 ( .IN1(n13790), .IN2(m2s3_cyc), .IN3(n34595), .QN(n30610) );
  NAND3X0 U24754 ( .IN1(n13738), .IN2(m3s3_cyc), .IN3(n34564), .QN(n30576) );
  NAND2X0 U24755 ( .IN1(n30610), .IN2(n30576), .QN(n30541) );
  NAND3X0 U24756 ( .IN1(n13902), .IN2(m0s3_cyc), .IN3(n34485), .QN(n30591) );
  NAND3X0 U24757 ( .IN1(n13842), .IN2(m1s3_cyc), .IN3(n34486), .QN(n30580) );
  NAND2X0 U24758 ( .IN1(n30591), .IN2(n30580), .QN(n30560) );
  NOR2X0 U24759 ( .IN1(n30541), .IN2(n30560), .QN(n30548) );
  NAND3X0 U24760 ( .IN1(n13686), .IN2(m4s3_cyc), .IN3(n34487), .QN(n30549) );
  INVX0 U24761 ( .INP(n30549), .ZN(n30597) );
  NAND3X0 U24762 ( .IN1(n13634), .IN2(m5s3_cyc), .IN3(n34551), .QN(n30577) );
  INVX0 U24763 ( .INP(n30577), .ZN(n30618) );
  NAND3X0 U24764 ( .IN1(n13582), .IN2(m6s3_cyc), .IN3(n34488), .QN(n30594) );
  NAND3X0 U24765 ( .IN1(n13530), .IN2(m7s3_cyc), .IN3(n34489), .QN(n30579) );
  NAND2X0 U24766 ( .IN1(n30594), .IN2(n30579), .QN(n30557) );
  NOR3X0 U24767 ( .IN1(n30597), .IN2(n30618), .IN3(n30557), .QN(n30544) );
  NAND2X0 U24768 ( .IN1(n30548), .IN2(n30544), .QN(n34095) );
  INVX0 U24769 ( .INP(n34095), .ZN(n21802) );
  NAND3X0 U24770 ( .IN1(m0s3_cyc), .IN2(n34309), .IN3(n34485), .QN(n30408) );
  NAND3X0 U24771 ( .IN1(m1s3_cyc), .IN2(n34310), .IN3(n34486), .QN(n30375) );
  NAND2X0 U24772 ( .IN1(n30408), .IN2(n30375), .QN(n30353) );
  NAND2X0 U24773 ( .IN1(m3s3_cyc), .IN2(n34564), .QN(n21797) );
  NOR2X0 U24774 ( .IN1(n13738), .IN2(n21797), .QN(n30393) );
  NAND2X0 U24775 ( .IN1(m2s3_cyc), .IN2(n34595), .QN(n21798) );
  NOR2X0 U24776 ( .IN1(n13790), .IN2(n21798), .QN(n30386) );
  NOR2X0 U24777 ( .IN1(n30393), .IN2(n30386), .QN(n30344) );
  INVX0 U24778 ( .INP(n30344), .ZN(n30345) );
  NOR2X0 U24779 ( .IN1(n30353), .IN2(n30345), .QN(n21799) );
  NAND3X0 U24780 ( .IN1(m4s3_cyc), .IN2(n34236), .IN3(n34487), .QN(n30388) );
  NAND3X0 U24781 ( .IN1(m5s3_cyc), .IN2(n34361), .IN3(n34551), .QN(n30365) );
  NAND2X0 U24782 ( .IN1(n30388), .IN2(n30365), .QN(n30347) );
  NAND3X0 U24783 ( .IN1(m6s3_cyc), .IN2(n34311), .IN3(n34488), .QN(n30398) );
  NAND3X0 U24784 ( .IN1(m7s3_cyc), .IN2(n34312), .IN3(n34489), .QN(n30374) );
  NAND2X0 U24785 ( .IN1(n30398), .IN2(n30374), .QN(n30340) );
  NOR2X0 U24786 ( .IN1(n30347), .IN2(n30340), .QN(n30336) );
  NAND3X0 U24787 ( .IN1(n21799), .IN2(n30336), .IN3(\s3/next ), .QN(n34094) );
  AO221X1 U24788 ( .IN1(n21802), .IN2(n21801), .IN3(n21802), .IN4(n21800), 
        .IN5(n34094), .Q(n21803) );
  NAND2X0 U24789 ( .IN1(n34688), .IN2(n21803), .QN(n21804) );
  NOR2X0 U24790 ( .IN1(n21805), .IN2(n21804), .QN(n17593) );
  NOR2X0 U24791 ( .IN1(\s2/next ), .IN2(\s2/msel/pri_out [1]), .QN(n21812) );
  NAND3X0 U24792 ( .IN1(n13581), .IN2(m6s2_cyc), .IN3(n34576), .QN(n30312) );
  NAND2X0 U24793 ( .IN1(m7s2_cyc), .IN2(n34641), .QN(n21809) );
  NOR2X0 U24794 ( .IN1(n34478), .IN2(n21809), .QN(n30286) );
  INVX0 U24795 ( .INP(n30286), .ZN(n30283) );
  NAND2X0 U24796 ( .IN1(n30312), .IN2(n30283), .QN(n30251) );
  NAND3X0 U24797 ( .IN1(n13685), .IN2(m4s2_cyc), .IN3(n34373), .QN(n30296) );
  NAND3X0 U24798 ( .IN1(n13633), .IN2(m5s2_cyc), .IN3(n34484), .QN(n30289) );
  NAND2X0 U24799 ( .IN1(n30296), .IN2(n30289), .QN(n30252) );
  NOR2X0 U24800 ( .IN1(n30251), .IN2(n30252), .QN(n34088) );
  NAND3X0 U24801 ( .IN1(n13900), .IN2(m0s2_cyc), .IN3(n34523), .QN(n30297) );
  NAND3X0 U24802 ( .IN1(n13841), .IN2(m1s2_cyc), .IN3(n34524), .QN(n30284) );
  NAND2X0 U24803 ( .IN1(n30297), .IN2(n30284), .QN(n30247) );
  NAND2X0 U24804 ( .IN1(m3s2_cyc), .IN2(n34647), .QN(n21806) );
  NOR2X0 U24805 ( .IN1(n34479), .IN2(n21806), .QN(n30260) );
  INVX0 U24806 ( .INP(n30260), .ZN(n30280) );
  NAND3X0 U24807 ( .IN1(n13789), .IN2(m2s2_cyc), .IN3(n34563), .QN(n30314) );
  NAND2X0 U24808 ( .IN1(n30280), .IN2(n30314), .QN(n30254) );
  NOR2X0 U24809 ( .IN1(n30247), .IN2(n30254), .QN(n34089) );
  NAND3X0 U24810 ( .IN1(m0s2_cyc), .IN2(n34308), .IN3(n34523), .QN(n30073) );
  NAND3X0 U24811 ( .IN1(m1s2_cyc), .IN2(n34337), .IN3(n34524), .QN(n30051) );
  NAND2X0 U24812 ( .IN1(n30073), .IN2(n30051), .QN(n30023) );
  INVX0 U24813 ( .INP(n30023), .ZN(n30039) );
  NOR2X0 U24814 ( .IN1(n13737), .IN2(n21806), .QN(n30012) );
  NAND2X0 U24815 ( .IN1(m2s2_cyc), .IN2(n34563), .QN(n21807) );
  NOR2X0 U24816 ( .IN1(n13789), .IN2(n21807), .QN(n30087) );
  NOR2X0 U24817 ( .IN1(n30012), .IN2(n30087), .QN(n30024) );
  NAND2X0 U24818 ( .IN1(n30039), .IN2(n30024), .QN(n30017) );
  NAND3X0 U24819 ( .IN1(m5s2_cyc), .IN2(n34307), .IN3(n34484), .QN(n30061) );
  INVX0 U24820 ( .INP(n30061), .ZN(n30044) );
  AND3X1 U24821 ( .IN1(m4s2_cyc), .IN2(n34605), .IN3(n34373), .Q(n30070) );
  NOR2X0 U24822 ( .IN1(n30044), .IN2(n30070), .QN(n30038) );
  NAND2X0 U24823 ( .IN1(m6s2_cyc), .IN2(n34576), .QN(n21808) );
  NOR2X0 U24824 ( .IN1(n13581), .IN2(n21808), .QN(n30082) );
  NOR2X0 U24825 ( .IN1(n13529), .IN2(n21809), .QN(n30055) );
  NOR2X0 U24826 ( .IN1(n30082), .IN2(n30055), .QN(n30036) );
  NAND2X0 U24827 ( .IN1(n30038), .IN2(n30036), .QN(n30020) );
  NOR3X0 U24828 ( .IN1(n30017), .IN2(n30020), .IN3(n34667), .QN(n34092) );
  NAND3X0 U24829 ( .IN1(n34088), .IN2(n34089), .IN3(n34092), .QN(n21810) );
  NAND2X0 U24830 ( .IN1(n34681), .IN2(n21810), .QN(n21811) );
  NOR2X0 U24831 ( .IN1(n21812), .IN2(n21811), .QN(n17594) );
  NOR2X0 U24832 ( .IN1(\s0/next ), .IN2(\s0/msel/pri_out [0]), .QN(n21822) );
  NAND3X0 U24833 ( .IN1(n13631), .IN2(m5s0_cyc), .IN3(n34520), .QN(n29697) );
  INVX0 U24834 ( .INP(n29697), .ZN(n29664) );
  NAND3X0 U24835 ( .IN1(n13683), .IN2(m4s0_cyc), .IN3(n34519), .QN(n29647) );
  INVX0 U24836 ( .INP(n29647), .ZN(n29704) );
  NOR2X0 U24837 ( .IN1(n29664), .IN2(n29704), .QN(n29644) );
  NAND3X0 U24838 ( .IN1(n13579), .IN2(m6s0_cyc), .IN3(n34575), .QN(n29654) );
  NAND3X0 U24839 ( .IN1(n13527), .IN2(m7s0_cyc), .IN3(n34562), .QN(n29685) );
  NAND2X0 U24840 ( .IN1(n29654), .IN2(n29685), .QN(n29646) );
  INVX0 U24841 ( .INP(n29646), .ZN(n29634) );
  NAND2X0 U24842 ( .IN1(n29644), .IN2(n29634), .QN(n29640) );
  NAND3X0 U24843 ( .IN1(n13896), .IN2(m0s0_cyc), .IN3(n34572), .QN(n29695) );
  NAND3X0 U24844 ( .IN1(n13839), .IN2(m1s0_cyc), .IN3(n34573), .QN(n29686) );
  NAND2X0 U24845 ( .IN1(n29695), .IN2(n29686), .QN(n29661) );
  NAND3X0 U24846 ( .IN1(n13735), .IN2(m3s0_cyc), .IN3(n34561), .QN(n29680) );
  INVX0 U24847 ( .INP(n29680), .ZN(n29637) );
  NAND3X0 U24848 ( .IN1(n13787), .IN2(m2s0_cyc), .IN3(n34574), .QN(n29716) );
  INVX0 U24849 ( .INP(n29716), .ZN(n29688) );
  NOR2X0 U24850 ( .IN1(n29637), .IN2(n29688), .QN(n29660) );
  NAND2X0 U24851 ( .IN1(n29645), .IN2(n29660), .QN(n29635) );
  NOR2X0 U24852 ( .IN1(n29640), .IN2(n29635), .QN(n34067) );
  NAND3X0 U24853 ( .IN1(n13761), .IN2(m2s0_cyc), .IN3(n34612), .QN(n29526) );
  INVX0 U24854 ( .INP(n29526), .ZN(n29514) );
  NAND3X0 U24855 ( .IN1(n13709), .IN2(m3s0_cyc), .IN3(n34613), .QN(n29507) );
  INVX0 U24856 ( .INP(n29507), .ZN(n29520) );
  NOR2X0 U24857 ( .IN1(n29514), .IN2(n29520), .QN(n29485) );
  NAND3X0 U24858 ( .IN1(n13865), .IN2(m0s0_cyc), .IN3(n34623), .QN(n29527) );
  NAND3X0 U24859 ( .IN1(n13813), .IN2(m1s0_cyc), .IN3(n34624), .QN(n29509) );
  NAND2X0 U24860 ( .IN1(n29527), .IN2(n29509), .QN(n29487) );
  INVX0 U24861 ( .INP(n29487), .ZN(n29481) );
  NAND2X0 U24862 ( .IN1(n29485), .IN2(n29481), .QN(n29472) );
  NAND3X0 U24863 ( .IN1(n13553), .IN2(m6s0_cyc), .IN3(n34614), .QN(n29519) );
  NAND3X0 U24864 ( .IN1(n13471), .IN2(m7s0_cyc), .IN3(n34625), .QN(n29508) );
  NAND2X0 U24865 ( .IN1(n29519), .IN2(n29508), .QN(n29490) );
  INVX0 U24866 ( .INP(n29490), .ZN(n29482) );
  NAND3X0 U24867 ( .IN1(n13657), .IN2(m4s0_cyc), .IN3(n34304), .QN(n29506) );
  NAND3X0 U24868 ( .IN1(n13605), .IN2(m5s0_cyc), .IN3(n34305), .QN(n29515) );
  NAND2X0 U24869 ( .IN1(n29506), .IN2(n29515), .QN(n29486) );
  INVX0 U24870 ( .INP(n29486), .ZN(n29480) );
  NAND2X0 U24871 ( .IN1(n29482), .IN2(n29480), .QN(n29475) );
  NAND2X0 U24872 ( .IN1(m1s0_cyc), .IN2(n34573), .QN(n21813) );
  NOR2X0 U24873 ( .IN1(n13839), .IN2(n21813), .QN(n29461) );
  NAND2X0 U24874 ( .IN1(m0s0_cyc), .IN2(n34572), .QN(n21814) );
  NOR2X0 U24875 ( .IN1(n13896), .IN2(n21814), .QN(n29459) );
  NOR2X0 U24876 ( .IN1(n29461), .IN2(n29459), .QN(n29397) );
  NAND2X0 U24877 ( .IN1(m3s0_cyc), .IN2(n34561), .QN(n21815) );
  NOR2X0 U24878 ( .IN1(n13735), .IN2(n21815), .QN(n29433) );
  NAND2X0 U24879 ( .IN1(m2s0_cyc), .IN2(n34574), .QN(n21816) );
  NOR2X0 U24880 ( .IN1(n13787), .IN2(n21816), .QN(n29460) );
  NOR2X0 U24881 ( .IN1(n29433), .IN2(n29460), .QN(n29400) );
  NAND3X0 U24882 ( .IN1(m4s0_cyc), .IN2(n34304), .IN3(n34519), .QN(n29422) );
  NAND3X0 U24883 ( .IN1(m5s0_cyc), .IN2(n34305), .IN3(n34520), .QN(n29431) );
  NAND2X0 U24884 ( .IN1(n29422), .IN2(n29431), .QN(n29408) );
  NAND2X0 U24885 ( .IN1(m6s0_cyc), .IN2(n34575), .QN(n21817) );
  NOR2X0 U24886 ( .IN1(n13579), .IN2(n21817), .QN(n29436) );
  NAND2X0 U24887 ( .IN1(m7s0_cyc), .IN2(n34562), .QN(n21818) );
  NOR2X0 U24888 ( .IN1(n13527), .IN2(n21818), .QN(n29445) );
  NOR2X0 U24889 ( .IN1(n29436), .IN2(n29445), .QN(n29398) );
  INVX0 U24890 ( .INP(n29398), .ZN(n21819) );
  NOR2X0 U24891 ( .IN1(n29408), .IN2(n21819), .QN(n29394) );
  NAND4X0 U24892 ( .IN1(n29397), .IN2(n29400), .IN3(n29394), .IN4(\s0/next ), 
        .QN(n34068) );
  AO221X1 U24893 ( .IN1(n34067), .IN2(n29472), .IN3(n34067), .IN4(n29475), 
        .IN5(n34068), .Q(n21820) );
  NAND2X0 U24894 ( .IN1(n34693), .IN2(n21820), .QN(n21821) );
  NOR2X0 U24895 ( .IN1(n21822), .IN2(n21821), .QN(n17599) );
  INVX0 U24896 ( .INP(m0s0_addr[28]), .ZN(n28912) );
  INVX0 U24897 ( .INP(m0s0_addr[29]), .ZN(n28925) );
  NAND2X0 U24898 ( .IN1(n28912), .IN2(n28925), .QN(n21827) );
  INVX0 U24899 ( .INP(m0s0_addr[31]), .ZN(n28950) );
  INVX0 U24900 ( .INP(m0s0_addr[30]), .ZN(n28931) );
  NAND2X0 U24901 ( .IN1(n28950), .IN2(n28931), .QN(n21832) );
  OR2X1 U24902 ( .IN1(n21827), .IN2(n21832), .Q(n23157) );
  NAND2X0 U24903 ( .IN1(m0s0_addr[31]), .IN2(m0s0_addr[30]), .QN(n21824) );
  NAND2X0 U24904 ( .IN1(n28925), .IN2(m0s0_addr[28]), .QN(n21825) );
  NOR2X0 U24905 ( .IN1(n21824), .IN2(n21825), .QN(n29238) );
  INVX0 U24906 ( .INP(n29238), .ZN(n23131) );
  OA22X1 U24907 ( .IN1(n23157), .IN2(n22204), .IN3(n23131), .IN4(n21823), .Q(
        n21843) );
  NAND2X0 U24908 ( .IN1(n28912), .IN2(m0s0_addr[29]), .QN(n21833) );
  NAND2X0 U24909 ( .IN1(n28931), .IN2(m0s0_addr[31]), .QN(n21826) );
  OR2X1 U24910 ( .IN1(n21833), .IN2(n21826), .Q(n23161) );
  NAND2X0 U24911 ( .IN1(m0s0_addr[28]), .IN2(m0s0_addr[29]), .QN(n21829) );
  NOR2X0 U24912 ( .IN1(n21829), .IN2(n21832), .QN(n29248) );
  INVX0 U24913 ( .INP(n29248), .ZN(n23167) );
  OA22X1 U24914 ( .IN1(n23161), .IN2(n22207), .IN3(n23167), .IN4(n22206), .Q(
        n21842) );
  NOR2X0 U24915 ( .IN1(n21829), .IN2(n21826), .QN(n29240) );
  OR2X1 U24916 ( .IN1(n21824), .IN2(n21833), .Q(n23127) );
  INVX0 U24917 ( .INP(n23127), .ZN(n29237) );
  AO22X1 U24918 ( .IN1(n29240), .IN2(m0s11_data_i[0]), .IN3(n29237), .IN4(
        m0s14_data_i[0]), .Q(n21839) );
  OR2X1 U24919 ( .IN1(n21824), .IN2(n21827), .Q(n23153) );
  INVX0 U24920 ( .INP(n23153), .ZN(n29239) );
  NAND2X0 U24921 ( .IN1(m0s0_addr[30]), .IN2(n28950), .QN(n21828) );
  OR2X1 U24922 ( .IN1(n21833), .IN2(n21828), .Q(n23139) );
  INVX0 U24923 ( .INP(n23139), .ZN(n29245) );
  AO22X1 U24924 ( .IN1(n29239), .IN2(m0s12_data_i[0]), .IN3(n29245), .IN4(
        m0s6_data_i[0]), .Q(n21838) );
  NOR2X0 U24925 ( .IN1(n21827), .IN2(n21826), .QN(n29243) );
  NOR2X0 U24926 ( .IN1(n21832), .IN2(n21825), .QN(n29250) );
  AO22X1 U24927 ( .IN1(n29243), .IN2(m0s8_data_i[0]), .IN3(n29250), .IN4(
        m0s1_data_i[0]), .Q(n21837) );
  OR2X1 U24928 ( .IN1(n21828), .IN2(n21825), .Q(n23135) );
  INVX0 U24929 ( .INP(n23135), .ZN(n29246) );
  NOR2X0 U24930 ( .IN1(n21826), .IN2(n21825), .QN(n29242) );
  AO22X1 U24931 ( .IN1(n29246), .IN2(m0s5_data_i[0]), .IN3(n29242), .IN4(
        m0s9_data_i[0]), .Q(n21831) );
  NOR2X0 U24932 ( .IN1(n21827), .IN2(n21828), .QN(n29247) );
  NOR2X0 U24933 ( .IN1(n21829), .IN2(n21828), .QN(n29244) );
  AO22X1 U24934 ( .IN1(n29247), .IN2(m0s4_data_i[0]), .IN3(n29244), .IN4(
        m0s7_data_i[0]), .Q(n21830) );
  NOR2X0 U24935 ( .IN1(n21831), .IN2(n21830), .QN(n21835) );
  NOR2X0 U24936 ( .IN1(n21833), .IN2(n21832), .QN(n29249) );
  NAND2X0 U24937 ( .IN1(n29249), .IN2(m0s2_data_i[0]), .QN(n21834) );
  NAND2X0 U24938 ( .IN1(n21835), .IN2(n21834), .QN(n21836) );
  NOR4X0 U24939 ( .IN1(n21839), .IN2(n21838), .IN3(n21837), .IN4(n21836), .QN(
        n21841) );
  INVX0 U24940 ( .INP(n22021), .ZN(n29236) );
  NAND2X0 U24941 ( .IN1(n29236), .IN2(n22218), .QN(n21840) );
  NAND4X0 U24942 ( .IN1(n21843), .IN2(n21842), .IN3(n21841), .IN4(n21840), 
        .QN(m0_data_o[0]) );
  INVX0 U24943 ( .INP(n23161), .ZN(n29241) );
  AO22X1 U24944 ( .IN1(n29241), .IN2(m0s10_data_i[1]), .IN3(n29249), .IN4(
        m0s2_data_i[1]), .Q(n21846) );
  INVX0 U24945 ( .INP(n29240), .ZN(n23149) );
  AO22X1 U24946 ( .IN1(n29240), .IN2(m0s11_data_i[1]), .IN3(n29243), .IN4(
        m0s8_data_i[1]), .Q(n21845) );
  INVX0 U24947 ( .INP(n23157), .ZN(n29252) );
  AO22X1 U24948 ( .IN1(n29252), .IN2(m0s0_data_i[1]), .IN3(n29247), .IN4(
        m0s4_data_i[1]), .Q(n21844) );
  NOR3X0 U24949 ( .IN1(n21846), .IN2(n21845), .IN3(n21844), .QN(n21854) );
  AO22X1 U24950 ( .IN1(n29239), .IN2(m0s12_data_i[1]), .IN3(n29237), .IN4(
        m0s14_data_i[1]), .Q(n21850) );
  AO22X1 U24951 ( .IN1(n29248), .IN2(m0s3_data_i[1]), .IN3(n29246), .IN4(
        m0s5_data_i[1]), .Q(n21849) );
  AO22X1 U24952 ( .IN1(n29245), .IN2(m0s6_data_i[1]), .IN3(n29238), .IN4(
        m0s13_data_i[1]), .Q(n21848) );
  AO22X1 U24953 ( .IN1(n29250), .IN2(m0s1_data_i[1]), .IN3(n29244), .IN4(
        m0s7_data_i[1]), .Q(n21847) );
  NOR4X0 U24954 ( .IN1(n21850), .IN2(n21849), .IN3(n21848), .IN4(n21847), .QN(
        n21853) );
  NAND2X0 U24955 ( .IN1(n29236), .IN2(n22235), .QN(n21852) );
  NAND2X0 U24956 ( .IN1(n29242), .IN2(m0s9_data_i[1]), .QN(n21851) );
  NAND4X0 U24957 ( .IN1(n21854), .IN2(n21853), .IN3(n21852), .IN4(n21851), 
        .QN(m0_data_o[1]) );
  AO22X1 U24958 ( .IN1(n29245), .IN2(m0s6_data_i[2]), .IN3(n29240), .IN4(
        m0s11_data_i[2]), .Q(n21857) );
  AO22X1 U24959 ( .IN1(n29250), .IN2(m0s1_data_i[2]), .IN3(n29246), .IN4(
        m0s5_data_i[2]), .Q(n21856) );
  AO22X1 U24960 ( .IN1(n29237), .IN2(m0s14_data_i[2]), .IN3(n29249), .IN4(
        m0s2_data_i[2]), .Q(n21855) );
  NOR3X0 U24961 ( .IN1(n21857), .IN2(n21856), .IN3(n21855), .QN(n21865) );
  AO22X1 U24962 ( .IN1(n29248), .IN2(m0s3_data_i[2]), .IN3(n29244), .IN4(
        m0s7_data_i[2]), .Q(n21861) );
  AO22X1 U24963 ( .IN1(n29239), .IN2(m0s12_data_i[2]), .IN3(n29242), .IN4(
        m0s9_data_i[2]), .Q(n21860) );
  AO22X1 U24964 ( .IN1(n29241), .IN2(m0s10_data_i[2]), .IN3(n29238), .IN4(
        m0s13_data_i[2]), .Q(n21859) );
  AO22X1 U24965 ( .IN1(n29243), .IN2(m0s8_data_i[2]), .IN3(n29247), .IN4(
        m0s4_data_i[2]), .Q(n21858) );
  NOR4X0 U24966 ( .IN1(n21861), .IN2(n21860), .IN3(n21859), .IN4(n21858), .QN(
        n21864) );
  NAND2X0 U24967 ( .IN1(n29236), .IN2(n22247), .QN(n21863) );
  NAND2X0 U24968 ( .IN1(n29252), .IN2(m0s0_data_i[2]), .QN(n21862) );
  NAND4X0 U24969 ( .IN1(n21865), .IN2(n21864), .IN3(n21863), .IN4(n21862), 
        .QN(m0_data_o[2]) );
  AO22X1 U24970 ( .IN1(n29242), .IN2(m0s9_data_i[3]), .IN3(n29247), .IN4(
        m0s4_data_i[3]), .Q(n21868) );
  AO22X1 U24971 ( .IN1(n29252), .IN2(m0s0_data_i[3]), .IN3(n29243), .IN4(
        m0s8_data_i[3]), .Q(n21867) );
  AO22X1 U24972 ( .IN1(n29237), .IN2(m0s14_data_i[3]), .IN3(n29241), .IN4(
        m0s10_data_i[3]), .Q(n21866) );
  NOR3X0 U24973 ( .IN1(n21868), .IN2(n21867), .IN3(n21866), .QN(n21876) );
  AO22X1 U24974 ( .IN1(n29239), .IN2(m0s12_data_i[3]), .IN3(n29248), .IN4(
        m0s3_data_i[3]), .Q(n21872) );
  AO22X1 U24975 ( .IN1(n29240), .IN2(m0s11_data_i[3]), .IN3(n29244), .IN4(
        m0s7_data_i[3]), .Q(n21871) );
  AO22X1 U24976 ( .IN1(n29245), .IN2(m0s6_data_i[3]), .IN3(n29249), .IN4(
        m0s2_data_i[3]), .Q(n21870) );
  AO22X1 U24977 ( .IN1(n29250), .IN2(m0s1_data_i[3]), .IN3(n29246), .IN4(
        m0s5_data_i[3]), .Q(n21869) );
  NOR4X0 U24978 ( .IN1(n21872), .IN2(n21871), .IN3(n21870), .IN4(n21869), .QN(
        n21875) );
  NAND2X0 U24979 ( .IN1(n29236), .IN2(n22646), .QN(n21874) );
  NAND2X0 U24980 ( .IN1(n29238), .IN2(m0s13_data_i[3]), .QN(n21873) );
  NAND4X0 U24981 ( .IN1(n21876), .IN2(n21875), .IN3(n21874), .IN4(n21873), 
        .QN(m0_data_o[3]) );
  AO22X1 U24982 ( .IN1(n29243), .IN2(m0s8_data_i[4]), .IN3(n29242), .IN4(
        m0s9_data_i[4]), .Q(n21879) );
  AO22X1 U24983 ( .IN1(n29240), .IN2(m0s11_data_i[4]), .IN3(n29241), .IN4(
        m0s10_data_i[4]), .Q(n21878) );
  AO22X1 U24984 ( .IN1(n29237), .IN2(m0s14_data_i[4]), .IN3(n29252), .IN4(
        m0s0_data_i[4]), .Q(n21877) );
  NOR3X0 U24985 ( .IN1(n21879), .IN2(n21878), .IN3(n21877), .QN(n21887) );
  AO22X1 U24986 ( .IN1(n29239), .IN2(m0s12_data_i[4]), .IN3(n29250), .IN4(
        m0s1_data_i[4]), .Q(n21883) );
  AO22X1 U24987 ( .IN1(n29248), .IN2(m0s3_data_i[4]), .IN3(n29246), .IN4(
        m0s5_data_i[4]), .Q(n21882) );
  AO22X1 U24988 ( .IN1(n29247), .IN2(m0s4_data_i[4]), .IN3(n29244), .IN4(
        m0s7_data_i[4]), .Q(n21881) );
  AO22X1 U24989 ( .IN1(n29245), .IN2(m0s6_data_i[4]), .IN3(n29249), .IN4(
        m0s2_data_i[4]), .Q(n21880) );
  NOR4X0 U24990 ( .IN1(n21883), .IN2(n21882), .IN3(n21881), .IN4(n21880), .QN(
        n21886) );
  NAND2X0 U24991 ( .IN1(n29236), .IN2(n22663), .QN(n21885) );
  NAND2X0 U24992 ( .IN1(n29238), .IN2(m0s13_data_i[4]), .QN(n21884) );
  NAND4X0 U24993 ( .IN1(n21887), .IN2(n21886), .IN3(n21885), .IN4(n21884), 
        .QN(m0_data_o[4]) );
  AO22X1 U24994 ( .IN1(n29239), .IN2(m0s12_data_i[5]), .IN3(n29246), .IN4(
        m0s5_data_i[5]), .Q(n21890) );
  AO22X1 U24995 ( .IN1(n29243), .IN2(m0s8_data_i[5]), .IN3(n29242), .IN4(
        m0s9_data_i[5]), .Q(n21889) );
  AO22X1 U24996 ( .IN1(n29240), .IN2(m0s11_data_i[5]), .IN3(n29244), .IN4(
        m0s7_data_i[5]), .Q(n21888) );
  NOR3X0 U24997 ( .IN1(n21890), .IN2(n21889), .IN3(n21888), .QN(n21898) );
  AO22X1 U24998 ( .IN1(n29252), .IN2(m0s0_data_i[5]), .IN3(n29249), .IN4(
        m0s2_data_i[5]), .Q(n21894) );
  AO22X1 U24999 ( .IN1(n29245), .IN2(m0s6_data_i[5]), .IN3(n29241), .IN4(
        m0s10_data_i[5]), .Q(n21893) );
  AO22X1 U25000 ( .IN1(n29237), .IN2(m0s14_data_i[5]), .IN3(n29238), .IN4(
        m0s13_data_i[5]), .Q(n21892) );
  AO22X1 U25001 ( .IN1(n29248), .IN2(m0s3_data_i[5]), .IN3(n29247), .IN4(
        m0s4_data_i[5]), .Q(n21891) );
  NOR4X0 U25002 ( .IN1(n21894), .IN2(n21893), .IN3(n21892), .IN4(n21891), .QN(
        n21897) );
  NAND2X0 U25003 ( .IN1(n29236), .IN2(n22680), .QN(n21896) );
  NAND2X0 U25004 ( .IN1(n29250), .IN2(m0s1_data_i[5]), .QN(n21895) );
  NAND4X0 U25005 ( .IN1(n21898), .IN2(n21897), .IN3(n21896), .IN4(n21895), 
        .QN(m0_data_o[5]) );
  AO22X1 U25006 ( .IN1(n29252), .IN2(m0s0_data_i[6]), .IN3(n29247), .IN4(
        m0s4_data_i[6]), .Q(n21901) );
  AO22X1 U25007 ( .IN1(n29237), .IN2(m0s14_data_i[6]), .IN3(n29248), .IN4(
        m0s3_data_i[6]), .Q(n21900) );
  AO22X1 U25008 ( .IN1(n29240), .IN2(m0s11_data_i[6]), .IN3(n29250), .IN4(
        m0s1_data_i[6]), .Q(n21899) );
  NOR3X0 U25009 ( .IN1(n21901), .IN2(n21900), .IN3(n21899), .QN(n21909) );
  AO22X1 U25010 ( .IN1(n29243), .IN2(m0s8_data_i[6]), .IN3(n29244), .IN4(
        m0s7_data_i[6]), .Q(n21905) );
  AO22X1 U25011 ( .IN1(n29239), .IN2(m0s12_data_i[6]), .IN3(n29246), .IN4(
        m0s5_data_i[6]), .Q(n21904) );
  AO22X1 U25012 ( .IN1(n29245), .IN2(m0s6_data_i[6]), .IN3(n29249), .IN4(
        m0s2_data_i[6]), .Q(n21903) );
  AO22X1 U25013 ( .IN1(n29241), .IN2(m0s10_data_i[6]), .IN3(n29242), .IN4(
        m0s9_data_i[6]), .Q(n21902) );
  NOR4X0 U25014 ( .IN1(n21905), .IN2(n21904), .IN3(n21903), .IN4(n21902), .QN(
        n21908) );
  NAND2X0 U25015 ( .IN1(n29236), .IN2(n22697), .QN(n21907) );
  NAND2X0 U25016 ( .IN1(n29238), .IN2(m0s13_data_i[6]), .QN(n21906) );
  NAND4X0 U25017 ( .IN1(n21909), .IN2(n21908), .IN3(n21907), .IN4(n21906), 
        .QN(m0_data_o[6]) );
  AO22X1 U25018 ( .IN1(n29240), .IN2(m0s11_data_i[7]), .IN3(n29237), .IN4(
        m0s14_data_i[7]), .Q(n21912) );
  AO22X1 U25019 ( .IN1(n29241), .IN2(m0s10_data_i[7]), .IN3(n29248), .IN4(
        m0s3_data_i[7]), .Q(n21911) );
  AO22X1 U25020 ( .IN1(n29238), .IN2(m0s13_data_i[7]), .IN3(n29249), .IN4(
        m0s2_data_i[7]), .Q(n21910) );
  NOR3X0 U25021 ( .IN1(n21912), .IN2(n21911), .IN3(n21910), .QN(n21920) );
  AO22X1 U25022 ( .IN1(n29239), .IN2(m0s12_data_i[7]), .IN3(n29242), .IN4(
        m0s9_data_i[7]), .Q(n21916) );
  AO22X1 U25023 ( .IN1(n29246), .IN2(m0s5_data_i[7]), .IN3(n29247), .IN4(
        m0s4_data_i[7]), .Q(n21915) );
  AO22X1 U25024 ( .IN1(n29243), .IN2(m0s8_data_i[7]), .IN3(n29250), .IN4(
        m0s1_data_i[7]), .Q(n21914) );
  AO22X1 U25025 ( .IN1(n29252), .IN2(m0s0_data_i[7]), .IN3(n29244), .IN4(
        m0s7_data_i[7]), .Q(n21913) );
  NOR4X0 U25026 ( .IN1(n21916), .IN2(n21915), .IN3(n21914), .IN4(n21913), .QN(
        n21919) );
  NAND2X0 U25027 ( .IN1(n29236), .IN2(n22714), .QN(n21918) );
  NAND2X0 U25028 ( .IN1(n29245), .IN2(m0s6_data_i[7]), .QN(n21917) );
  NAND4X0 U25029 ( .IN1(n21920), .IN2(n21919), .IN3(n21918), .IN4(n21917), 
        .QN(m0_data_o[7]) );
  AO22X1 U25030 ( .IN1(n29238), .IN2(m0s13_data_i[8]), .IN3(n29243), .IN4(
        m0s8_data_i[8]), .Q(n21923) );
  AO22X1 U25031 ( .IN1(n29248), .IN2(m0s3_data_i[8]), .IN3(n29249), .IN4(
        m0s2_data_i[8]), .Q(n21922) );
  AO22X1 U25032 ( .IN1(n29237), .IN2(m0s14_data_i[8]), .IN3(n29242), .IN4(
        m0s9_data_i[8]), .Q(n21921) );
  NOR3X0 U25033 ( .IN1(n21923), .IN2(n21922), .IN3(n21921), .QN(n21931) );
  AO22X1 U25034 ( .IN1(n29246), .IN2(m0s5_data_i[8]), .IN3(n29244), .IN4(
        m0s7_data_i[8]), .Q(n21927) );
  AO22X1 U25035 ( .IN1(n29239), .IN2(m0s12_data_i[8]), .IN3(n29240), .IN4(
        m0s11_data_i[8]), .Q(n21926) );
  AO22X1 U25036 ( .IN1(n29245), .IN2(m0s6_data_i[8]), .IN3(n29250), .IN4(
        m0s1_data_i[8]), .Q(n21925) );
  AO22X1 U25037 ( .IN1(n29241), .IN2(m0s10_data_i[8]), .IN3(n29247), .IN4(
        m0s4_data_i[8]), .Q(n21924) );
  NOR4X0 U25038 ( .IN1(n21927), .IN2(n21926), .IN3(n21925), .IN4(n21924), .QN(
        n21930) );
  NAND2X0 U25039 ( .IN1(n29236), .IN2(n22731), .QN(n21929) );
  NAND2X0 U25040 ( .IN1(n29252), .IN2(m0s0_data_i[8]), .QN(n21928) );
  NAND4X0 U25041 ( .IN1(n21931), .IN2(n21930), .IN3(n21929), .IN4(n21928), 
        .QN(m0_data_o[8]) );
  AO22X1 U25042 ( .IN1(n29246), .IN2(m0s5_data_i[9]), .IN3(n29247), .IN4(
        m0s4_data_i[9]), .Q(n21934) );
  AO22X1 U25043 ( .IN1(n29252), .IN2(m0s0_data_i[9]), .IN3(n29244), .IN4(
        m0s7_data_i[9]), .Q(n21933) );
  AO22X1 U25044 ( .IN1(n29237), .IN2(m0s14_data_i[9]), .IN3(n29250), .IN4(
        m0s1_data_i[9]), .Q(n21932) );
  NOR3X0 U25045 ( .IN1(n21934), .IN2(n21933), .IN3(n21932), .QN(n21942) );
  AO22X1 U25046 ( .IN1(n29241), .IN2(m0s10_data_i[9]), .IN3(n29249), .IN4(
        m0s2_data_i[9]), .Q(n21938) );
  AO22X1 U25047 ( .IN1(n29248), .IN2(m0s3_data_i[9]), .IN3(n29242), .IN4(
        m0s9_data_i[9]), .Q(n21937) );
  AO22X1 U25048 ( .IN1(n29238), .IN2(m0s13_data_i[9]), .IN3(n29243), .IN4(
        m0s8_data_i[9]), .Q(n21936) );
  AO22X1 U25049 ( .IN1(n29239), .IN2(m0s12_data_i[9]), .IN3(n29245), .IN4(
        m0s6_data_i[9]), .Q(n21935) );
  NOR4X0 U25050 ( .IN1(n21938), .IN2(n21937), .IN3(n21936), .IN4(n21935), .QN(
        n21941) );
  NAND2X0 U25051 ( .IN1(n29236), .IN2(n22993), .QN(n21940) );
  NAND2X0 U25052 ( .IN1(n29240), .IN2(m0s11_data_i[9]), .QN(n21939) );
  NAND4X0 U25053 ( .IN1(n21942), .IN2(n21941), .IN3(n21940), .IN4(n21939), 
        .QN(m0_data_o[9]) );
  AO22X1 U25054 ( .IN1(n29237), .IN2(m0s14_data_i[10]), .IN3(n29243), .IN4(
        m0s8_data_i[10]), .Q(n21945) );
  AO22X1 U25055 ( .IN1(n29252), .IN2(m0s0_data_i[10]), .IN3(n29246), .IN4(
        m0s5_data_i[10]), .Q(n21944) );
  AO22X1 U25056 ( .IN1(n29241), .IN2(m0s10_data_i[10]), .IN3(n29249), .IN4(
        m0s2_data_i[10]), .Q(n21943) );
  NOR3X0 U25057 ( .IN1(n21945), .IN2(n21944), .IN3(n21943), .QN(n21953) );
  AO22X1 U25058 ( .IN1(n29240), .IN2(m0s11_data_i[10]), .IN3(n29244), .IN4(
        m0s7_data_i[10]), .Q(n21949) );
  AO22X1 U25059 ( .IN1(n29238), .IN2(m0s13_data_i[10]), .IN3(n29242), .IN4(
        m0s9_data_i[10]), .Q(n21948) );
  AO22X1 U25060 ( .IN1(n29248), .IN2(m0s3_data_i[10]), .IN3(n29250), .IN4(
        m0s1_data_i[10]), .Q(n21947) );
  AO22X1 U25061 ( .IN1(n29239), .IN2(m0s12_data_i[10]), .IN3(n29245), .IN4(
        m0s6_data_i[10]), .Q(n21946) );
  NOR4X0 U25062 ( .IN1(n21949), .IN2(n21948), .IN3(n21947), .IN4(n21946), .QN(
        n21952) );
  NAND2X0 U25063 ( .IN1(n29236), .IN2(n22763), .QN(n21951) );
  NAND2X0 U25064 ( .IN1(n29247), .IN2(m0s4_data_i[10]), .QN(n21950) );
  NAND4X0 U25065 ( .IN1(n21953), .IN2(n21952), .IN3(n21951), .IN4(n21950), 
        .QN(m0_data_o[10]) );
  AO22X1 U25066 ( .IN1(n29252), .IN2(m0s0_data_i[11]), .IN3(n29244), .IN4(
        m0s7_data_i[11]), .Q(n21956) );
  AO22X1 U25067 ( .IN1(n29241), .IN2(m0s10_data_i[11]), .IN3(n29247), .IN4(
        m0s4_data_i[11]), .Q(n21955) );
  AO22X1 U25068 ( .IN1(n29243), .IN2(m0s8_data_i[11]), .IN3(n29246), .IN4(
        m0s5_data_i[11]), .Q(n21954) );
  NOR3X0 U25069 ( .IN1(n21956), .IN2(n21955), .IN3(n21954), .QN(n21964) );
  AO22X1 U25070 ( .IN1(n29245), .IN2(m0s6_data_i[11]), .IN3(n29250), .IN4(
        m0s1_data_i[11]), .Q(n21960) );
  AO22X1 U25071 ( .IN1(n29239), .IN2(m0s12_data_i[11]), .IN3(n29238), .IN4(
        m0s13_data_i[11]), .Q(n21959) );
  AO22X1 U25072 ( .IN1(n29248), .IN2(m0s3_data_i[11]), .IN3(n29249), .IN4(
        m0s2_data_i[11]), .Q(n21958) );
  AO22X1 U25073 ( .IN1(n29237), .IN2(m0s14_data_i[11]), .IN3(n29242), .IN4(
        m0s9_data_i[11]), .Q(n21957) );
  NOR4X0 U25074 ( .IN1(n21960), .IN2(n21959), .IN3(n21958), .IN4(n21957), .QN(
        n21963) );
  NAND2X0 U25075 ( .IN1(n29236), .IN2(n23013), .QN(n21962) );
  NAND2X0 U25076 ( .IN1(n29240), .IN2(m0s11_data_i[11]), .QN(n21961) );
  NAND4X0 U25077 ( .IN1(n21964), .IN2(n21963), .IN3(n21962), .IN4(n21961), 
        .QN(m0_data_o[11]) );
  AO22X1 U25078 ( .IN1(n29239), .IN2(m0s12_data_i[12]), .IN3(n29240), .IN4(
        m0s11_data_i[12]), .Q(n21967) );
  AO22X1 U25079 ( .IN1(n29238), .IN2(m0s13_data_i[12]), .IN3(n29247), .IN4(
        m0s4_data_i[12]), .Q(n21966) );
  AO22X1 U25080 ( .IN1(n29248), .IN2(m0s3_data_i[12]), .IN3(n29246), .IN4(
        m0s5_data_i[12]), .Q(n21965) );
  NOR3X0 U25081 ( .IN1(n21967), .IN2(n21966), .IN3(n21965), .QN(n21975) );
  AO22X1 U25082 ( .IN1(n29237), .IN2(m0s14_data_i[12]), .IN3(n29249), .IN4(
        m0s2_data_i[12]), .Q(n21971) );
  AO22X1 U25083 ( .IN1(n29241), .IN2(m0s10_data_i[12]), .IN3(n29243), .IN4(
        m0s8_data_i[12]), .Q(n21970) );
  AO22X1 U25084 ( .IN1(n29245), .IN2(m0s6_data_i[12]), .IN3(n29252), .IN4(
        m0s0_data_i[12]), .Q(n21969) );
  AO22X1 U25085 ( .IN1(n29242), .IN2(m0s9_data_i[12]), .IN3(n29244), .IN4(
        m0s7_data_i[12]), .Q(n21968) );
  NOR4X0 U25086 ( .IN1(n21971), .IN2(n21970), .IN3(n21969), .IN4(n21968), .QN(
        n21974) );
  NAND2X0 U25087 ( .IN1(n29236), .IN2(n23034), .QN(n21973) );
  NAND2X0 U25088 ( .IN1(n29250), .IN2(m0s1_data_i[12]), .QN(n21972) );
  NAND4X0 U25089 ( .IN1(n21975), .IN2(n21974), .IN3(n21973), .IN4(n21972), 
        .QN(m0_data_o[12]) );
  AO22X1 U25090 ( .IN1(n29239), .IN2(m0s12_data_i[13]), .IN3(n29246), .IN4(
        m0s5_data_i[13]), .Q(n21978) );
  AO22X1 U25091 ( .IN1(n29248), .IN2(m0s3_data_i[13]), .IN3(n29250), .IN4(
        m0s1_data_i[13]), .Q(n21977) );
  AO22X1 U25092 ( .IN1(n29237), .IN2(m0s14_data_i[13]), .IN3(n29242), .IN4(
        m0s9_data_i[13]), .Q(n21976) );
  NOR3X0 U25093 ( .IN1(n21978), .IN2(n21977), .IN3(n21976), .QN(n21986) );
  AO22X1 U25094 ( .IN1(n29252), .IN2(m0s0_data_i[13]), .IN3(n29238), .IN4(
        m0s13_data_i[13]), .Q(n21982) );
  AO22X1 U25095 ( .IN1(n29245), .IN2(m0s6_data_i[13]), .IN3(n29244), .IN4(
        m0s7_data_i[13]), .Q(n21981) );
  AO22X1 U25096 ( .IN1(n29240), .IN2(m0s11_data_i[13]), .IN3(n29247), .IN4(
        m0s4_data_i[13]), .Q(n21980) );
  AO22X1 U25097 ( .IN1(n29241), .IN2(m0s10_data_i[13]), .IN3(n29243), .IN4(
        m0s8_data_i[13]), .Q(n21979) );
  NOR4X0 U25098 ( .IN1(n21982), .IN2(n21981), .IN3(n21980), .IN4(n21979), .QN(
        n21985) );
  NAND2X0 U25099 ( .IN1(n29236), .IN2(n23053), .QN(n21984) );
  NAND2X0 U25100 ( .IN1(n29249), .IN2(m0s2_data_i[13]), .QN(n21983) );
  NAND4X0 U25101 ( .IN1(n21986), .IN2(n21985), .IN3(n21984), .IN4(n21983), 
        .QN(m0_data_o[13]) );
  AO22X1 U25102 ( .IN1(n29237), .IN2(m0s14_data_i[14]), .IN3(n29247), .IN4(
        m0s4_data_i[14]), .Q(n21989) );
  AO22X1 U25103 ( .IN1(n29240), .IN2(m0s11_data_i[14]), .IN3(n29238), .IN4(
        m0s13_data_i[14]), .Q(n21988) );
  AO22X1 U25104 ( .IN1(n29239), .IN2(m0s12_data_i[14]), .IN3(n29246), .IN4(
        m0s5_data_i[14]), .Q(n21987) );
  NOR3X0 U25105 ( .IN1(n21989), .IN2(n21988), .IN3(n21987), .QN(n21997) );
  AO22X1 U25106 ( .IN1(n29243), .IN2(m0s8_data_i[14]), .IN3(n29250), .IN4(
        m0s1_data_i[14]), .Q(n21993) );
  AO22X1 U25107 ( .IN1(n29245), .IN2(m0s6_data_i[14]), .IN3(n29252), .IN4(
        m0s0_data_i[14]), .Q(n21992) );
  AO22X1 U25108 ( .IN1(n29249), .IN2(m0s2_data_i[14]), .IN3(n29244), .IN4(
        m0s7_data_i[14]), .Q(n21991) );
  AO22X1 U25109 ( .IN1(n29241), .IN2(m0s10_data_i[14]), .IN3(n29248), .IN4(
        m0s3_data_i[14]), .Q(n21990) );
  NOR4X0 U25110 ( .IN1(n21993), .IN2(n21992), .IN3(n21991), .IN4(n21990), .QN(
        n21996) );
  NAND2X0 U25111 ( .IN1(n29236), .IN2(n23078), .QN(n21995) );
  NAND2X0 U25112 ( .IN1(n29242), .IN2(m0s9_data_i[14]), .QN(n21994) );
  NAND4X0 U25113 ( .IN1(n21997), .IN2(n21996), .IN3(n21995), .IN4(n21994), 
        .QN(m0_data_o[14]) );
  AO22X1 U25114 ( .IN1(n29241), .IN2(m0s10_data_i[15]), .IN3(n29252), .IN4(
        m0s0_data_i[15]), .Q(n22000) );
  AO22X1 U25115 ( .IN1(n29239), .IN2(m0s12_data_i[15]), .IN3(n29246), .IN4(
        m0s5_data_i[15]), .Q(n21999) );
  AO22X1 U25116 ( .IN1(n29238), .IN2(m0s13_data_i[15]), .IN3(n29247), .IN4(
        m0s4_data_i[15]), .Q(n21998) );
  NOR3X0 U25117 ( .IN1(n22000), .IN2(n21999), .IN3(n21998), .QN(n22008) );
  AO22X1 U25118 ( .IN1(n29249), .IN2(m0s2_data_i[15]), .IN3(n29244), .IN4(
        m0s7_data_i[15]), .Q(n22004) );
  AO22X1 U25119 ( .IN1(n29237), .IN2(m0s14_data_i[15]), .IN3(n29248), .IN4(
        m0s3_data_i[15]), .Q(n22003) );
  AO22X1 U25120 ( .IN1(n29240), .IN2(m0s11_data_i[15]), .IN3(n29250), .IN4(
        m0s1_data_i[15]), .Q(n22002) );
  AO22X1 U25121 ( .IN1(n29245), .IN2(m0s6_data_i[15]), .IN3(n29242), .IN4(
        m0s9_data_i[15]), .Q(n22001) );
  NOR4X0 U25122 ( .IN1(n22004), .IN2(n22003), .IN3(n22002), .IN4(n22001), .QN(
        n22007) );
  NAND2X0 U25123 ( .IN1(n29236), .IN2(n23103), .QN(n22006) );
  NAND2X0 U25124 ( .IN1(n29243), .IN2(m0s8_data_i[15]), .QN(n22005) );
  NAND4X0 U25125 ( .IN1(n22008), .IN2(n22007), .IN3(n22006), .IN4(n22005), 
        .QN(m0_data_o[15]) );
  OA22X1 U25126 ( .IN1(n23131), .IN2(n22010), .IN3(n23135), .IN4(n22009), .Q(
        n22025) );
  OA22X1 U25127 ( .IN1(n23153), .IN2(n22012), .IN3(n23149), .IN4(n22011), .Q(
        n22024) );
  AO22X1 U25128 ( .IN1(n29249), .IN2(m0s2_data_i[16]), .IN3(n29244), .IN4(
        m0s7_data_i[16]), .Q(n22020) );
  AO22X1 U25129 ( .IN1(n29237), .IN2(m0s14_data_i[16]), .IN3(n29248), .IN4(
        m0s3_data_i[16]), .Q(n22019) );
  AO22X1 U25130 ( .IN1(n29250), .IN2(m0s1_data_i[16]), .IN3(n29247), .IN4(
        m0s4_data_i[16]), .Q(n22018) );
  AO22X1 U25131 ( .IN1(n29252), .IN2(m0s0_data_i[16]), .IN3(n29243), .IN4(
        m0s8_data_i[16]), .Q(n22014) );
  AO22X1 U25132 ( .IN1(n29241), .IN2(m0s10_data_i[16]), .IN3(n29242), .IN4(
        m0s9_data_i[16]), .Q(n22013) );
  NOR2X0 U25133 ( .IN1(n22014), .IN2(n22013), .QN(n22016) );
  NAND2X0 U25134 ( .IN1(n29245), .IN2(m0s6_data_i[16]), .QN(n22015) );
  NAND2X0 U25135 ( .IN1(n22016), .IN2(n22015), .QN(n22017) );
  NOR4X0 U25136 ( .IN1(n22020), .IN2(n22019), .IN3(n22018), .IN4(n22017), .QN(
        n22023) );
  NOR2X0 U25137 ( .IN1(n23501), .IN2(n22021), .QN(n22198) );
  NAND2X0 U25138 ( .IN1(s15_data_i[16]), .IN2(n22198), .QN(n22022) );
  NAND4X0 U25139 ( .IN1(n22025), .IN2(n22024), .IN3(n22023), .IN4(n22022), 
        .QN(m0_data_o[16]) );
  AO22X1 U25140 ( .IN1(n29252), .IN2(m0s0_data_i[17]), .IN3(n29243), .IN4(
        m0s8_data_i[17]), .Q(n22028) );
  AO22X1 U25141 ( .IN1(n29241), .IN2(m0s10_data_i[17]), .IN3(n29246), .IN4(
        m0s5_data_i[17]), .Q(n22027) );
  AO22X1 U25142 ( .IN1(n29245), .IN2(m0s6_data_i[17]), .IN3(n29240), .IN4(
        m0s11_data_i[17]), .Q(n22026) );
  NOR3X0 U25143 ( .IN1(n22028), .IN2(n22027), .IN3(n22026), .QN(n22036) );
  AO22X1 U25144 ( .IN1(n29237), .IN2(m0s14_data_i[17]), .IN3(n29242), .IN4(
        m0s9_data_i[17]), .Q(n22032) );
  AO22X1 U25145 ( .IN1(n29239), .IN2(m0s12_data_i[17]), .IN3(n29244), .IN4(
        m0s7_data_i[17]), .Q(n22031) );
  AO22X1 U25146 ( .IN1(n29248), .IN2(m0s3_data_i[17]), .IN3(n29250), .IN4(
        m0s1_data_i[17]), .Q(n22030) );
  AO22X1 U25147 ( .IN1(n29249), .IN2(m0s2_data_i[17]), .IN3(n29247), .IN4(
        m0s4_data_i[17]), .Q(n22029) );
  NOR4X0 U25148 ( .IN1(n22032), .IN2(n22031), .IN3(n22030), .IN4(n22029), .QN(
        n22035) );
  NAND2X0 U25149 ( .IN1(n22198), .IN2(s15_data_i[17]), .QN(n22034) );
  NAND2X0 U25150 ( .IN1(n29238), .IN2(m0s13_data_i[17]), .QN(n22033) );
  NAND4X0 U25151 ( .IN1(n22036), .IN2(n22035), .IN3(n22034), .IN4(n22033), 
        .QN(m0_data_o[17]) );
  AOI22X1 U25152 ( .IN1(n29246), .IN2(m0s5_data_i[18]), .IN3(n29244), .IN4(
        m0s7_data_i[18]), .QN(n22049) );
  INVX0 U25153 ( .INP(n29250), .ZN(n22178) );
  OA22X1 U25154 ( .IN1(n23153), .IN2(n22410), .IN3(n22178), .IN4(n22037), .Q(
        n22048) );
  AO22X1 U25155 ( .IN1(n29242), .IN2(m0s9_data_i[18]), .IN3(n29247), .IN4(
        m0s4_data_i[18]), .Q(n22045) );
  AO22X1 U25156 ( .IN1(n29245), .IN2(m0s6_data_i[18]), .IN3(n29237), .IN4(
        m0s14_data_i[18]), .Q(n22044) );
  AO22X1 U25157 ( .IN1(n29248), .IN2(m0s3_data_i[18]), .IN3(n29238), .IN4(
        m0s13_data_i[18]), .Q(n22043) );
  AO22X1 U25158 ( .IN1(n29241), .IN2(m0s10_data_i[18]), .IN3(n29249), .IN4(
        m0s2_data_i[18]), .Q(n22039) );
  AO22X1 U25159 ( .IN1(n29240), .IN2(m0s11_data_i[18]), .IN3(n29243), .IN4(
        m0s8_data_i[18]), .Q(n22038) );
  NOR2X0 U25160 ( .IN1(n22039), .IN2(n22038), .QN(n22041) );
  NAND2X0 U25161 ( .IN1(n29252), .IN2(m0s0_data_i[18]), .QN(n22040) );
  NAND2X0 U25162 ( .IN1(n22041), .IN2(n22040), .QN(n22042) );
  NOR4X0 U25163 ( .IN1(n22045), .IN2(n22044), .IN3(n22043), .IN4(n22042), .QN(
        n22047) );
  NAND2X0 U25164 ( .IN1(n22198), .IN2(s15_data_i[18]), .QN(n22046) );
  NAND4X0 U25165 ( .IN1(n22049), .IN2(n22048), .IN3(n22047), .IN4(n22046), 
        .QN(m0_data_o[18]) );
  OA22X1 U25166 ( .IN1(n23153), .IN2(n22434), .IN3(n23167), .IN4(n22431), .Q(
        n22062) );
  OA22X1 U25167 ( .IN1(n23157), .IN2(n22433), .IN3(n23135), .IN4(n22050), .Q(
        n22061) );
  AO22X1 U25168 ( .IN1(n29242), .IN2(m0s9_data_i[19]), .IN3(n29244), .IN4(
        m0s7_data_i[19]), .Q(n22058) );
  AO22X1 U25169 ( .IN1(n29237), .IN2(m0s14_data_i[19]), .IN3(n29247), .IN4(
        m0s4_data_i[19]), .Q(n22057) );
  AO22X1 U25170 ( .IN1(n29249), .IN2(m0s2_data_i[19]), .IN3(n29250), .IN4(
        m0s1_data_i[19]), .Q(n22056) );
  AO22X1 U25171 ( .IN1(n29245), .IN2(m0s6_data_i[19]), .IN3(n29241), .IN4(
        m0s10_data_i[19]), .Q(n22052) );
  AO22X1 U25172 ( .IN1(n29238), .IN2(m0s13_data_i[19]), .IN3(n29243), .IN4(
        m0s8_data_i[19]), .Q(n22051) );
  NOR2X0 U25173 ( .IN1(n22052), .IN2(n22051), .QN(n22054) );
  NAND2X0 U25174 ( .IN1(n29240), .IN2(m0s11_data_i[19]), .QN(n22053) );
  NAND2X0 U25175 ( .IN1(n22054), .IN2(n22053), .QN(n22055) );
  NOR4X0 U25176 ( .IN1(n22058), .IN2(n22057), .IN3(n22056), .IN4(n22055), .QN(
        n22060) );
  NAND2X0 U25177 ( .IN1(n22198), .IN2(s15_data_i[19]), .QN(n22059) );
  NAND4X0 U25178 ( .IN1(n22062), .IN2(n22061), .IN3(n22060), .IN4(n22059), 
        .QN(m0_data_o[19]) );
  OA22X1 U25179 ( .IN1(n23149), .IN2(n22450), .IN3(n23157), .IN4(n22451), .Q(
        n22074) );
  OA22X1 U25180 ( .IN1(n23127), .IN2(n22453), .IN3(n23135), .IN4(n22448), .Q(
        n22073) );
  AO22X1 U25181 ( .IN1(n29248), .IN2(m0s3_data_i[20]), .IN3(n29238), .IN4(
        m0s13_data_i[20]), .Q(n22070) );
  AO22X1 U25182 ( .IN1(n29242), .IN2(m0s9_data_i[20]), .IN3(n29247), .IN4(
        m0s4_data_i[20]), .Q(n22069) );
  AO22X1 U25183 ( .IN1(n29243), .IN2(m0s8_data_i[20]), .IN3(n29244), .IN4(
        m0s7_data_i[20]), .Q(n22068) );
  AO22X1 U25184 ( .IN1(n29249), .IN2(m0s2_data_i[20]), .IN3(n29250), .IN4(
        m0s1_data_i[20]), .Q(n22064) );
  AO22X1 U25185 ( .IN1(n29239), .IN2(m0s12_data_i[20]), .IN3(n29241), .IN4(
        m0s10_data_i[20]), .Q(n22063) );
  NOR2X0 U25186 ( .IN1(n22064), .IN2(n22063), .QN(n22066) );
  NAND2X0 U25187 ( .IN1(n29245), .IN2(m0s6_data_i[20]), .QN(n22065) );
  NAND2X0 U25188 ( .IN1(n22066), .IN2(n22065), .QN(n22067) );
  NOR4X0 U25189 ( .IN1(n22070), .IN2(n22069), .IN3(n22068), .IN4(n22067), .QN(
        n22072) );
  NAND2X0 U25190 ( .IN1(n22198), .IN2(s15_data_i[20]), .QN(n22071) );
  NAND4X0 U25191 ( .IN1(n22074), .IN2(n22073), .IN3(n22072), .IN4(n22071), 
        .QN(m0_data_o[20]) );
  AO22X1 U25192 ( .IN1(n29239), .IN2(m0s12_data_i[21]), .IN3(n29244), .IN4(
        m0s7_data_i[21]), .Q(n22077) );
  AO22X1 U25193 ( .IN1(n29245), .IN2(m0s6_data_i[21]), .IN3(n29243), .IN4(
        m0s8_data_i[21]), .Q(n22076) );
  AO22X1 U25194 ( .IN1(n29240), .IN2(m0s11_data_i[21]), .IN3(n29241), .IN4(
        m0s10_data_i[21]), .Q(n22075) );
  NOR3X0 U25195 ( .IN1(n22077), .IN2(n22076), .IN3(n22075), .QN(n22085) );
  AO22X1 U25196 ( .IN1(n29248), .IN2(m0s3_data_i[21]), .IN3(n29247), .IN4(
        m0s4_data_i[21]), .Q(n22081) );
  AO22X1 U25197 ( .IN1(n29252), .IN2(m0s0_data_i[21]), .IN3(n29238), .IN4(
        m0s13_data_i[21]), .Q(n22080) );
  AO22X1 U25198 ( .IN1(n29246), .IN2(m0s5_data_i[21]), .IN3(n29242), .IN4(
        m0s9_data_i[21]), .Q(n22079) );
  AO22X1 U25199 ( .IN1(n29237), .IN2(m0s14_data_i[21]), .IN3(n29250), .IN4(
        m0s1_data_i[21]), .Q(n22078) );
  NOR4X0 U25200 ( .IN1(n22081), .IN2(n22080), .IN3(n22079), .IN4(n22078), .QN(
        n22084) );
  NAND2X0 U25201 ( .IN1(n22198), .IN2(s15_data_i[21]), .QN(n22083) );
  NAND2X0 U25202 ( .IN1(n29249), .IN2(m0s2_data_i[21]), .QN(n22082) );
  NAND4X0 U25203 ( .IN1(n22085), .IN2(n22084), .IN3(n22083), .IN4(n22082), 
        .QN(m0_data_o[21]) );
  AO22X1 U25204 ( .IN1(n29252), .IN2(m0s0_data_i[22]), .IN3(n29246), .IN4(
        m0s5_data_i[22]), .Q(n22088) );
  AO22X1 U25205 ( .IN1(n29238), .IN2(m0s13_data_i[22]), .IN3(n29242), .IN4(
        m0s9_data_i[22]), .Q(n22087) );
  AO22X1 U25206 ( .IN1(n29241), .IN2(m0s10_data_i[22]), .IN3(n29249), .IN4(
        m0s2_data_i[22]), .Q(n22086) );
  NOR3X0 U25207 ( .IN1(n22088), .IN2(n22087), .IN3(n22086), .QN(n22096) );
  AO22X1 U25208 ( .IN1(n29239), .IN2(m0s12_data_i[22]), .IN3(n29248), .IN4(
        m0s3_data_i[22]), .Q(n22092) );
  AO22X1 U25209 ( .IN1(n29245), .IN2(m0s6_data_i[22]), .IN3(n29243), .IN4(
        m0s8_data_i[22]), .Q(n22091) );
  AO22X1 U25210 ( .IN1(n29237), .IN2(m0s14_data_i[22]), .IN3(n29250), .IN4(
        m0s1_data_i[22]), .Q(n22090) );
  AO22X1 U25211 ( .IN1(n29240), .IN2(m0s11_data_i[22]), .IN3(n29247), .IN4(
        m0s4_data_i[22]), .Q(n22089) );
  NOR4X0 U25212 ( .IN1(n22092), .IN2(n22091), .IN3(n22090), .IN4(n22089), .QN(
        n22095) );
  NAND2X0 U25213 ( .IN1(n22198), .IN2(s15_data_i[22]), .QN(n22094) );
  NAND2X0 U25214 ( .IN1(n29244), .IN2(m0s7_data_i[22]), .QN(n22093) );
  NAND4X0 U25215 ( .IN1(n22096), .IN2(n22095), .IN3(n22094), .IN4(n22093), 
        .QN(m0_data_o[22]) );
  AO22X1 U25216 ( .IN1(n29239), .IN2(m0s12_data_i[23]), .IN3(n29237), .IN4(
        m0s14_data_i[23]), .Q(n22099) );
  AO22X1 U25217 ( .IN1(n29252), .IN2(m0s0_data_i[23]), .IN3(n29244), .IN4(
        m0s7_data_i[23]), .Q(n22098) );
  AO22X1 U25218 ( .IN1(n29248), .IN2(m0s3_data_i[23]), .IN3(n29243), .IN4(
        m0s8_data_i[23]), .Q(n22097) );
  NOR3X0 U25219 ( .IN1(n22099), .IN2(n22098), .IN3(n22097), .QN(n22107) );
  AO22X1 U25220 ( .IN1(n29245), .IN2(m0s6_data_i[23]), .IN3(n29250), .IN4(
        m0s1_data_i[23]), .Q(n22103) );
  AO22X1 U25221 ( .IN1(n29246), .IN2(m0s5_data_i[23]), .IN3(n29242), .IN4(
        m0s9_data_i[23]), .Q(n22102) );
  AO22X1 U25222 ( .IN1(n29238), .IN2(m0s13_data_i[23]), .IN3(n29247), .IN4(
        m0s4_data_i[23]), .Q(n22101) );
  AO22X1 U25223 ( .IN1(n29240), .IN2(m0s11_data_i[23]), .IN3(n29241), .IN4(
        m0s10_data_i[23]), .Q(n22100) );
  NOR4X0 U25224 ( .IN1(n22103), .IN2(n22102), .IN3(n22101), .IN4(n22100), .QN(
        n22106) );
  NAND2X0 U25225 ( .IN1(n22198), .IN2(s15_data_i[23]), .QN(n22105) );
  NAND2X0 U25226 ( .IN1(n29249), .IN2(m0s2_data_i[23]), .QN(n22104) );
  NAND4X0 U25227 ( .IN1(n22107), .IN2(n22106), .IN3(n22105), .IN4(n22104), 
        .QN(m0_data_o[23]) );
  AO22X1 U25228 ( .IN1(n29240), .IN2(m0s11_data_i[24]), .IN3(n29248), .IN4(
        m0s3_data_i[24]), .Q(n22110) );
  AO22X1 U25229 ( .IN1(n29242), .IN2(m0s9_data_i[24]), .IN3(n29244), .IN4(
        m0s7_data_i[24]), .Q(n22109) );
  AO22X1 U25230 ( .IN1(n29245), .IN2(m0s6_data_i[24]), .IN3(n29250), .IN4(
        m0s1_data_i[24]), .Q(n22108) );
  NOR3X0 U25231 ( .IN1(n22110), .IN2(n22109), .IN3(n22108), .QN(n22118) );
  AO22X1 U25232 ( .IN1(n29237), .IN2(m0s14_data_i[24]), .IN3(n29249), .IN4(
        m0s2_data_i[24]), .Q(n22114) );
  AO22X1 U25233 ( .IN1(n29241), .IN2(m0s10_data_i[24]), .IN3(n29238), .IN4(
        m0s13_data_i[24]), .Q(n22113) );
  AO22X1 U25234 ( .IN1(n29252), .IN2(m0s0_data_i[24]), .IN3(n29246), .IN4(
        m0s5_data_i[24]), .Q(n22112) );
  AO22X1 U25235 ( .IN1(n29239), .IN2(m0s12_data_i[24]), .IN3(n29247), .IN4(
        m0s4_data_i[24]), .Q(n22111) );
  NOR4X0 U25236 ( .IN1(n22114), .IN2(n22113), .IN3(n22112), .IN4(n22111), .QN(
        n22117) );
  NAND2X0 U25237 ( .IN1(n22198), .IN2(s15_data_i[24]), .QN(n22116) );
  NAND2X0 U25238 ( .IN1(n29243), .IN2(m0s8_data_i[24]), .QN(n22115) );
  NAND4X0 U25239 ( .IN1(n22118), .IN2(n22117), .IN3(n22116), .IN4(n22115), 
        .QN(m0_data_o[24]) );
  OA22X1 U25240 ( .IN1(n23127), .IN2(n22524), .IN3(n23167), .IN4(n22521), .Q(
        n22131) );
  OA22X1 U25241 ( .IN1(n23139), .IN2(n22119), .IN3(n23161), .IN4(n22523), .Q(
        n22130) );
  AO22X1 U25242 ( .IN1(n29250), .IN2(m0s1_data_i[25]), .IN3(n29242), .IN4(
        m0s9_data_i[25]), .Q(n22127) );
  AO22X1 U25243 ( .IN1(n29239), .IN2(m0s12_data_i[25]), .IN3(n29252), .IN4(
        m0s0_data_i[25]), .Q(n22126) );
  AO22X1 U25244 ( .IN1(n29240), .IN2(m0s11_data_i[25]), .IN3(n29249), .IN4(
        m0s2_data_i[25]), .Q(n22125) );
  AO22X1 U25245 ( .IN1(n29243), .IN2(m0s8_data_i[25]), .IN3(n29247), .IN4(
        m0s4_data_i[25]), .Q(n22121) );
  AO22X1 U25246 ( .IN1(n29238), .IN2(m0s13_data_i[25]), .IN3(n29246), .IN4(
        m0s5_data_i[25]), .Q(n22120) );
  NOR2X0 U25247 ( .IN1(n22121), .IN2(n22120), .QN(n22123) );
  NAND2X0 U25248 ( .IN1(n29244), .IN2(m0s7_data_i[25]), .QN(n22122) );
  NAND2X0 U25249 ( .IN1(n22123), .IN2(n22122), .QN(n22124) );
  NOR4X0 U25250 ( .IN1(n22127), .IN2(n22126), .IN3(n22125), .IN4(n22124), .QN(
        n22129) );
  NAND2X0 U25251 ( .IN1(n22198), .IN2(s15_data_i[25]), .QN(n22128) );
  NAND4X0 U25252 ( .IN1(n22131), .IN2(n22130), .IN3(n22129), .IN4(n22128), 
        .QN(m0_data_o[25]) );
  AO22X1 U25253 ( .IN1(n29252), .IN2(m0s0_data_i[26]), .IN3(n29250), .IN4(
        m0s1_data_i[26]), .Q(n22134) );
  AO22X1 U25254 ( .IN1(n29239), .IN2(m0s12_data_i[26]), .IN3(n29238), .IN4(
        m0s13_data_i[26]), .Q(n22133) );
  AO22X1 U25255 ( .IN1(n29240), .IN2(m0s11_data_i[26]), .IN3(n29242), .IN4(
        m0s9_data_i[26]), .Q(n22132) );
  NOR3X0 U25256 ( .IN1(n22134), .IN2(n22133), .IN3(n22132), .QN(n22142) );
  AO22X1 U25257 ( .IN1(n29237), .IN2(m0s14_data_i[26]), .IN3(n29249), .IN4(
        m0s2_data_i[26]), .Q(n22138) );
  AO22X1 U25258 ( .IN1(n29247), .IN2(m0s4_data_i[26]), .IN3(n29244), .IN4(
        m0s7_data_i[26]), .Q(n22137) );
  AO22X1 U25259 ( .IN1(n29245), .IN2(m0s6_data_i[26]), .IN3(n29241), .IN4(
        m0s10_data_i[26]), .Q(n22136) );
  AO22X1 U25260 ( .IN1(n29243), .IN2(m0s8_data_i[26]), .IN3(n29246), .IN4(
        m0s5_data_i[26]), .Q(n22135) );
  NOR4X0 U25261 ( .IN1(n22138), .IN2(n22137), .IN3(n22136), .IN4(n22135), .QN(
        n22141) );
  NAND2X0 U25262 ( .IN1(n22198), .IN2(s15_data_i[26]), .QN(n22140) );
  NAND2X0 U25263 ( .IN1(n29248), .IN2(m0s3_data_i[26]), .QN(n22139) );
  NAND4X0 U25264 ( .IN1(n22142), .IN2(n22141), .IN3(n22140), .IN4(n22139), 
        .QN(m0_data_o[26]) );
  AO22X1 U25265 ( .IN1(n29248), .IN2(m0s3_data_i[27]), .IN3(n29243), .IN4(
        m0s8_data_i[27]), .Q(n22145) );
  AO22X1 U25266 ( .IN1(n29245), .IN2(m0s6_data_i[27]), .IN3(n29244), .IN4(
        m0s7_data_i[27]), .Q(n22144) );
  AO22X1 U25267 ( .IN1(n29238), .IN2(m0s13_data_i[27]), .IN3(n29250), .IN4(
        m0s1_data_i[27]), .Q(n22143) );
  NOR3X0 U25268 ( .IN1(n22145), .IN2(n22144), .IN3(n22143), .QN(n22153) );
  AO22X1 U25269 ( .IN1(n29241), .IN2(m0s10_data_i[27]), .IN3(n29247), .IN4(
        m0s4_data_i[27]), .Q(n22149) );
  AO22X1 U25270 ( .IN1(n29237), .IN2(m0s14_data_i[27]), .IN3(n29242), .IN4(
        m0s9_data_i[27]), .Q(n22148) );
  AO22X1 U25271 ( .IN1(n29252), .IN2(m0s0_data_i[27]), .IN3(n29246), .IN4(
        m0s5_data_i[27]), .Q(n22147) );
  AO22X1 U25272 ( .IN1(n29240), .IN2(m0s11_data_i[27]), .IN3(n29249), .IN4(
        m0s2_data_i[27]), .Q(n22146) );
  NOR4X0 U25273 ( .IN1(n22149), .IN2(n22148), .IN3(n22147), .IN4(n22146), .QN(
        n22152) );
  NAND2X0 U25274 ( .IN1(n22198), .IN2(s15_data_i[27]), .QN(n22151) );
  NAND2X0 U25275 ( .IN1(n29239), .IN2(m0s12_data_i[27]), .QN(n22150) );
  NAND4X0 U25276 ( .IN1(n22153), .IN2(n22152), .IN3(n22151), .IN4(n22150), 
        .QN(m0_data_o[27]) );
  OA22X1 U25277 ( .IN1(n23153), .IN2(n22935), .IN3(n23139), .IN4(n22940), .Q(
        n22165) );
  OA22X1 U25278 ( .IN1(n23131), .IN2(n22932), .IN3(n22178), .IN4(n22941), .Q(
        n22164) );
  AO22X1 U25279 ( .IN1(n29248), .IN2(m0s3_data_i[28]), .IN3(n29247), .IN4(
        m0s4_data_i[28]), .Q(n22161) );
  AO22X1 U25280 ( .IN1(n29237), .IN2(m0s14_data_i[28]), .IN3(n29243), .IN4(
        m0s8_data_i[28]), .Q(n22160) );
  AO22X1 U25281 ( .IN1(n29240), .IN2(m0s11_data_i[28]), .IN3(n29252), .IN4(
        m0s0_data_i[28]), .Q(n22159) );
  AO22X1 U25282 ( .IN1(n29249), .IN2(m0s2_data_i[28]), .IN3(n29244), .IN4(
        m0s7_data_i[28]), .Q(n22155) );
  AO22X1 U25283 ( .IN1(n29246), .IN2(m0s5_data_i[28]), .IN3(n29242), .IN4(
        m0s9_data_i[28]), .Q(n22154) );
  NOR2X0 U25284 ( .IN1(n22155), .IN2(n22154), .QN(n22157) );
  NAND2X0 U25285 ( .IN1(n29241), .IN2(m0s10_data_i[28]), .QN(n22156) );
  NAND2X0 U25286 ( .IN1(n22157), .IN2(n22156), .QN(n22158) );
  NOR4X0 U25287 ( .IN1(n22161), .IN2(n22160), .IN3(n22159), .IN4(n22158), .QN(
        n22163) );
  NAND2X0 U25288 ( .IN1(n22198), .IN2(s15_data_i[28]), .QN(n22162) );
  NAND4X0 U25289 ( .IN1(n22165), .IN2(n22164), .IN3(n22163), .IN4(n22162), 
        .QN(m0_data_o[28]) );
  AO22X1 U25290 ( .IN1(n29237), .IN2(m0s14_data_i[29]), .IN3(n29252), .IN4(
        m0s0_data_i[29]), .Q(n22168) );
  AO22X1 U25291 ( .IN1(n29248), .IN2(m0s3_data_i[29]), .IN3(n29238), .IN4(
        m0s13_data_i[29]), .Q(n22167) );
  AO22X1 U25292 ( .IN1(n29241), .IN2(m0s10_data_i[29]), .IN3(n29249), .IN4(
        m0s2_data_i[29]), .Q(n22166) );
  NOR3X0 U25293 ( .IN1(n22168), .IN2(n22167), .IN3(n22166), .QN(n22176) );
  AO22X1 U25294 ( .IN1(n29245), .IN2(m0s6_data_i[29]), .IN3(n29247), .IN4(
        m0s4_data_i[29]), .Q(n22172) );
  AO22X1 U25295 ( .IN1(n29239), .IN2(m0s12_data_i[29]), .IN3(n29240), .IN4(
        m0s11_data_i[29]), .Q(n22171) );
  AO22X1 U25296 ( .IN1(n29242), .IN2(m0s9_data_i[29]), .IN3(n29244), .IN4(
        m0s7_data_i[29]), .Q(n22170) );
  AO22X1 U25297 ( .IN1(n29243), .IN2(m0s8_data_i[29]), .IN3(n29246), .IN4(
        m0s5_data_i[29]), .Q(n22169) );
  NOR4X0 U25298 ( .IN1(n22172), .IN2(n22171), .IN3(n22170), .IN4(n22169), .QN(
        n22175) );
  NAND2X0 U25299 ( .IN1(n22198), .IN2(s15_data_i[29]), .QN(n22174) );
  NAND2X0 U25300 ( .IN1(n29250), .IN2(m0s1_data_i[29]), .QN(n22173) );
  NAND4X0 U25301 ( .IN1(n22176), .IN2(n22175), .IN3(n22174), .IN4(n22173), 
        .QN(m0_data_o[29]) );
  OA22X1 U25302 ( .IN1(n23127), .IN2(n22597), .IN3(n23157), .IN4(n22177), .Q(
        n22190) );
  OA22X1 U25303 ( .IN1(n23131), .IN2(n22602), .IN3(n22178), .IN4(n22601), .Q(
        n22189) );
  AO22X1 U25304 ( .IN1(n29239), .IN2(m0s12_data_i[30]), .IN3(n29242), .IN4(
        m0s9_data_i[30]), .Q(n22186) );
  AO22X1 U25305 ( .IN1(n29248), .IN2(m0s3_data_i[30]), .IN3(n29244), .IN4(
        m0s7_data_i[30]), .Q(n22185) );
  AO22X1 U25306 ( .IN1(n29245), .IN2(m0s6_data_i[30]), .IN3(n29241), .IN4(
        m0s10_data_i[30]), .Q(n22184) );
  AO22X1 U25307 ( .IN1(n29243), .IN2(m0s8_data_i[30]), .IN3(n29246), .IN4(
        m0s5_data_i[30]), .Q(n22180) );
  AO22X1 U25308 ( .IN1(n29249), .IN2(m0s2_data_i[30]), .IN3(n29247), .IN4(
        m0s4_data_i[30]), .Q(n22179) );
  NOR2X0 U25309 ( .IN1(n22180), .IN2(n22179), .QN(n22182) );
  NAND2X0 U25310 ( .IN1(n29240), .IN2(m0s11_data_i[30]), .QN(n22181) );
  NAND2X0 U25311 ( .IN1(n22182), .IN2(n22181), .QN(n22183) );
  NOR4X0 U25312 ( .IN1(n22186), .IN2(n22185), .IN3(n22184), .IN4(n22183), .QN(
        n22188) );
  NAND2X0 U25313 ( .IN1(n22198), .IN2(s15_data_i[30]), .QN(n22187) );
  NAND4X0 U25314 ( .IN1(n22190), .IN2(n22189), .IN3(n22188), .IN4(n22187), 
        .QN(m0_data_o[30]) );
  AO22X1 U25315 ( .IN1(n29239), .IN2(m0s12_data_i[31]), .IN3(n29244), .IN4(
        m0s7_data_i[31]), .Q(n22193) );
  AO22X1 U25316 ( .IN1(n29237), .IN2(m0s14_data_i[31]), .IN3(n29243), .IN4(
        m0s8_data_i[31]), .Q(n22192) );
  AO22X1 U25317 ( .IN1(n29238), .IN2(m0s13_data_i[31]), .IN3(n29242), .IN4(
        m0s9_data_i[31]), .Q(n22191) );
  NOR3X0 U25318 ( .IN1(n22193), .IN2(n22192), .IN3(n22191), .QN(n22202) );
  AO22X1 U25319 ( .IN1(n29252), .IN2(m0s0_data_i[31]), .IN3(n29246), .IN4(
        m0s5_data_i[31]), .Q(n22197) );
  AO22X1 U25320 ( .IN1(n29245), .IN2(m0s6_data_i[31]), .IN3(n29247), .IN4(
        m0s4_data_i[31]), .Q(n22196) );
  AO22X1 U25321 ( .IN1(n29248), .IN2(m0s3_data_i[31]), .IN3(n29250), .IN4(
        m0s1_data_i[31]), .Q(n22195) );
  AO22X1 U25322 ( .IN1(n29241), .IN2(m0s10_data_i[31]), .IN3(n29249), .IN4(
        m0s2_data_i[31]), .Q(n22194) );
  NOR4X0 U25323 ( .IN1(n22197), .IN2(n22196), .IN3(n22195), .IN4(n22194), .QN(
        n22201) );
  NAND2X0 U25324 ( .IN1(n22198), .IN2(s15_data_i[31]), .QN(n22200) );
  NAND2X0 U25325 ( .IN1(n29240), .IN2(m0s11_data_i[31]), .QN(n22199) );
  NAND4X0 U25326 ( .IN1(n22202), .IN2(n22201), .IN3(n22200), .IN4(n22199), 
        .QN(m0_data_o[31]) );
  INVX0 U25327 ( .INP(n29271), .ZN(n22569) );
  OA22X1 U25328 ( .IN1(n22204), .IN2(n22569), .IN3(n22203), .IN4(n22567), .Q(
        n22222) );
  OA22X1 U25329 ( .IN1(n22206), .IN2(n23235), .IN3(n22205), .IN4(n22620), .Q(
        n22221) );
  INVX0 U25330 ( .INP(n22584), .ZN(n29263) );
  AO22X1 U25331 ( .IN1(m0s5_data_i[0]), .IN2(n29265), .IN3(m0s7_data_i[0]), 
        .IN4(n29263), .Q(n22216) );
  INVX0 U25332 ( .INP(n23232), .ZN(n29264) );
  AO22X1 U25333 ( .IN1(m0s6_data_i[0]), .IN2(n29264), .IN3(m0s13_data_i[0]), 
        .IN4(n29257), .Q(n22215) );
  INVX0 U25334 ( .INP(n23238), .ZN(n29269) );
  INVX0 U25335 ( .INP(n22582), .ZN(n29261) );
  AO22X1 U25336 ( .IN1(m0s1_data_i[0]), .IN2(n29269), .IN3(m0s9_data_i[0]), 
        .IN4(n29261), .Q(n22214) );
  OA22X1 U25337 ( .IN1(n22208), .IN2(n23223), .IN3(n22207), .IN4(n22599), .Q(
        n22212) );
  NAND2X0 U25338 ( .IN1(m0s8_data_i[0]), .IN2(n29262), .QN(n22211) );
  INVX0 U25339 ( .INP(n23241), .ZN(n29256) );
  NAND2X0 U25340 ( .IN1(m0s14_data_i[0]), .IN2(n29256), .QN(n22210) );
  INVX0 U25341 ( .INP(n23226), .ZN(n29258) );
  NAND2X0 U25342 ( .IN1(m0s12_data_i[0]), .IN2(n29258), .QN(n22209) );
  NAND4X0 U25343 ( .IN1(n22212), .IN2(n22211), .IN3(n22210), .IN4(n22209), 
        .QN(n22213) );
  NOR4X0 U25344 ( .IN1(n22216), .IN2(n22215), .IN3(n22214), .IN4(n22213), .QN(
        n22220) );
  INVX0 U25345 ( .INP(n22217), .ZN(n29255) );
  NAND2X0 U25346 ( .IN1(n29255), .IN2(n22218), .QN(n22219) );
  NAND4X0 U25347 ( .IN1(n22222), .IN2(n22221), .IN3(n22220), .IN4(n22219), 
        .QN(m1_data_o[0]) );
  OA22X1 U25348 ( .IN1(n22224), .IN2(n23241), .IN3(n22223), .IN4(n22569), .Q(
        n22239) );
  OA22X1 U25349 ( .IN1(n22226), .IN2(n22584), .IN3(n22225), .IN4(n22620), .Q(
        n22238) );
  AO22X1 U25350 ( .IN1(m0s3_data_i[1]), .IN2(n29267), .IN3(m0s9_data_i[1]), 
        .IN4(n29261), .Q(n22234) );
  INVX0 U25351 ( .INP(n22567), .ZN(n29266) );
  AO22X1 U25352 ( .IN1(m0s1_data_i[1]), .IN2(n29269), .IN3(m0s4_data_i[1]), 
        .IN4(n29266), .Q(n22233) );
  AO22X1 U25353 ( .IN1(m0s5_data_i[1]), .IN2(n29265), .IN3(m0s6_data_i[1]), 
        .IN4(n29264), .Q(n22232) );
  INVX0 U25354 ( .INP(n22599), .ZN(n29260) );
  AO22X1 U25355 ( .IN1(m0s12_data_i[1]), .IN2(n29258), .IN3(m0s10_data_i[1]), 
        .IN4(n29260), .Q(n22228) );
  AO22X1 U25356 ( .IN1(m0s8_data_i[1]), .IN2(n29262), .IN3(m0s11_data_i[1]), 
        .IN4(n29259), .Q(n22227) );
  NOR2X0 U25357 ( .IN1(n22228), .IN2(n22227), .QN(n22230) );
  NAND2X0 U25358 ( .IN1(m0s13_data_i[1]), .IN2(n29257), .QN(n22229) );
  NAND2X0 U25359 ( .IN1(n22230), .IN2(n22229), .QN(n22231) );
  NOR4X0 U25360 ( .IN1(n22234), .IN2(n22233), .IN3(n22232), .IN4(n22231), .QN(
        n22237) );
  NAND2X0 U25361 ( .IN1(n29255), .IN2(n22235), .QN(n22236) );
  NAND4X0 U25362 ( .IN1(n22239), .IN2(n22238), .IN3(n22237), .IN4(n22236), 
        .QN(m1_data_o[1]) );
  AO22X1 U25363 ( .IN1(m0s7_data_i[2]), .IN2(n29263), .IN3(m0s0_data_i[2]), 
        .IN4(n29271), .Q(n22242) );
  AO22X1 U25364 ( .IN1(m0s13_data_i[2]), .IN2(n29257), .IN3(m0s11_data_i[2]), 
        .IN4(n29259), .Q(n22241) );
  AO22X1 U25365 ( .IN1(m0s3_data_i[2]), .IN2(n29267), .IN3(m0s1_data_i[2]), 
        .IN4(n29269), .Q(n22240) );
  NOR3X0 U25366 ( .IN1(n22242), .IN2(n22241), .IN3(n22240), .QN(n22251) );
  INVX0 U25367 ( .INP(n22620), .ZN(n29268) );
  AO22X1 U25368 ( .IN1(m0s8_data_i[2]), .IN2(n29262), .IN3(m0s2_data_i[2]), 
        .IN4(n29268), .Q(n22246) );
  AO22X1 U25369 ( .IN1(m0s4_data_i[2]), .IN2(n29266), .IN3(m0s6_data_i[2]), 
        .IN4(n29264), .Q(n22245) );
  AO22X1 U25370 ( .IN1(m0s9_data_i[2]), .IN2(n29261), .IN3(m0s14_data_i[2]), 
        .IN4(n29256), .Q(n22244) );
  AO22X1 U25371 ( .IN1(m0s12_data_i[2]), .IN2(n29258), .IN3(m0s10_data_i[2]), 
        .IN4(n29260), .Q(n22243) );
  NOR4X0 U25372 ( .IN1(n22246), .IN2(n22245), .IN3(n22244), .IN4(n22243), .QN(
        n22250) );
  NAND2X0 U25373 ( .IN1(n29255), .IN2(n22247), .QN(n22249) );
  NAND2X0 U25374 ( .IN1(m0s5_data_i[2]), .IN2(n29265), .QN(n22248) );
  NAND4X0 U25375 ( .IN1(n22251), .IN2(n22250), .IN3(n22249), .IN4(n22248), 
        .QN(m1_data_o[2]) );
  AO22X1 U25376 ( .IN1(m0s1_data_i[3]), .IN2(n29269), .IN3(m0s0_data_i[3]), 
        .IN4(n29271), .Q(n22254) );
  AO22X1 U25377 ( .IN1(m0s11_data_i[3]), .IN2(n29259), .IN3(m0s6_data_i[3]), 
        .IN4(n29264), .Q(n22253) );
  AO22X1 U25378 ( .IN1(m0s3_data_i[3]), .IN2(n29267), .IN3(m0s4_data_i[3]), 
        .IN4(n29266), .Q(n22252) );
  NOR3X0 U25379 ( .IN1(n22254), .IN2(n22253), .IN3(n22252), .QN(n22262) );
  AO22X1 U25380 ( .IN1(m0s12_data_i[3]), .IN2(n29258), .IN3(m0s2_data_i[3]), 
        .IN4(n29268), .Q(n22258) );
  AO22X1 U25381 ( .IN1(m0s5_data_i[3]), .IN2(n29265), .IN3(m0s14_data_i[3]), 
        .IN4(n29256), .Q(n22257) );
  AO22X1 U25382 ( .IN1(m0s7_data_i[3]), .IN2(n29263), .IN3(m0s10_data_i[3]), 
        .IN4(n29260), .Q(n22256) );
  AO22X1 U25383 ( .IN1(m0s9_data_i[3]), .IN2(n29261), .IN3(m0s8_data_i[3]), 
        .IN4(n29262), .Q(n22255) );
  NOR4X0 U25384 ( .IN1(n22258), .IN2(n22257), .IN3(n22256), .IN4(n22255), .QN(
        n22261) );
  NAND2X0 U25385 ( .IN1(n29255), .IN2(n22646), .QN(n22260) );
  NAND2X0 U25386 ( .IN1(m0s13_data_i[3]), .IN2(n29257), .QN(n22259) );
  NAND4X0 U25387 ( .IN1(n22262), .IN2(n22261), .IN3(n22260), .IN4(n22259), 
        .QN(m1_data_o[3]) );
  AO22X1 U25388 ( .IN1(m0s12_data_i[4]), .IN2(n29258), .IN3(m0s2_data_i[4]), 
        .IN4(n29268), .Q(n22265) );
  AO22X1 U25389 ( .IN1(m0s4_data_i[4]), .IN2(n29266), .IN3(m0s9_data_i[4]), 
        .IN4(n29261), .Q(n22264) );
  AO22X1 U25390 ( .IN1(m0s5_data_i[4]), .IN2(n29265), .IN3(m0s10_data_i[4]), 
        .IN4(n29260), .Q(n22263) );
  NOR3X0 U25391 ( .IN1(n22265), .IN2(n22264), .IN3(n22263), .QN(n22273) );
  AO22X1 U25392 ( .IN1(m0s6_data_i[4]), .IN2(n29264), .IN3(m0s8_data_i[4]), 
        .IN4(n29262), .Q(n22269) );
  AO22X1 U25393 ( .IN1(m0s11_data_i[4]), .IN2(n29259), .IN3(m0s0_data_i[4]), 
        .IN4(n29271), .Q(n22268) );
  AO22X1 U25394 ( .IN1(m0s13_data_i[4]), .IN2(n29257), .IN3(m0s14_data_i[4]), 
        .IN4(n29256), .Q(n22267) );
  AO22X1 U25395 ( .IN1(m0s3_data_i[4]), .IN2(n29267), .IN3(m0s7_data_i[4]), 
        .IN4(n29263), .Q(n22266) );
  NOR4X0 U25396 ( .IN1(n22269), .IN2(n22268), .IN3(n22267), .IN4(n22266), .QN(
        n22272) );
  NAND2X0 U25397 ( .IN1(n29255), .IN2(n22663), .QN(n22271) );
  NAND2X0 U25398 ( .IN1(m0s1_data_i[4]), .IN2(n29269), .QN(n22270) );
  NAND4X0 U25399 ( .IN1(n22273), .IN2(n22272), .IN3(n22271), .IN4(n22270), 
        .QN(m1_data_o[4]) );
  AO22X1 U25400 ( .IN1(m0s14_data_i[5]), .IN2(n29256), .IN3(m0s1_data_i[5]), 
        .IN4(n29269), .Q(n22276) );
  AO22X1 U25401 ( .IN1(m0s10_data_i[5]), .IN2(n29260), .IN3(m0s3_data_i[5]), 
        .IN4(n29267), .Q(n22275) );
  AO22X1 U25402 ( .IN1(m0s6_data_i[5]), .IN2(n29264), .IN3(m0s0_data_i[5]), 
        .IN4(n29271), .Q(n22274) );
  NOR3X0 U25403 ( .IN1(n22276), .IN2(n22275), .IN3(n22274), .QN(n22284) );
  AO22X1 U25404 ( .IN1(m0s7_data_i[5]), .IN2(n29263), .IN3(m0s11_data_i[5]), 
        .IN4(n29259), .Q(n22280) );
  AO22X1 U25405 ( .IN1(m0s4_data_i[5]), .IN2(n29266), .IN3(m0s5_data_i[5]), 
        .IN4(n29265), .Q(n22279) );
  AO22X1 U25406 ( .IN1(m0s12_data_i[5]), .IN2(n29258), .IN3(m0s9_data_i[5]), 
        .IN4(n29261), .Q(n22278) );
  AO22X1 U25407 ( .IN1(m0s2_data_i[5]), .IN2(n29268), .IN3(m0s8_data_i[5]), 
        .IN4(n29262), .Q(n22277) );
  NOR4X0 U25408 ( .IN1(n22280), .IN2(n22279), .IN3(n22278), .IN4(n22277), .QN(
        n22283) );
  NAND2X0 U25409 ( .IN1(n29255), .IN2(n22680), .QN(n22282) );
  NAND2X0 U25410 ( .IN1(m0s13_data_i[5]), .IN2(n29257), .QN(n22281) );
  NAND4X0 U25411 ( .IN1(n22284), .IN2(n22283), .IN3(n22282), .IN4(n22281), 
        .QN(m1_data_o[5]) );
  AO22X1 U25412 ( .IN1(m0s12_data_i[6]), .IN2(n29258), .IN3(m0s7_data_i[6]), 
        .IN4(n29263), .Q(n22287) );
  AO22X1 U25413 ( .IN1(m0s14_data_i[6]), .IN2(n29256), .IN3(m0s1_data_i[6]), 
        .IN4(n29269), .Q(n22286) );
  AO22X1 U25414 ( .IN1(m0s6_data_i[6]), .IN2(n29264), .IN3(m0s11_data_i[6]), 
        .IN4(n29259), .Q(n22285) );
  NOR3X0 U25415 ( .IN1(n22287), .IN2(n22286), .IN3(n22285), .QN(n22295) );
  AO22X1 U25416 ( .IN1(m0s10_data_i[6]), .IN2(n29260), .IN3(m0s0_data_i[6]), 
        .IN4(n29271), .Q(n22291) );
  AO22X1 U25417 ( .IN1(m0s5_data_i[6]), .IN2(n29265), .IN3(m0s9_data_i[6]), 
        .IN4(n29261), .Q(n22290) );
  AO22X1 U25418 ( .IN1(m0s8_data_i[6]), .IN2(n29262), .IN3(m0s13_data_i[6]), 
        .IN4(n29257), .Q(n22289) );
  AO22X1 U25419 ( .IN1(m0s2_data_i[6]), .IN2(n29268), .IN3(m0s4_data_i[6]), 
        .IN4(n29266), .Q(n22288) );
  NOR4X0 U25420 ( .IN1(n22291), .IN2(n22290), .IN3(n22289), .IN4(n22288), .QN(
        n22294) );
  NAND2X0 U25421 ( .IN1(n29255), .IN2(n22697), .QN(n22293) );
  NAND2X0 U25422 ( .IN1(m0s3_data_i[6]), .IN2(n29267), .QN(n22292) );
  NAND4X0 U25423 ( .IN1(n22295), .IN2(n22294), .IN3(n22293), .IN4(n22292), 
        .QN(m1_data_o[6]) );
  AO22X1 U25424 ( .IN1(m0s12_data_i[7]), .IN2(n29258), .IN3(m0s0_data_i[7]), 
        .IN4(n29271), .Q(n22298) );
  AO22X1 U25425 ( .IN1(m0s11_data_i[7]), .IN2(n29259), .IN3(m0s2_data_i[7]), 
        .IN4(n29268), .Q(n22297) );
  AO22X1 U25426 ( .IN1(m0s6_data_i[7]), .IN2(n29264), .IN3(m0s14_data_i[7]), 
        .IN4(n29256), .Q(n22296) );
  NOR3X0 U25427 ( .IN1(n22298), .IN2(n22297), .IN3(n22296), .QN(n22306) );
  AO22X1 U25428 ( .IN1(m0s3_data_i[7]), .IN2(n29267), .IN3(m0s13_data_i[7]), 
        .IN4(n29257), .Q(n22302) );
  AO22X1 U25429 ( .IN1(m0s1_data_i[7]), .IN2(n29269), .IN3(m0s10_data_i[7]), 
        .IN4(n29260), .Q(n22301) );
  AO22X1 U25430 ( .IN1(m0s4_data_i[7]), .IN2(n29266), .IN3(m0s7_data_i[7]), 
        .IN4(n29263), .Q(n22300) );
  AO22X1 U25431 ( .IN1(m0s5_data_i[7]), .IN2(n29265), .IN3(m0s9_data_i[7]), 
        .IN4(n29261), .Q(n22299) );
  NOR4X0 U25432 ( .IN1(n22302), .IN2(n22301), .IN3(n22300), .IN4(n22299), .QN(
        n22305) );
  NAND2X0 U25433 ( .IN1(n29255), .IN2(n22714), .QN(n22304) );
  NAND2X0 U25434 ( .IN1(m0s8_data_i[7]), .IN2(n29262), .QN(n22303) );
  NAND4X0 U25435 ( .IN1(n22306), .IN2(n22305), .IN3(n22304), .IN4(n22303), 
        .QN(m1_data_o[7]) );
  AO22X1 U25436 ( .IN1(m0s12_data_i[8]), .IN2(n29258), .IN3(m0s0_data_i[8]), 
        .IN4(n29271), .Q(n22309) );
  AO22X1 U25437 ( .IN1(m0s11_data_i[8]), .IN2(n29259), .IN3(m0s2_data_i[8]), 
        .IN4(n29268), .Q(n22308) );
  AO22X1 U25438 ( .IN1(m0s14_data_i[8]), .IN2(n29256), .IN3(m0s9_data_i[8]), 
        .IN4(n29261), .Q(n22307) );
  NOR3X0 U25439 ( .IN1(n22309), .IN2(n22308), .IN3(n22307), .QN(n22317) );
  AO22X1 U25440 ( .IN1(m0s1_data_i[8]), .IN2(n29269), .IN3(m0s3_data_i[8]), 
        .IN4(n29267), .Q(n22313) );
  AO22X1 U25441 ( .IN1(m0s5_data_i[8]), .IN2(n29265), .IN3(m0s6_data_i[8]), 
        .IN4(n29264), .Q(n22312) );
  AO22X1 U25442 ( .IN1(m0s13_data_i[8]), .IN2(n29257), .IN3(m0s8_data_i[8]), 
        .IN4(n29262), .Q(n22311) );
  AO22X1 U25443 ( .IN1(m0s7_data_i[8]), .IN2(n29263), .IN3(m0s10_data_i[8]), 
        .IN4(n29260), .Q(n22310) );
  NOR4X0 U25444 ( .IN1(n22313), .IN2(n22312), .IN3(n22311), .IN4(n22310), .QN(
        n22316) );
  NAND2X0 U25445 ( .IN1(n29255), .IN2(n22731), .QN(n22315) );
  NAND2X0 U25446 ( .IN1(m0s4_data_i[8]), .IN2(n29266), .QN(n22314) );
  NAND4X0 U25447 ( .IN1(n22317), .IN2(n22316), .IN3(n22315), .IN4(n22314), 
        .QN(m1_data_o[8]) );
  AO22X1 U25448 ( .IN1(m0s3_data_i[9]), .IN2(n29267), .IN3(m0s11_data_i[9]), 
        .IN4(n29259), .Q(n22320) );
  AO22X1 U25449 ( .IN1(m0s9_data_i[9]), .IN2(n29261), .IN3(m0s4_data_i[9]), 
        .IN4(n29266), .Q(n22319) );
  AO22X1 U25450 ( .IN1(m0s8_data_i[9]), .IN2(n29262), .IN3(m0s14_data_i[9]), 
        .IN4(n29256), .Q(n22318) );
  NOR3X0 U25451 ( .IN1(n22320), .IN2(n22319), .IN3(n22318), .QN(n22328) );
  AO22X1 U25452 ( .IN1(m0s12_data_i[9]), .IN2(n29258), .IN3(m0s5_data_i[9]), 
        .IN4(n29265), .Q(n22324) );
  AO22X1 U25453 ( .IN1(m0s10_data_i[9]), .IN2(n29260), .IN3(m0s7_data_i[9]), 
        .IN4(n29263), .Q(n22323) );
  AO22X1 U25454 ( .IN1(m0s13_data_i[9]), .IN2(n29257), .IN3(m0s0_data_i[9]), 
        .IN4(n29271), .Q(n22322) );
  AO22X1 U25455 ( .IN1(m0s6_data_i[9]), .IN2(n29264), .IN3(m0s1_data_i[9]), 
        .IN4(n29269), .Q(n22321) );
  NOR4X0 U25456 ( .IN1(n22324), .IN2(n22323), .IN3(n22322), .IN4(n22321), .QN(
        n22327) );
  NAND2X0 U25457 ( .IN1(n29255), .IN2(n22993), .QN(n22326) );
  NAND2X0 U25458 ( .IN1(m0s2_data_i[9]), .IN2(n29268), .QN(n22325) );
  NAND4X0 U25459 ( .IN1(n22328), .IN2(n22327), .IN3(n22326), .IN4(n22325), 
        .QN(m1_data_o[9]) );
  OA22X1 U25460 ( .IN1(n22329), .IN2(n23241), .IN3(n22749), .IN4(n22620), .Q(
        n22341) );
  OA22X1 U25461 ( .IN1(n22753), .IN2(n22567), .IN3(n22751), .IN4(n22599), .Q(
        n22340) );
  AO22X1 U25462 ( .IN1(m0s8_data_i[10]), .IN2(n29262), .IN3(m0s0_data_i[10]), 
        .IN4(n29271), .Q(n22337) );
  AO22X1 U25463 ( .IN1(m0s7_data_i[10]), .IN2(n29263), .IN3(m0s3_data_i[10]), 
        .IN4(n29267), .Q(n22336) );
  AO22X1 U25464 ( .IN1(m0s6_data_i[10]), .IN2(n29264), .IN3(m0s5_data_i[10]), 
        .IN4(n29265), .Q(n22335) );
  AO22X1 U25465 ( .IN1(m0s13_data_i[10]), .IN2(n29257), .IN3(m0s11_data_i[10]), 
        .IN4(n29259), .Q(n22331) );
  AO22X1 U25466 ( .IN1(m0s12_data_i[10]), .IN2(n29258), .IN3(m0s1_data_i[10]), 
        .IN4(n29269), .Q(n22330) );
  NOR2X0 U25467 ( .IN1(n22331), .IN2(n22330), .QN(n22333) );
  NAND2X0 U25468 ( .IN1(m0s9_data_i[10]), .IN2(n29261), .QN(n22332) );
  NAND2X0 U25469 ( .IN1(n22333), .IN2(n22332), .QN(n22334) );
  NOR4X0 U25470 ( .IN1(n22337), .IN2(n22336), .IN3(n22335), .IN4(n22334), .QN(
        n22339) );
  NAND2X0 U25471 ( .IN1(n29255), .IN2(n22763), .QN(n22338) );
  NAND4X0 U25472 ( .IN1(n22341), .IN2(n22340), .IN3(n22339), .IN4(n22338), 
        .QN(m1_data_o[10]) );
  AO22X1 U25473 ( .IN1(m0s12_data_i[11]), .IN2(n29258), .IN3(m0s7_data_i[11]), 
        .IN4(n29263), .Q(n22344) );
  AO22X1 U25474 ( .IN1(m0s13_data_i[11]), .IN2(n29257), .IN3(m0s6_data_i[11]), 
        .IN4(n29264), .Q(n22343) );
  AO22X1 U25475 ( .IN1(m0s11_data_i[11]), .IN2(n29259), .IN3(m0s10_data_i[11]), 
        .IN4(n29260), .Q(n22342) );
  NOR3X0 U25476 ( .IN1(n22344), .IN2(n22343), .IN3(n22342), .QN(n22352) );
  AO22X1 U25477 ( .IN1(m0s14_data_i[11]), .IN2(n29256), .IN3(m0s0_data_i[11]), 
        .IN4(n29271), .Q(n22348) );
  AO22X1 U25478 ( .IN1(m0s3_data_i[11]), .IN2(n29267), .IN3(m0s5_data_i[11]), 
        .IN4(n29265), .Q(n22347) );
  AO22X1 U25479 ( .IN1(m0s2_data_i[11]), .IN2(n29268), .IN3(m0s4_data_i[11]), 
        .IN4(n29266), .Q(n22346) );
  AO22X1 U25480 ( .IN1(m0s1_data_i[11]), .IN2(n29269), .IN3(m0s9_data_i[11]), 
        .IN4(n29261), .Q(n22345) );
  NOR4X0 U25481 ( .IN1(n22348), .IN2(n22347), .IN3(n22346), .IN4(n22345), .QN(
        n22351) );
  NAND2X0 U25482 ( .IN1(n29255), .IN2(n23013), .QN(n22350) );
  NAND2X0 U25483 ( .IN1(m0s8_data_i[11]), .IN2(n29262), .QN(n22349) );
  NAND4X0 U25484 ( .IN1(n22352), .IN2(n22351), .IN3(n22350), .IN4(n22349), 
        .QN(m1_data_o[11]) );
  AO22X1 U25485 ( .IN1(m0s9_data_i[12]), .IN2(n29261), .IN3(m0s0_data_i[12]), 
        .IN4(n29271), .Q(n22355) );
  AO22X1 U25486 ( .IN1(m0s4_data_i[12]), .IN2(n29266), .IN3(m0s13_data_i[12]), 
        .IN4(n29257), .Q(n22354) );
  AO22X1 U25487 ( .IN1(m0s11_data_i[12]), .IN2(n29259), .IN3(m0s3_data_i[12]), 
        .IN4(n29267), .Q(n22353) );
  NOR3X0 U25488 ( .IN1(n22355), .IN2(n22354), .IN3(n22353), .QN(n22363) );
  AO22X1 U25489 ( .IN1(m0s8_data_i[12]), .IN2(n29262), .IN3(m0s5_data_i[12]), 
        .IN4(n29265), .Q(n22359) );
  AO22X1 U25490 ( .IN1(m0s7_data_i[12]), .IN2(n29263), .IN3(m0s6_data_i[12]), 
        .IN4(n29264), .Q(n22358) );
  AO22X1 U25491 ( .IN1(m0s10_data_i[12]), .IN2(n29260), .IN3(m0s12_data_i[12]), 
        .IN4(n29258), .Q(n22357) );
  AO22X1 U25492 ( .IN1(m0s2_data_i[12]), .IN2(n29268), .IN3(m0s1_data_i[12]), 
        .IN4(n29269), .Q(n22356) );
  NOR4X0 U25493 ( .IN1(n22359), .IN2(n22358), .IN3(n22357), .IN4(n22356), .QN(
        n22362) );
  NAND2X0 U25494 ( .IN1(n29255), .IN2(n23034), .QN(n22361) );
  NAND2X0 U25495 ( .IN1(m0s14_data_i[12]), .IN2(n29256), .QN(n22360) );
  NAND4X0 U25496 ( .IN1(n22363), .IN2(n22362), .IN3(n22361), .IN4(n22360), 
        .QN(m1_data_o[12]) );
  AO22X1 U25497 ( .IN1(m0s4_data_i[13]), .IN2(n29266), .IN3(m0s5_data_i[13]), 
        .IN4(n29265), .Q(n22366) );
  AO22X1 U25498 ( .IN1(m0s1_data_i[13]), .IN2(n29269), .IN3(m0s14_data_i[13]), 
        .IN4(n29256), .Q(n22365) );
  AO22X1 U25499 ( .IN1(m0s10_data_i[13]), .IN2(n29260), .IN3(m0s9_data_i[13]), 
        .IN4(n29261), .Q(n22364) );
  NOR3X0 U25500 ( .IN1(n22366), .IN2(n22365), .IN3(n22364), .QN(n22374) );
  AO22X1 U25501 ( .IN1(m0s7_data_i[13]), .IN2(n29263), .IN3(m0s11_data_i[13]), 
        .IN4(n29259), .Q(n22370) );
  AO22X1 U25502 ( .IN1(m0s6_data_i[13]), .IN2(n29264), .IN3(m0s3_data_i[13]), 
        .IN4(n29267), .Q(n22369) );
  AO22X1 U25503 ( .IN1(m0s8_data_i[13]), .IN2(n29262), .IN3(m0s2_data_i[13]), 
        .IN4(n29268), .Q(n22368) );
  AO22X1 U25504 ( .IN1(m0s13_data_i[13]), .IN2(n29257), .IN3(m0s12_data_i[13]), 
        .IN4(n29258), .Q(n22367) );
  NOR4X0 U25505 ( .IN1(n22370), .IN2(n22369), .IN3(n22368), .IN4(n22367), .QN(
        n22373) );
  NAND2X0 U25506 ( .IN1(n29255), .IN2(n23053), .QN(n22372) );
  NAND2X0 U25507 ( .IN1(m0s0_data_i[13]), .IN2(n29271), .QN(n22371) );
  NAND4X0 U25508 ( .IN1(n22374), .IN2(n22373), .IN3(n22372), .IN4(n22371), 
        .QN(m1_data_o[13]) );
  AO22X1 U25509 ( .IN1(m0s5_data_i[14]), .IN2(n29265), .IN3(m0s12_data_i[14]), 
        .IN4(n29258), .Q(n22377) );
  AO22X1 U25510 ( .IN1(m0s2_data_i[14]), .IN2(n29268), .IN3(m0s7_data_i[14]), 
        .IN4(n29263), .Q(n22376) );
  AO22X1 U25511 ( .IN1(m0s9_data_i[14]), .IN2(n29261), .IN3(m0s4_data_i[14]), 
        .IN4(n29266), .Q(n22375) );
  NOR3X0 U25512 ( .IN1(n22377), .IN2(n22376), .IN3(n22375), .QN(n22385) );
  AO22X1 U25513 ( .IN1(m0s8_data_i[14]), .IN2(n29262), .IN3(m0s14_data_i[14]), 
        .IN4(n29256), .Q(n22381) );
  AO22X1 U25514 ( .IN1(m0s0_data_i[14]), .IN2(n29271), .IN3(m0s3_data_i[14]), 
        .IN4(n29267), .Q(n22380) );
  AO22X1 U25515 ( .IN1(m0s10_data_i[14]), .IN2(n29260), .IN3(m0s13_data_i[14]), 
        .IN4(n29257), .Q(n22379) );
  AO22X1 U25516 ( .IN1(m0s6_data_i[14]), .IN2(n29264), .IN3(m0s11_data_i[14]), 
        .IN4(n29259), .Q(n22378) );
  NOR4X0 U25517 ( .IN1(n22381), .IN2(n22380), .IN3(n22379), .IN4(n22378), .QN(
        n22384) );
  NAND2X0 U25518 ( .IN1(n29255), .IN2(n23078), .QN(n22383) );
  NAND2X0 U25519 ( .IN1(m0s1_data_i[14]), .IN2(n29269), .QN(n22382) );
  NAND4X0 U25520 ( .IN1(n22385), .IN2(n22384), .IN3(n22383), .IN4(n22382), 
        .QN(m1_data_o[14]) );
  AO22X1 U25521 ( .IN1(m0s14_data_i[15]), .IN2(n29256), .IN3(m0s10_data_i[15]), 
        .IN4(n29260), .Q(n22388) );
  AO22X1 U25522 ( .IN1(m0s11_data_i[15]), .IN2(n29259), .IN3(m0s8_data_i[15]), 
        .IN4(n29262), .Q(n22387) );
  AO22X1 U25523 ( .IN1(m0s2_data_i[15]), .IN2(n29268), .IN3(m0s9_data_i[15]), 
        .IN4(n29261), .Q(n22386) );
  NOR3X0 U25524 ( .IN1(n22388), .IN2(n22387), .IN3(n22386), .QN(n22396) );
  AO22X1 U25525 ( .IN1(m0s7_data_i[15]), .IN2(n29263), .IN3(m0s4_data_i[15]), 
        .IN4(n29266), .Q(n22392) );
  AO22X1 U25526 ( .IN1(m0s6_data_i[15]), .IN2(n29264), .IN3(m0s0_data_i[15]), 
        .IN4(n29271), .Q(n22391) );
  AO22X1 U25527 ( .IN1(m0s3_data_i[15]), .IN2(n29267), .IN3(m0s5_data_i[15]), 
        .IN4(n29265), .Q(n22390) );
  AO22X1 U25528 ( .IN1(m0s12_data_i[15]), .IN2(n29258), .IN3(m0s13_data_i[15]), 
        .IN4(n29257), .Q(n22389) );
  NOR4X0 U25529 ( .IN1(n22392), .IN2(n22391), .IN3(n22390), .IN4(n22389), .QN(
        n22395) );
  NAND2X0 U25530 ( .IN1(n29255), .IN2(n23103), .QN(n22394) );
  NAND2X0 U25531 ( .IN1(m0s1_data_i[15]), .IN2(n29269), .QN(n22393) );
  NAND4X0 U25532 ( .IN1(n22396), .IN2(n22395), .IN3(n22394), .IN4(n22393), 
        .QN(m1_data_o[15]) );
  OA22X1 U25533 ( .IN1(n23235), .IN2(n22830), .IN3(n22599), .IN4(n22834), .Q(
        n22409) );
  INVX0 U25534 ( .INP(n29262), .ZN(n22493) );
  OA22X1 U25535 ( .IN1(n22493), .IN2(n22397), .IN3(n23226), .IN4(n22837), .Q(
        n22408) );
  AO22X1 U25536 ( .IN1(n29257), .IN2(m0s13_data_i[17]), .IN3(n29259), .IN4(
        m0s11_data_i[17]), .Q(n22405) );
  AO22X1 U25537 ( .IN1(n29269), .IN2(m0s1_data_i[17]), .IN3(n29256), .IN4(
        m0s14_data_i[17]), .Q(n22404) );
  AO22X1 U25538 ( .IN1(n29266), .IN2(m0s4_data_i[17]), .IN3(n29265), .IN4(
        m0s5_data_i[17]), .Q(n22403) );
  AO22X1 U25539 ( .IN1(n29271), .IN2(m0s0_data_i[17]), .IN3(n29264), .IN4(
        m0s6_data_i[17]), .Q(n22399) );
  AO22X1 U25540 ( .IN1(n29268), .IN2(m0s2_data_i[17]), .IN3(n29261), .IN4(
        m0s9_data_i[17]), .Q(n22398) );
  NOR2X0 U25541 ( .IN1(n22399), .IN2(n22398), .QN(n22401) );
  NAND2X0 U25542 ( .IN1(n29263), .IN2(m0s7_data_i[17]), .QN(n22400) );
  NAND2X0 U25543 ( .IN1(n22401), .IN2(n22400), .QN(n22402) );
  NOR4X0 U25544 ( .IN1(n22405), .IN2(n22404), .IN3(n22403), .IN4(n22402), .QN(
        n22407) );
  NAND2X0 U25545 ( .IN1(s15_data_i[17]), .IN2(n22629), .QN(n22406) );
  NAND4X0 U25546 ( .IN1(n22409), .IN2(n22408), .IN3(n22407), .IN4(n22406), 
        .QN(m1_data_o[17]) );
  OA22X1 U25547 ( .IN1(n22584), .IN2(n22411), .IN3(n23226), .IN4(n22410), .Q(
        n22427) );
  OA22X1 U25548 ( .IN1(n23235), .IN2(n22413), .IN3(n23232), .IN4(n22412), .Q(
        n22426) );
  AO22X1 U25549 ( .IN1(n29268), .IN2(m0s2_data_i[18]), .IN3(n29269), .IN4(
        m0s1_data_i[18]), .Q(n22423) );
  AO22X1 U25550 ( .IN1(n29266), .IN2(m0s4_data_i[18]), .IN3(n29256), .IN4(
        m0s14_data_i[18]), .Q(n22422) );
  AO22X1 U25551 ( .IN1(n29259), .IN2(m0s11_data_i[18]), .IN3(n29260), .IN4(
        m0s10_data_i[18]), .Q(n22421) );
  OA22X1 U25552 ( .IN1(n22569), .IN2(n22415), .IN3(n23229), .IN4(n22414), .Q(
        n22419) );
  NAND2X0 U25553 ( .IN1(n29262), .IN2(m0s8_data_i[18]), .QN(n22418) );
  NAND2X0 U25554 ( .IN1(n29261), .IN2(m0s9_data_i[18]), .QN(n22417) );
  NAND2X0 U25555 ( .IN1(n29257), .IN2(m0s13_data_i[18]), .QN(n22416) );
  NAND4X0 U25556 ( .IN1(n22419), .IN2(n22418), .IN3(n22417), .IN4(n22416), 
        .QN(n22420) );
  NOR4X0 U25557 ( .IN1(n22423), .IN2(n22422), .IN3(n22421), .IN4(n22420), .QN(
        n22425) );
  NAND2X0 U25558 ( .IN1(s15_data_i[18]), .IN2(n22629), .QN(n22424) );
  NAND4X0 U25559 ( .IN1(n22427), .IN2(n22426), .IN3(n22425), .IN4(n22424), 
        .QN(m1_data_o[18]) );
  OA22X1 U25560 ( .IN1(n22582), .IN2(n22429), .IN3(n23241), .IN4(n22428), .Q(
        n22446) );
  OA22X1 U25561 ( .IN1(n23235), .IN2(n22431), .IN3(n22554), .IN4(n22430), .Q(
        n22445) );
  AO22X1 U25562 ( .IN1(n29262), .IN2(m0s8_data_i[19]), .IN3(n29269), .IN4(
        m0s1_data_i[19]), .Q(n22442) );
  AO22X1 U25563 ( .IN1(n29268), .IN2(m0s2_data_i[19]), .IN3(n29266), .IN4(
        m0s4_data_i[19]), .Q(n22441) );
  AO22X1 U25564 ( .IN1(n29264), .IN2(m0s6_data_i[19]), .IN3(n29259), .IN4(
        m0s11_data_i[19]), .Q(n22440) );
  OA22X1 U25565 ( .IN1(n22569), .IN2(n22433), .IN3(n22599), .IN4(n22432), .Q(
        n22438) );
  OA22X1 U25566 ( .IN1(n22584), .IN2(n22435), .IN3(n23226), .IN4(n22434), .Q(
        n22437) );
  NAND2X0 U25567 ( .IN1(n29265), .IN2(m0s5_data_i[19]), .QN(n22436) );
  NAND3X0 U25568 ( .IN1(n22438), .IN2(n22437), .IN3(n22436), .QN(n22439) );
  NOR4X0 U25569 ( .IN1(n22442), .IN2(n22441), .IN3(n22440), .IN4(n22439), .QN(
        n22444) );
  NAND2X0 U25570 ( .IN1(s15_data_i[19]), .IN2(n22629), .QN(n22443) );
  NAND4X0 U25571 ( .IN1(n22446), .IN2(n22445), .IN3(n22444), .IN4(n22443), 
        .QN(m1_data_o[19]) );
  OA22X1 U25572 ( .IN1(n23229), .IN2(n22448), .IN3(n22582), .IN4(n22447), .Q(
        n22465) );
  OA22X1 U25573 ( .IN1(n23223), .IN2(n22450), .IN3(n23226), .IN4(n22449), .Q(
        n22464) );
  AO22X1 U25574 ( .IN1(n29266), .IN2(m0s4_data_i[20]), .IN3(n29263), .IN4(
        m0s7_data_i[20]), .Q(n22461) );
  AO22X1 U25575 ( .IN1(n29269), .IN2(m0s1_data_i[20]), .IN3(n29260), .IN4(
        m0s10_data_i[20]), .Q(n22460) );
  AO22X1 U25576 ( .IN1(n29257), .IN2(m0s13_data_i[20]), .IN3(n29262), .IN4(
        m0s8_data_i[20]), .Q(n22459) );
  OA22X1 U25577 ( .IN1(n22620), .IN2(n22452), .IN3(n22569), .IN4(n22451), .Q(
        n22457) );
  OA22X1 U25578 ( .IN1(n23232), .IN2(n22454), .IN3(n23241), .IN4(n22453), .Q(
        n22456) );
  NAND2X0 U25579 ( .IN1(n29267), .IN2(m0s3_data_i[20]), .QN(n22455) );
  NAND3X0 U25580 ( .IN1(n22457), .IN2(n22456), .IN3(n22455), .QN(n22458) );
  NOR4X0 U25581 ( .IN1(n22461), .IN2(n22460), .IN3(n22459), .IN4(n22458), .QN(
        n22463) );
  NAND2X0 U25582 ( .IN1(s15_data_i[20]), .IN2(n22629), .QN(n22462) );
  NAND4X0 U25583 ( .IN1(n22465), .IN2(n22464), .IN3(n22463), .IN4(n22462), 
        .QN(m1_data_o[20]) );
  OA22X1 U25584 ( .IN1(n22569), .IN2(n22853), .IN3(n22567), .IN4(n22850), .Q(
        n22478) );
  OA22X1 U25585 ( .IN1(n22620), .IN2(n22856), .IN3(n23238), .IN4(n22466), .Q(
        n22477) );
  AO22X1 U25586 ( .IN1(n29264), .IN2(m0s6_data_i[21]), .IN3(n29260), .IN4(
        m0s10_data_i[21]), .Q(n22474) );
  AO22X1 U25587 ( .IN1(n29257), .IN2(m0s13_data_i[21]), .IN3(n29259), .IN4(
        m0s11_data_i[21]), .Q(n22473) );
  AO22X1 U25588 ( .IN1(n29267), .IN2(m0s3_data_i[21]), .IN3(n29265), .IN4(
        m0s5_data_i[21]), .Q(n22472) );
  AO22X1 U25589 ( .IN1(n29263), .IN2(m0s7_data_i[21]), .IN3(n29261), .IN4(
        m0s9_data_i[21]), .Q(n22468) );
  AO22X1 U25590 ( .IN1(n29262), .IN2(m0s8_data_i[21]), .IN3(n29256), .IN4(
        m0s14_data_i[21]), .Q(n22467) );
  NOR2X0 U25591 ( .IN1(n22468), .IN2(n22467), .QN(n22470) );
  NAND2X0 U25592 ( .IN1(n29258), .IN2(m0s12_data_i[21]), .QN(n22469) );
  NAND2X0 U25593 ( .IN1(n22470), .IN2(n22469), .QN(n22471) );
  NOR4X0 U25594 ( .IN1(n22474), .IN2(n22473), .IN3(n22472), .IN4(n22471), .QN(
        n22476) );
  NAND2X0 U25595 ( .IN1(s15_data_i[21]), .IN2(n22629), .QN(n22475) );
  NAND4X0 U25596 ( .IN1(n22478), .IN2(n22477), .IN3(n22476), .IN4(n22475), 
        .QN(m1_data_o[21]) );
  OA22X1 U25597 ( .IN1(n22493), .IN2(n22873), .IN3(n23226), .IN4(n22875), .Q(
        n22490) );
  OA22X1 U25598 ( .IN1(n22620), .IN2(n22870), .IN3(n23235), .IN4(n22871), .Q(
        n22489) );
  AO22X1 U25599 ( .IN1(n29271), .IN2(m0s0_data_i[22]), .IN3(n29269), .IN4(
        m0s1_data_i[22]), .Q(n22486) );
  AO22X1 U25600 ( .IN1(n29266), .IN2(m0s4_data_i[22]), .IN3(n29257), .IN4(
        m0s13_data_i[22]), .Q(n22485) );
  AO22X1 U25601 ( .IN1(n29263), .IN2(m0s7_data_i[22]), .IN3(n29261), .IN4(
        m0s9_data_i[22]), .Q(n22484) );
  AO22X1 U25602 ( .IN1(n29264), .IN2(m0s6_data_i[22]), .IN3(n29259), .IN4(
        m0s11_data_i[22]), .Q(n22480) );
  AO22X1 U25603 ( .IN1(n29265), .IN2(m0s5_data_i[22]), .IN3(n29260), .IN4(
        m0s10_data_i[22]), .Q(n22479) );
  NOR2X0 U25604 ( .IN1(n22480), .IN2(n22479), .QN(n22482) );
  NAND2X0 U25605 ( .IN1(n29256), .IN2(m0s14_data_i[22]), .QN(n22481) );
  NAND2X0 U25606 ( .IN1(n22482), .IN2(n22481), .QN(n22483) );
  NOR4X0 U25607 ( .IN1(n22486), .IN2(n22485), .IN3(n22484), .IN4(n22483), .QN(
        n22488) );
  NAND2X0 U25608 ( .IN1(s15_data_i[22]), .IN2(n22629), .QN(n22487) );
  NAND4X0 U25609 ( .IN1(n22490), .IN2(n22489), .IN3(n22488), .IN4(n22487), 
        .QN(m1_data_o[22]) );
  OA22X1 U25610 ( .IN1(n22493), .IN2(n22492), .IN3(n23238), .IN4(n22491), .Q(
        n22507) );
  OA22X1 U25611 ( .IN1(n22584), .IN2(n22495), .IN3(n22599), .IN4(n22494), .Q(
        n22506) );
  AO22X1 U25612 ( .IN1(n29267), .IN2(m0s3_data_i[23]), .IN3(n29265), .IN4(
        m0s5_data_i[23]), .Q(n22503) );
  AO22X1 U25613 ( .IN1(n29268), .IN2(m0s2_data_i[23]), .IN3(n29256), .IN4(
        m0s14_data_i[23]), .Q(n22502) );
  AO22X1 U25614 ( .IN1(n29271), .IN2(m0s0_data_i[23]), .IN3(n29257), .IN4(
        m0s13_data_i[23]), .Q(n22501) );
  AO22X1 U25615 ( .IN1(n29261), .IN2(m0s9_data_i[23]), .IN3(n29259), .IN4(
        m0s11_data_i[23]), .Q(n22497) );
  AO22X1 U25616 ( .IN1(n29264), .IN2(m0s6_data_i[23]), .IN3(n29258), .IN4(
        m0s12_data_i[23]), .Q(n22496) );
  NOR2X0 U25617 ( .IN1(n22497), .IN2(n22496), .QN(n22499) );
  NAND2X0 U25618 ( .IN1(n29266), .IN2(m0s4_data_i[23]), .QN(n22498) );
  NAND2X0 U25619 ( .IN1(n22499), .IN2(n22498), .QN(n22500) );
  NOR4X0 U25620 ( .IN1(n22503), .IN2(n22502), .IN3(n22501), .IN4(n22500), .QN(
        n22505) );
  NAND2X0 U25621 ( .IN1(s15_data_i[23]), .IN2(n22629), .QN(n22504) );
  NAND4X0 U25622 ( .IN1(n22507), .IN2(n22506), .IN3(n22505), .IN4(n22504), 
        .QN(m1_data_o[23]) );
  OA22X1 U25623 ( .IN1(n22554), .IN2(n22888), .IN3(n23241), .IN4(n22893), .Q(
        n22519) );
  OA22X1 U25624 ( .IN1(n22584), .IN2(n22891), .IN3(n23238), .IN4(n22896), .Q(
        n22518) );
  AO22X1 U25625 ( .IN1(n29271), .IN2(m0s0_data_i[24]), .IN3(n29265), .IN4(
        m0s5_data_i[24]), .Q(n22515) );
  AO22X1 U25626 ( .IN1(n29267), .IN2(m0s3_data_i[24]), .IN3(n29260), .IN4(
        m0s10_data_i[24]), .Q(n22514) );
  AO22X1 U25627 ( .IN1(n29261), .IN2(m0s9_data_i[24]), .IN3(n29259), .IN4(
        m0s11_data_i[24]), .Q(n22513) );
  AO22X1 U25628 ( .IN1(n29268), .IN2(m0s2_data_i[24]), .IN3(n29262), .IN4(
        m0s8_data_i[24]), .Q(n22509) );
  AO22X1 U25629 ( .IN1(n29266), .IN2(m0s4_data_i[24]), .IN3(n29264), .IN4(
        m0s6_data_i[24]), .Q(n22508) );
  NOR2X0 U25630 ( .IN1(n22509), .IN2(n22508), .QN(n22511) );
  NAND2X0 U25631 ( .IN1(n29258), .IN2(m0s12_data_i[24]), .QN(n22510) );
  NAND2X0 U25632 ( .IN1(n22511), .IN2(n22510), .QN(n22512) );
  NOR4X0 U25633 ( .IN1(n22515), .IN2(n22514), .IN3(n22513), .IN4(n22512), .QN(
        n22517) );
  NAND2X0 U25634 ( .IN1(s15_data_i[24]), .IN2(n22629), .QN(n22516) );
  NAND4X0 U25635 ( .IN1(n22519), .IN2(n22518), .IN3(n22517), .IN4(n22516), 
        .QN(m1_data_o[24]) );
  OA22X1 U25636 ( .IN1(n23235), .IN2(n22521), .IN3(n22582), .IN4(n22520), .Q(
        n22537) );
  OA22X1 U25637 ( .IN1(n22599), .IN2(n22523), .IN3(n23226), .IN4(n22522), .Q(
        n22536) );
  AO22X1 U25638 ( .IN1(n29268), .IN2(m0s2_data_i[25]), .IN3(n29264), .IN4(
        m0s6_data_i[25]), .Q(n22533) );
  AO22X1 U25639 ( .IN1(n29266), .IN2(m0s4_data_i[25]), .IN3(n29269), .IN4(
        m0s1_data_i[25]), .Q(n22532) );
  AO22X1 U25640 ( .IN1(n29271), .IN2(m0s0_data_i[25]), .IN3(n29259), .IN4(
        m0s11_data_i[25]), .Q(n22531) );
  OA22X1 U25641 ( .IN1(n23229), .IN2(n22525), .IN3(n23241), .IN4(n22524), .Q(
        n22529) );
  NAND2X0 U25642 ( .IN1(n29263), .IN2(m0s7_data_i[25]), .QN(n22528) );
  NAND2X0 U25643 ( .IN1(n29257), .IN2(m0s13_data_i[25]), .QN(n22527) );
  NAND2X0 U25644 ( .IN1(n29262), .IN2(m0s8_data_i[25]), .QN(n22526) );
  NAND4X0 U25645 ( .IN1(n22529), .IN2(n22528), .IN3(n22527), .IN4(n22526), 
        .QN(n22530) );
  NOR4X0 U25646 ( .IN1(n22533), .IN2(n22532), .IN3(n22531), .IN4(n22530), .QN(
        n22535) );
  NAND2X0 U25647 ( .IN1(s15_data_i[25]), .IN2(n22629), .QN(n22534) );
  NAND4X0 U25648 ( .IN1(n22537), .IN2(n22536), .IN3(n22535), .IN4(n22534), 
        .QN(m1_data_o[25]) );
  OA22X1 U25649 ( .IN1(n23232), .IN2(n22539), .IN3(n22493), .IN4(n22538), .Q(
        n22553) );
  OA22X1 U25650 ( .IN1(n23223), .IN2(n22541), .IN3(n22599), .IN4(n22540), .Q(
        n22552) );
  AO22X1 U25651 ( .IN1(n29268), .IN2(m0s2_data_i[26]), .IN3(n29266), .IN4(
        m0s4_data_i[26]), .Q(n22549) );
  AO22X1 U25652 ( .IN1(n29261), .IN2(m0s9_data_i[26]), .IN3(n29258), .IN4(
        m0s12_data_i[26]), .Q(n22548) );
  AO22X1 U25653 ( .IN1(n29271), .IN2(m0s0_data_i[26]), .IN3(n29256), .IN4(
        m0s14_data_i[26]), .Q(n22547) );
  AO22X1 U25654 ( .IN1(n29257), .IN2(m0s13_data_i[26]), .IN3(n29265), .IN4(
        m0s5_data_i[26]), .Q(n22543) );
  AO22X1 U25655 ( .IN1(n29267), .IN2(m0s3_data_i[26]), .IN3(n29269), .IN4(
        m0s1_data_i[26]), .Q(n22542) );
  NOR2X0 U25656 ( .IN1(n22543), .IN2(n22542), .QN(n22545) );
  NAND2X0 U25657 ( .IN1(n29263), .IN2(m0s7_data_i[26]), .QN(n22544) );
  NAND2X0 U25658 ( .IN1(n22545), .IN2(n22544), .QN(n22546) );
  NOR4X0 U25659 ( .IN1(n22549), .IN2(n22548), .IN3(n22547), .IN4(n22546), .QN(
        n22551) );
  NAND2X0 U25660 ( .IN1(s15_data_i[26]), .IN2(n22629), .QN(n22550) );
  NAND4X0 U25661 ( .IN1(n22553), .IN2(n22552), .IN3(n22551), .IN4(n22550), 
        .QN(m1_data_o[26]) );
  OA22X1 U25662 ( .IN1(n22554), .IN2(n22918), .IN3(n22493), .IN4(n22913), .Q(
        n22566) );
  OA22X1 U25663 ( .IN1(n22620), .IN2(n22916), .IN3(n23238), .IN4(n22910), .Q(
        n22565) );
  AO22X1 U25664 ( .IN1(n29260), .IN2(m0s10_data_i[27]), .IN3(n29256), .IN4(
        m0s14_data_i[27]), .Q(n22562) );
  AO22X1 U25665 ( .IN1(n29265), .IN2(m0s5_data_i[27]), .IN3(n29258), .IN4(
        m0s12_data_i[27]), .Q(n22561) );
  AO22X1 U25666 ( .IN1(n29266), .IN2(m0s4_data_i[27]), .IN3(n29263), .IN4(
        m0s7_data_i[27]), .Q(n22560) );
  AO22X1 U25667 ( .IN1(n29264), .IN2(m0s6_data_i[27]), .IN3(n29259), .IN4(
        m0s11_data_i[27]), .Q(n22556) );
  AO22X1 U25668 ( .IN1(n29267), .IN2(m0s3_data_i[27]), .IN3(n29261), .IN4(
        m0s9_data_i[27]), .Q(n22555) );
  NOR2X0 U25669 ( .IN1(n22556), .IN2(n22555), .QN(n22558) );
  NAND2X0 U25670 ( .IN1(n29271), .IN2(m0s0_data_i[27]), .QN(n22557) );
  NAND2X0 U25671 ( .IN1(n22558), .IN2(n22557), .QN(n22559) );
  NOR4X0 U25672 ( .IN1(n22562), .IN2(n22561), .IN3(n22560), .IN4(n22559), .QN(
        n22564) );
  NAND2X0 U25673 ( .IN1(s15_data_i[27]), .IN2(n22629), .QN(n22563) );
  NAND4X0 U25674 ( .IN1(n22566), .IN2(n22565), .IN3(n22564), .IN4(n22563), 
        .QN(m1_data_o[27]) );
  OA22X1 U25675 ( .IN1(n23238), .IN2(n22941), .IN3(n22582), .IN4(n22934), .Q(
        n22581) );
  OA22X1 U25676 ( .IN1(n22569), .IN2(n22568), .IN3(n22567), .IN4(n22938), .Q(
        n22580) );
  AO22X1 U25677 ( .IN1(n29257), .IN2(m0s13_data_i[28]), .IN3(n29259), .IN4(
        m0s11_data_i[28]), .Q(n22577) );
  AO22X1 U25678 ( .IN1(n29267), .IN2(m0s3_data_i[28]), .IN3(n29263), .IN4(
        m0s7_data_i[28]), .Q(n22576) );
  AO22X1 U25679 ( .IN1(n29262), .IN2(m0s8_data_i[28]), .IN3(n29260), .IN4(
        m0s10_data_i[28]), .Q(n22575) );
  OA22X1 U25680 ( .IN1(n23232), .IN2(n22940), .IN3(n23226), .IN4(n22935), .Q(
        n22573) );
  NAND2X0 U25681 ( .IN1(n29256), .IN2(m0s14_data_i[28]), .QN(n22572) );
  NAND2X0 U25682 ( .IN1(n29265), .IN2(m0s5_data_i[28]), .QN(n22571) );
  NAND2X0 U25683 ( .IN1(n29268), .IN2(m0s2_data_i[28]), .QN(n22570) );
  NAND4X0 U25684 ( .IN1(n22573), .IN2(n22572), .IN3(n22571), .IN4(n22570), 
        .QN(n22574) );
  NOR4X0 U25685 ( .IN1(n22577), .IN2(n22576), .IN3(n22575), .IN4(n22574), .QN(
        n22579) );
  NAND2X0 U25686 ( .IN1(s15_data_i[28]), .IN2(n22629), .QN(n22578) );
  NAND4X0 U25687 ( .IN1(n22581), .IN2(n22580), .IN3(n22579), .IN4(n22578), 
        .QN(m1_data_o[28]) );
  OA22X1 U25688 ( .IN1(n22584), .IN2(n22583), .IN3(n22582), .IN4(n22955), .Q(
        n22596) );
  OA22X1 U25689 ( .IN1(n23232), .IN2(n22963), .IN3(n23226), .IN4(n22957), .Q(
        n22595) );
  AO22X1 U25690 ( .IN1(n29267), .IN2(m0s3_data_i[29]), .IN3(n29269), .IN4(
        m0s1_data_i[29]), .Q(n22592) );
  AO22X1 U25691 ( .IN1(n29271), .IN2(m0s0_data_i[29]), .IN3(n29256), .IN4(
        m0s14_data_i[29]), .Q(n22591) );
  AO22X1 U25692 ( .IN1(n29268), .IN2(m0s2_data_i[29]), .IN3(n29262), .IN4(
        m0s8_data_i[29]), .Q(n22590) );
  AO22X1 U25693 ( .IN1(n29259), .IN2(m0s11_data_i[29]), .IN3(n29260), .IN4(
        m0s10_data_i[29]), .Q(n22586) );
  AO22X1 U25694 ( .IN1(n29266), .IN2(m0s4_data_i[29]), .IN3(n29257), .IN4(
        m0s13_data_i[29]), .Q(n22585) );
  NOR2X0 U25695 ( .IN1(n22586), .IN2(n22585), .QN(n22588) );
  NAND2X0 U25696 ( .IN1(n29265), .IN2(m0s5_data_i[29]), .QN(n22587) );
  NAND2X0 U25697 ( .IN1(n22588), .IN2(n22587), .QN(n22589) );
  NOR4X0 U25698 ( .IN1(n22592), .IN2(n22591), .IN3(n22590), .IN4(n22589), .QN(
        n22594) );
  NAND2X0 U25699 ( .IN1(s15_data_i[29]), .IN2(n22629), .QN(n22593) );
  NAND4X0 U25700 ( .IN1(n22596), .IN2(n22595), .IN3(n22594), .IN4(n22593), 
        .QN(m1_data_o[29]) );
  OA22X1 U25701 ( .IN1(n22599), .IN2(n22598), .IN3(n23241), .IN4(n22597), .Q(
        n22615) );
  OA22X1 U25702 ( .IN1(n23238), .IN2(n22601), .IN3(n23226), .IN4(n22600), .Q(
        n22614) );
  AO22X1 U25703 ( .IN1(n29271), .IN2(m0s0_data_i[30]), .IN3(n29259), .IN4(
        m0s11_data_i[30]), .Q(n22611) );
  AO22X1 U25704 ( .IN1(n29266), .IN2(m0s4_data_i[30]), .IN3(n29265), .IN4(
        m0s5_data_i[30]), .Q(n22610) );
  AO22X1 U25705 ( .IN1(n29267), .IN2(m0s3_data_i[30]), .IN3(n29261), .IN4(
        m0s9_data_i[30]), .Q(n22609) );
  OA22X1 U25706 ( .IN1(n22620), .IN2(n22603), .IN3(n22554), .IN4(n22602), .Q(
        n22607) );
  NAND2X0 U25707 ( .IN1(n29264), .IN2(m0s6_data_i[30]), .QN(n22606) );
  NAND2X0 U25708 ( .IN1(n29263), .IN2(m0s7_data_i[30]), .QN(n22605) );
  NAND2X0 U25709 ( .IN1(n29262), .IN2(m0s8_data_i[30]), .QN(n22604) );
  NAND4X0 U25710 ( .IN1(n22607), .IN2(n22606), .IN3(n22605), .IN4(n22604), 
        .QN(n22608) );
  NOR4X0 U25711 ( .IN1(n22611), .IN2(n22610), .IN3(n22609), .IN4(n22608), .QN(
        n22613) );
  NAND2X0 U25712 ( .IN1(s15_data_i[30]), .IN2(n22629), .QN(n22612) );
  NAND4X0 U25713 ( .IN1(n22615), .IN2(n22614), .IN3(n22613), .IN4(n22612), 
        .QN(m1_data_o[30]) );
  OA22X1 U25714 ( .IN1(n23235), .IN2(n22617), .IN3(n23229), .IN4(n22616), .Q(
        n22633) );
  OA22X1 U25715 ( .IN1(n22620), .IN2(n22619), .IN3(n22554), .IN4(n22618), .Q(
        n22632) );
  AO22X1 U25716 ( .IN1(n29266), .IN2(m0s4_data_i[31]), .IN3(n29261), .IN4(
        m0s9_data_i[31]), .Q(n22628) );
  AO22X1 U25717 ( .IN1(n29259), .IN2(m0s11_data_i[31]), .IN3(n29260), .IN4(
        m0s10_data_i[31]), .Q(n22627) );
  AO22X1 U25718 ( .IN1(n29271), .IN2(m0s0_data_i[31]), .IN3(n29256), .IN4(
        m0s14_data_i[31]), .Q(n22626) );
  AO22X1 U25719 ( .IN1(n29262), .IN2(m0s8_data_i[31]), .IN3(n29269), .IN4(
        m0s1_data_i[31]), .Q(n22622) );
  AO22X1 U25720 ( .IN1(n29264), .IN2(m0s6_data_i[31]), .IN3(n29258), .IN4(
        m0s12_data_i[31]), .Q(n22621) );
  NOR2X0 U25721 ( .IN1(n22622), .IN2(n22621), .QN(n22624) );
  NAND2X0 U25722 ( .IN1(n29263), .IN2(m0s7_data_i[31]), .QN(n22623) );
  NAND2X0 U25723 ( .IN1(n22624), .IN2(n22623), .QN(n22625) );
  NOR4X0 U25724 ( .IN1(n22628), .IN2(n22627), .IN3(n22626), .IN4(n22625), .QN(
        n22631) );
  NAND2X0 U25725 ( .IN1(s15_data_i[31]), .IN2(n22629), .QN(n22630) );
  NAND4X0 U25726 ( .IN1(n22633), .IN2(n22632), .IN3(n22631), .IN4(n22630), 
        .QN(m1_data_o[31]) );
  OA22X1 U25727 ( .IN1(n22635), .IN2(n22958), .IN3(n22634), .IN4(n22939), .Q(
        n22650) );
  OA22X1 U25728 ( .IN1(n22637), .IN2(n22937), .IN3(n22636), .IN4(n22933), .Q(
        n22649) );
  AO22X1 U25729 ( .IN1(m0s6_data_i[3]), .IN2(n29283), .IN3(m0s14_data_i[3]), 
        .IN4(n29275), .Q(n22645) );
  AO22X1 U25730 ( .IN1(m0s2_data_i[3]), .IN2(n29287), .IN3(m0s10_data_i[3]), 
        .IN4(n29279), .Q(n22644) );
  AO22X1 U25731 ( .IN1(m0s3_data_i[3]), .IN2(n29286), .IN3(m0s9_data_i[3]), 
        .IN4(n29280), .Q(n22643) );
  AO22X1 U25732 ( .IN1(m0s11_data_i[3]), .IN2(n29278), .IN3(m0s7_data_i[3]), 
        .IN4(n29282), .Q(n22639) );
  INVX0 U25733 ( .INP(n22960), .ZN(n29288) );
  AO22X1 U25734 ( .IN1(m0s1_data_i[3]), .IN2(n29288), .IN3(m0s8_data_i[3]), 
        .IN4(n29281), .Q(n22638) );
  NOR2X0 U25735 ( .IN1(n22639), .IN2(n22638), .QN(n22641) );
  NAND2X0 U25736 ( .IN1(m0s0_data_i[3]), .IN2(n29290), .QN(n22640) );
  NAND2X0 U25737 ( .IN1(n22641), .IN2(n22640), .QN(n22642) );
  NOR4X0 U25738 ( .IN1(n22645), .IN2(n22644), .IN3(n22643), .IN4(n22642), .QN(
        n22648) );
  NAND2X0 U25739 ( .IN1(n29274), .IN2(n22646), .QN(n22647) );
  NAND4X0 U25740 ( .IN1(n22650), .IN2(n22649), .IN3(n22648), .IN4(n22647), 
        .QN(m2_data_o[3]) );
  OA22X1 U25741 ( .IN1(n22652), .IN2(n22917), .IN3(n22651), .IN4(n22939), .Q(
        n22667) );
  OA22X1 U25742 ( .IN1(n22654), .IN2(n22958), .IN3(n22653), .IN4(n22933), .Q(
        n22666) );
  AO22X1 U25743 ( .IN1(m0s5_data_i[4]), .IN2(n29284), .IN3(m0s14_data_i[4]), 
        .IN4(n29275), .Q(n22662) );
  AO22X1 U25744 ( .IN1(m0s9_data_i[4]), .IN2(n29280), .IN3(m0s8_data_i[4]), 
        .IN4(n29281), .Q(n22661) );
  AO22X1 U25745 ( .IN1(m0s1_data_i[4]), .IN2(n29288), .IN3(m0s7_data_i[4]), 
        .IN4(n29282), .Q(n22660) );
  AO22X1 U25746 ( .IN1(m0s6_data_i[4]), .IN2(n29283), .IN3(m0s11_data_i[4]), 
        .IN4(n29278), .Q(n22656) );
  AO22X1 U25747 ( .IN1(m0s3_data_i[4]), .IN2(n29286), .IN3(m0s10_data_i[4]), 
        .IN4(n29279), .Q(n22655) );
  NOR2X0 U25748 ( .IN1(n22656), .IN2(n22655), .QN(n22658) );
  NAND2X0 U25749 ( .IN1(m0s0_data_i[4]), .IN2(n29290), .QN(n22657) );
  NAND2X0 U25750 ( .IN1(n22658), .IN2(n22657), .QN(n22659) );
  NOR4X0 U25751 ( .IN1(n22662), .IN2(n22661), .IN3(n22660), .IN4(n22659), .QN(
        n22665) );
  NAND2X0 U25752 ( .IN1(n29274), .IN2(n22663), .QN(n22664) );
  NAND4X0 U25753 ( .IN1(n22667), .IN2(n22666), .IN3(n22665), .IN4(n22664), 
        .QN(m2_data_o[4]) );
  OA22X1 U25754 ( .IN1(n22669), .IN2(n22917), .IN3(n22668), .IN4(n22954), .Q(
        n22684) );
  OA22X1 U25755 ( .IN1(n22671), .IN2(n22933), .IN3(n22670), .IN4(n22909), .Q(
        n22683) );
  AO22X1 U25756 ( .IN1(m0s10_data_i[5]), .IN2(n29279), .IN3(m0s4_data_i[5]), 
        .IN4(n29285), .Q(n22679) );
  AO22X1 U25757 ( .IN1(m0s5_data_i[5]), .IN2(n29284), .IN3(m0s9_data_i[5]), 
        .IN4(n29280), .Q(n22678) );
  AO22X1 U25758 ( .IN1(m0s6_data_i[5]), .IN2(n29283), .IN3(m0s12_data_i[5]), 
        .IN4(n29277), .Q(n22677) );
  AO22X1 U25759 ( .IN1(m0s1_data_i[5]), .IN2(n29288), .IN3(m0s11_data_i[5]), 
        .IN4(n29278), .Q(n22673) );
  AO22X1 U25760 ( .IN1(m0s0_data_i[5]), .IN2(n29290), .IN3(m0s14_data_i[5]), 
        .IN4(n29275), .Q(n22672) );
  NOR2X0 U25761 ( .IN1(n22673), .IN2(n22672), .QN(n22675) );
  NAND2X0 U25762 ( .IN1(m0s8_data_i[5]), .IN2(n29281), .QN(n22674) );
  NAND2X0 U25763 ( .IN1(n22675), .IN2(n22674), .QN(n22676) );
  NOR4X0 U25764 ( .IN1(n22679), .IN2(n22678), .IN3(n22677), .IN4(n22676), .QN(
        n22682) );
  NAND2X0 U25765 ( .IN1(n29274), .IN2(n22680), .QN(n22681) );
  NAND4X0 U25766 ( .IN1(n22684), .IN2(n22683), .IN3(n22682), .IN4(n22681), 
        .QN(m2_data_o[5]) );
  OA22X1 U25767 ( .IN1(n22686), .IN2(n22962), .IN3(n22685), .IN4(n22954), .Q(
        n22701) );
  OA22X1 U25768 ( .IN1(n22688), .IN2(n22914), .IN3(n22687), .IN4(n22933), .Q(
        n22700) );
  AO22X1 U25769 ( .IN1(m0s5_data_i[6]), .IN2(n29284), .IN3(m0s9_data_i[6]), 
        .IN4(n29280), .Q(n22696) );
  AO22X1 U25770 ( .IN1(m0s7_data_i[6]), .IN2(n29282), .IN3(m0s14_data_i[6]), 
        .IN4(n29275), .Q(n22695) );
  AO22X1 U25771 ( .IN1(m0s11_data_i[6]), .IN2(n29278), .IN3(m0s1_data_i[6]), 
        .IN4(n29288), .Q(n22694) );
  AO22X1 U25772 ( .IN1(m0s12_data_i[6]), .IN2(n29277), .IN3(m0s4_data_i[6]), 
        .IN4(n29285), .Q(n22690) );
  AO22X1 U25773 ( .IN1(m0s6_data_i[6]), .IN2(n29283), .IN3(m0s2_data_i[6]), 
        .IN4(n29287), .Q(n22689) );
  NOR2X0 U25774 ( .IN1(n22690), .IN2(n22689), .QN(n22692) );
  NAND2X0 U25775 ( .IN1(m0s0_data_i[6]), .IN2(n29290), .QN(n22691) );
  NAND2X0 U25776 ( .IN1(n22692), .IN2(n22691), .QN(n22693) );
  NOR4X0 U25777 ( .IN1(n22696), .IN2(n22695), .IN3(n22694), .IN4(n22693), .QN(
        n22699) );
  NAND2X0 U25778 ( .IN1(n29274), .IN2(n22697), .QN(n22698) );
  NAND4X0 U25779 ( .IN1(n22701), .IN2(n22700), .IN3(n22699), .IN4(n22698), 
        .QN(m2_data_o[6]) );
  OA22X1 U25780 ( .IN1(n22703), .IN2(n22854), .IN3(n22702), .IN4(n22917), .Q(
        n22718) );
  OA22X1 U25781 ( .IN1(n22705), .IN2(n22939), .IN3(n22704), .IN4(n22958), .Q(
        n22717) );
  AO22X1 U25782 ( .IN1(m0s7_data_i[7]), .IN2(n29282), .IN3(m0s14_data_i[7]), 
        .IN4(n29275), .Q(n22713) );
  AO22X1 U25783 ( .IN1(m0s9_data_i[7]), .IN2(n29280), .IN3(m0s8_data_i[7]), 
        .IN4(n29281), .Q(n22712) );
  AO22X1 U25784 ( .IN1(m0s11_data_i[7]), .IN2(n29278), .IN3(m0s13_data_i[7]), 
        .IN4(n29276), .Q(n22711) );
  AO22X1 U25785 ( .IN1(m0s5_data_i[7]), .IN2(n29284), .IN3(m0s10_data_i[7]), 
        .IN4(n29279), .Q(n22707) );
  AO22X1 U25786 ( .IN1(m0s6_data_i[7]), .IN2(n29283), .IN3(m0s3_data_i[7]), 
        .IN4(n29286), .Q(n22706) );
  NOR2X0 U25787 ( .IN1(n22707), .IN2(n22706), .QN(n22709) );
  NAND2X0 U25788 ( .IN1(m0s1_data_i[7]), .IN2(n29288), .QN(n22708) );
  NAND2X0 U25789 ( .IN1(n22709), .IN2(n22708), .QN(n22710) );
  NOR4X0 U25790 ( .IN1(n22713), .IN2(n22712), .IN3(n22711), .IN4(n22710), .QN(
        n22716) );
  NAND2X0 U25791 ( .IN1(n29274), .IN2(n22714), .QN(n22715) );
  NAND4X0 U25792 ( .IN1(n22718), .IN2(n22717), .IN3(n22716), .IN4(n22715), 
        .QN(m2_data_o[7]) );
  OA22X1 U25793 ( .IN1(n22720), .IN2(n22909), .IN3(n22719), .IN4(n22914), .Q(
        n22735) );
  OA22X1 U25794 ( .IN1(n22722), .IN2(n22960), .IN3(n22721), .IN4(n22854), .Q(
        n22734) );
  AO22X1 U25795 ( .IN1(m0s11_data_i[8]), .IN2(n29278), .IN3(m0s3_data_i[8]), 
        .IN4(n29286), .Q(n22730) );
  AO22X1 U25796 ( .IN1(m0s12_data_i[8]), .IN2(n29277), .IN3(m0s6_data_i[8]), 
        .IN4(n29283), .Q(n22729) );
  AO22X1 U25797 ( .IN1(m0s2_data_i[8]), .IN2(n29287), .IN3(m0s14_data_i[8]), 
        .IN4(n29275), .Q(n22728) );
  AO22X1 U25798 ( .IN1(m0s4_data_i[8]), .IN2(n29285), .IN3(m0s13_data_i[8]), 
        .IN4(n29276), .Q(n22724) );
  AO22X1 U25799 ( .IN1(m0s10_data_i[8]), .IN2(n29279), .IN3(m0s9_data_i[8]), 
        .IN4(n29280), .Q(n22723) );
  NOR2X0 U25800 ( .IN1(n22724), .IN2(n22723), .QN(n22726) );
  NAND2X0 U25801 ( .IN1(m0s5_data_i[8]), .IN2(n29284), .QN(n22725) );
  NAND2X0 U25802 ( .IN1(n22726), .IN2(n22725), .QN(n22727) );
  NOR4X0 U25803 ( .IN1(n22730), .IN2(n22729), .IN3(n22728), .IN4(n22727), .QN(
        n22733) );
  NAND2X0 U25804 ( .IN1(n29274), .IN2(n22731), .QN(n22732) );
  NAND4X0 U25805 ( .IN1(n22735), .IN2(n22734), .IN3(n22733), .IN4(n22732), 
        .QN(m2_data_o[8]) );
  OA22X1 U25806 ( .IN1(n22979), .IN2(n22958), .IN3(n22983), .IN4(n22937), .Q(
        n22748) );
  OA22X1 U25807 ( .IN1(n22984), .IN2(n22956), .IN3(n22736), .IN4(n22909), .Q(
        n22747) );
  AO22X1 U25808 ( .IN1(m0s11_data_i[9]), .IN2(n29278), .IN3(m0s0_data_i[9]), 
        .IN4(n29290), .Q(n22744) );
  AO22X1 U25809 ( .IN1(m0s10_data_i[9]), .IN2(n29279), .IN3(m0s6_data_i[9]), 
        .IN4(n29283), .Q(n22743) );
  AO22X1 U25810 ( .IN1(m0s1_data_i[9]), .IN2(n29288), .IN3(m0s14_data_i[9]), 
        .IN4(n29275), .Q(n22742) );
  AO22X1 U25811 ( .IN1(m0s3_data_i[9]), .IN2(n29286), .IN3(m0s8_data_i[9]), 
        .IN4(n29281), .Q(n22738) );
  AO22X1 U25812 ( .IN1(m0s2_data_i[9]), .IN2(n29287), .IN3(m0s13_data_i[9]), 
        .IN4(n29276), .Q(n22737) );
  NOR2X0 U25813 ( .IN1(n22738), .IN2(n22737), .QN(n22740) );
  NAND2X0 U25814 ( .IN1(m0s4_data_i[9]), .IN2(n29285), .QN(n22739) );
  NAND2X0 U25815 ( .IN1(n22740), .IN2(n22739), .QN(n22741) );
  NOR4X0 U25816 ( .IN1(n22744), .IN2(n22743), .IN3(n22742), .IN4(n22741), .QN(
        n22746) );
  NAND2X0 U25817 ( .IN1(n29274), .IN2(n22993), .QN(n22745) );
  NAND4X0 U25818 ( .IN1(n22748), .IN2(n22747), .IN3(n22746), .IN4(n22745), 
        .QN(m2_data_o[9]) );
  OA22X1 U25819 ( .IN1(n22750), .IN2(n22909), .IN3(n22749), .IN4(n22917), .Q(
        n22767) );
  OA22X1 U25820 ( .IN1(n22752), .IN2(n22954), .IN3(n22751), .IN4(n22962), .Q(
        n22766) );
  AO22X1 U25821 ( .IN1(m0s14_data_i[10]), .IN2(n29275), .IN3(m0s0_data_i[10]), 
        .IN4(n29290), .Q(n22762) );
  AO22X1 U25822 ( .IN1(m0s8_data_i[10]), .IN2(n29281), .IN3(m0s5_data_i[10]), 
        .IN4(n29284), .Q(n22761) );
  AO22X1 U25823 ( .IN1(m0s13_data_i[10]), .IN2(n29276), .IN3(m0s6_data_i[10]), 
        .IN4(n29283), .Q(n22760) );
  OA22X1 U25824 ( .IN1(n22754), .IN2(n22958), .IN3(n22753), .IN4(n22939), .Q(
        n22758) );
  NAND2X0 U25825 ( .IN1(m0s9_data_i[10]), .IN2(n29280), .QN(n22757) );
  NAND2X0 U25826 ( .IN1(m0s11_data_i[10]), .IN2(n29278), .QN(n22756) );
  NAND2X0 U25827 ( .IN1(m0s1_data_i[10]), .IN2(n29288), .QN(n22755) );
  NAND4X0 U25828 ( .IN1(n22758), .IN2(n22757), .IN3(n22756), .IN4(n22755), 
        .QN(n22759) );
  NOR4X0 U25829 ( .IN1(n22762), .IN2(n22761), .IN3(n22760), .IN4(n22759), .QN(
        n22765) );
  NAND2X0 U25830 ( .IN1(n29274), .IN2(n22763), .QN(n22764) );
  NAND4X0 U25831 ( .IN1(n22767), .IN2(n22766), .IN3(n22765), .IN4(n22764), 
        .QN(m2_data_o[10]) );
  OA22X1 U25832 ( .IN1(n23004), .IN2(n22964), .IN3(n23000), .IN4(n22914), .Q(
        n22779) );
  OA22X1 U25833 ( .IN1(n23002), .IN2(n22954), .IN3(n23001), .IN4(n22931), .Q(
        n22778) );
  AO22X1 U25834 ( .IN1(m0s4_data_i[11]), .IN2(n29285), .IN3(m0s10_data_i[11]), 
        .IN4(n29279), .Q(n22775) );
  AO22X1 U25835 ( .IN1(m0s1_data_i[11]), .IN2(n29288), .IN3(m0s2_data_i[11]), 
        .IN4(n29287), .Q(n22774) );
  AO22X1 U25836 ( .IN1(m0s12_data_i[11]), .IN2(n29277), .IN3(m0s7_data_i[11]), 
        .IN4(n29282), .Q(n22773) );
  AO22X1 U25837 ( .IN1(m0s14_data_i[11]), .IN2(n29275), .IN3(m0s0_data_i[11]), 
        .IN4(n29290), .Q(n22769) );
  AO22X1 U25838 ( .IN1(m0s13_data_i[11]), .IN2(n29276), .IN3(m0s9_data_i[11]), 
        .IN4(n29280), .Q(n22768) );
  NOR2X0 U25839 ( .IN1(n22769), .IN2(n22768), .QN(n22771) );
  NAND2X0 U25840 ( .IN1(m0s5_data_i[11]), .IN2(n29284), .QN(n22770) );
  NAND2X0 U25841 ( .IN1(n22771), .IN2(n22770), .QN(n22772) );
  NOR4X0 U25842 ( .IN1(n22775), .IN2(n22774), .IN3(n22773), .IN4(n22772), .QN(
        n22777) );
  NAND2X0 U25843 ( .IN1(n29274), .IN2(n23013), .QN(n22776) );
  NAND4X0 U25844 ( .IN1(n22779), .IN2(n22778), .IN3(n22777), .IN4(n22776), 
        .QN(m2_data_o[11]) );
  OA22X1 U25845 ( .IN1(n23018), .IN2(n22931), .IN3(n23025), .IN4(n22958), .Q(
        n22792) );
  OA22X1 U25846 ( .IN1(n22780), .IN2(n22933), .IN3(n23023), .IN4(n22954), .Q(
        n22791) );
  AO22X1 U25847 ( .IN1(m0s8_data_i[12]), .IN2(n29281), .IN3(m0s10_data_i[12]), 
        .IN4(n29279), .Q(n22788) );
  AO22X1 U25848 ( .IN1(m0s9_data_i[12]), .IN2(n29280), .IN3(m0s1_data_i[12]), 
        .IN4(n29288), .Q(n22787) );
  AO22X1 U25849 ( .IN1(m0s6_data_i[12]), .IN2(n29283), .IN3(m0s4_data_i[12]), 
        .IN4(n29285), .Q(n22786) );
  AO22X1 U25850 ( .IN1(m0s0_data_i[12]), .IN2(n29290), .IN3(m0s5_data_i[12]), 
        .IN4(n29284), .Q(n22782) );
  AO22X1 U25851 ( .IN1(m0s14_data_i[12]), .IN2(n29275), .IN3(m0s7_data_i[12]), 
        .IN4(n29282), .Q(n22781) );
  NOR2X0 U25852 ( .IN1(n22782), .IN2(n22781), .QN(n22784) );
  NAND2X0 U25853 ( .IN1(m0s2_data_i[12]), .IN2(n29287), .QN(n22783) );
  NAND2X0 U25854 ( .IN1(n22784), .IN2(n22783), .QN(n22785) );
  NOR4X0 U25855 ( .IN1(n22788), .IN2(n22787), .IN3(n22786), .IN4(n22785), .QN(
        n22790) );
  NAND2X0 U25856 ( .IN1(n29274), .IN2(n23034), .QN(n22789) );
  NAND4X0 U25857 ( .IN1(n22792), .IN2(n22791), .IN3(n22790), .IN4(n22789), 
        .QN(m2_data_o[12]) );
  OA22X1 U25858 ( .IN1(n23044), .IN2(n22962), .IN3(n23040), .IN4(n22917), .Q(
        n22805) );
  OA22X1 U25859 ( .IN1(n23042), .IN2(n22854), .IN3(n22793), .IN4(n22954), .Q(
        n22804) );
  AO22X1 U25860 ( .IN1(m0s7_data_i[13]), .IN2(n29282), .IN3(m0s1_data_i[13]), 
        .IN4(n29288), .Q(n22801) );
  AO22X1 U25861 ( .IN1(m0s8_data_i[13]), .IN2(n29281), .IN3(m0s12_data_i[13]), 
        .IN4(n29277), .Q(n22800) );
  AO22X1 U25862 ( .IN1(m0s4_data_i[13]), .IN2(n29285), .IN3(m0s9_data_i[13]), 
        .IN4(n29280), .Q(n22799) );
  AO22X1 U25863 ( .IN1(m0s6_data_i[13]), .IN2(n29283), .IN3(m0s11_data_i[13]), 
        .IN4(n29278), .Q(n22795) );
  AO22X1 U25864 ( .IN1(m0s13_data_i[13]), .IN2(n29276), .IN3(m0s5_data_i[13]), 
        .IN4(n29284), .Q(n22794) );
  NOR2X0 U25865 ( .IN1(n22795), .IN2(n22794), .QN(n22797) );
  NAND2X0 U25866 ( .IN1(m0s14_data_i[13]), .IN2(n29275), .QN(n22796) );
  NAND2X0 U25867 ( .IN1(n22797), .IN2(n22796), .QN(n22798) );
  NOR4X0 U25868 ( .IN1(n22801), .IN2(n22800), .IN3(n22799), .IN4(n22798), .QN(
        n22803) );
  NAND2X0 U25869 ( .IN1(n29274), .IN2(n23053), .QN(n22802) );
  NAND4X0 U25870 ( .IN1(n22805), .IN2(n22804), .IN3(n22803), .IN4(n22802), 
        .QN(m2_data_o[13]) );
  OA22X1 U25871 ( .IN1(n23066), .IN2(n22854), .IN3(n23064), .IN4(n22939), .Q(
        n22817) );
  OA22X1 U25872 ( .IN1(n23061), .IN2(n22960), .IN3(n23068), .IN4(n22931), .Q(
        n22816) );
  AO22X1 U25873 ( .IN1(m0s14_data_i[14]), .IN2(n29275), .IN3(m0s13_data_i[14]), 
        .IN4(n29276), .Q(n22813) );
  AO22X1 U25874 ( .IN1(m0s3_data_i[14]), .IN2(n29286), .IN3(m0s5_data_i[14]), 
        .IN4(n29284), .Q(n22812) );
  AO22X1 U25875 ( .IN1(m0s6_data_i[14]), .IN2(n29283), .IN3(m0s2_data_i[14]), 
        .IN4(n29287), .Q(n22811) );
  AO22X1 U25876 ( .IN1(m0s8_data_i[14]), .IN2(n29281), .IN3(m0s10_data_i[14]), 
        .IN4(n29279), .Q(n22807) );
  AO22X1 U25877 ( .IN1(m0s7_data_i[14]), .IN2(n29282), .IN3(m0s9_data_i[14]), 
        .IN4(n29280), .Q(n22806) );
  NOR2X0 U25878 ( .IN1(n22807), .IN2(n22806), .QN(n22809) );
  NAND2X0 U25879 ( .IN1(m0s12_data_i[14]), .IN2(n29277), .QN(n22808) );
  NAND2X0 U25880 ( .IN1(n22809), .IN2(n22808), .QN(n22810) );
  NOR4X0 U25881 ( .IN1(n22813), .IN2(n22812), .IN3(n22811), .IN4(n22810), .QN(
        n22815) );
  NAND2X0 U25882 ( .IN1(n29274), .IN2(n23078), .QN(n22814) );
  NAND4X0 U25883 ( .IN1(n22817), .IN2(n22816), .IN3(n22815), .IN4(n22814), 
        .QN(m2_data_o[14]) );
  OA22X1 U25884 ( .IN1(n23092), .IN2(n22914), .IN3(n23088), .IN4(n22958), .Q(
        n22829) );
  OA22X1 U25885 ( .IN1(n23090), .IN2(n22954), .IN3(n23094), .IN4(n22909), .Q(
        n22828) );
  AO22X1 U25886 ( .IN1(m0s14_data_i[15]), .IN2(n29275), .IN3(m0s9_data_i[15]), 
        .IN4(n29280), .Q(n22825) );
  AO22X1 U25887 ( .IN1(m0s10_data_i[15]), .IN2(n29279), .IN3(m0s4_data_i[15]), 
        .IN4(n29285), .Q(n22824) );
  AO22X1 U25888 ( .IN1(m0s11_data_i[15]), .IN2(n29278), .IN3(m0s0_data_i[15]), 
        .IN4(n29290), .Q(n22823) );
  AO22X1 U25889 ( .IN1(m0s5_data_i[15]), .IN2(n29284), .IN3(m0s13_data_i[15]), 
        .IN4(n29276), .Q(n22819) );
  AO22X1 U25890 ( .IN1(m0s2_data_i[15]), .IN2(n29287), .IN3(m0s1_data_i[15]), 
        .IN4(n29288), .Q(n22818) );
  NOR2X0 U25891 ( .IN1(n22819), .IN2(n22818), .QN(n22821) );
  NAND2X0 U25892 ( .IN1(m0s6_data_i[15]), .IN2(n29283), .QN(n22820) );
  NAND2X0 U25893 ( .IN1(n22821), .IN2(n22820), .QN(n22822) );
  NOR4X0 U25894 ( .IN1(n22825), .IN2(n22824), .IN3(n22823), .IN4(n22822), .QN(
        n22827) );
  NAND2X0 U25895 ( .IN1(n29274), .IN2(n23103), .QN(n22826) );
  NAND4X0 U25896 ( .IN1(n22829), .IN2(n22828), .IN3(n22827), .IN4(n22826), 
        .QN(m2_data_o[15]) );
  OA22X1 U25897 ( .IN1(n22909), .IN2(n22831), .IN3(n22954), .IN4(n22830), .Q(
        n22848) );
  OA22X1 U25898 ( .IN1(n22939), .IN2(n22833), .IN3(n22931), .IN4(n22832), .Q(
        n22847) );
  AO22X1 U25899 ( .IN1(n29288), .IN2(m0s1_data_i[17]), .IN3(n29275), .IN4(
        m0s14_data_i[17]), .Q(n22844) );
  AO22X1 U25900 ( .IN1(n29287), .IN2(m0s2_data_i[17]), .IN3(n29290), .IN4(
        m0s0_data_i[17]), .Q(n22843) );
  AO22X1 U25901 ( .IN1(n29283), .IN2(m0s6_data_i[17]), .IN3(n29284), .IN4(
        m0s5_data_i[17]), .Q(n22842) );
  OA22X1 U25902 ( .IN1(n22956), .IN2(n22835), .IN3(n22962), .IN4(n22834), .Q(
        n22840) );
  OA22X1 U25903 ( .IN1(n22958), .IN2(n22837), .IN3(n22933), .IN4(n22836), .Q(
        n22839) );
  NAND2X0 U25904 ( .IN1(n29281), .IN2(m0s8_data_i[17]), .QN(n22838) );
  NAND3X0 U25905 ( .IN1(n22840), .IN2(n22839), .IN3(n22838), .QN(n22841) );
  NOR4X0 U25906 ( .IN1(n22844), .IN2(n22843), .IN3(n22842), .IN4(n22841), .QN(
        n22846) );
  NAND2X0 U25907 ( .IN1(s15_data_i[17]), .IN2(n22973), .QN(n22845) );
  NAND4X0 U25908 ( .IN1(n22848), .IN2(n22847), .IN3(n22846), .IN4(n22845), 
        .QN(m2_data_o[17]) );
  OA22X1 U25909 ( .IN1(n22939), .IN2(n22850), .IN3(n22962), .IN4(n22849), .Q(
        n22868) );
  OA22X1 U25910 ( .IN1(n22958), .IN2(n22852), .IN3(n22937), .IN4(n22851), .Q(
        n22867) );
  AO22X1 U25911 ( .IN1(n29281), .IN2(m0s8_data_i[21]), .IN3(n29275), .IN4(
        m0s14_data_i[21]), .Q(n22864) );
  AO22X1 U25912 ( .IN1(n29276), .IN2(m0s13_data_i[21]), .IN3(n29286), .IN4(
        m0s3_data_i[21]), .Q(n22863) );
  AO22X1 U25913 ( .IN1(n29280), .IN2(m0s9_data_i[21]), .IN3(n29278), .IN4(
        m0s11_data_i[21]), .Q(n22862) );
  OA22X1 U25914 ( .IN1(n22964), .IN2(n22855), .IN3(n22854), .IN4(n22853), .Q(
        n22860) );
  OA22X1 U25915 ( .IN1(n22909), .IN2(n22857), .IN3(n22917), .IN4(n22856), .Q(
        n22859) );
  NAND2X0 U25916 ( .IN1(n29288), .IN2(m0s1_data_i[21]), .QN(n22858) );
  NAND3X0 U25917 ( .IN1(n22860), .IN2(n22859), .IN3(n22858), .QN(n22861) );
  NOR4X0 U25918 ( .IN1(n22864), .IN2(n22863), .IN3(n22862), .IN4(n22861), .QN(
        n22866) );
  NAND2X0 U25919 ( .IN1(s15_data_i[21]), .IN2(n22973), .QN(n22865) );
  NAND4X0 U25920 ( .IN1(n22868), .IN2(n22867), .IN3(n22866), .IN4(n22865), 
        .QN(m2_data_o[21]) );
  OA22X1 U25921 ( .IN1(n22917), .IN2(n22870), .IN3(n22962), .IN4(n22869), .Q(
        n22887) );
  OA22X1 U25922 ( .IN1(n22964), .IN2(n22872), .IN3(n22954), .IN4(n22871), .Q(
        n22886) );
  AO22X1 U25923 ( .IN1(n29280), .IN2(m0s9_data_i[22]), .IN3(n29284), .IN4(
        m0s5_data_i[22]), .Q(n22883) );
  AO22X1 U25924 ( .IN1(n29278), .IN2(m0s11_data_i[22]), .IN3(n29290), .IN4(
        m0s0_data_i[22]), .Q(n22882) );
  AO22X1 U25925 ( .IN1(n29288), .IN2(m0s1_data_i[22]), .IN3(n29275), .IN4(
        m0s14_data_i[22]), .Q(n22881) );
  OA22X1 U25926 ( .IN1(n22909), .IN2(n22874), .IN3(n22914), .IN4(n22873), .Q(
        n22879) );
  OA22X1 U25927 ( .IN1(n22939), .IN2(n22876), .IN3(n22958), .IN4(n22875), .Q(
        n22878) );
  NAND2X0 U25928 ( .IN1(n29276), .IN2(m0s13_data_i[22]), .QN(n22877) );
  NAND3X0 U25929 ( .IN1(n22879), .IN2(n22878), .IN3(n22877), .QN(n22880) );
  NOR4X0 U25930 ( .IN1(n22883), .IN2(n22882), .IN3(n22881), .IN4(n22880), .QN(
        n22885) );
  NAND2X0 U25931 ( .IN1(s15_data_i[22]), .IN2(n22973), .QN(n22884) );
  NAND4X0 U25932 ( .IN1(n22887), .IN2(n22886), .IN3(n22885), .IN4(n22884), 
        .QN(m2_data_o[22]) );
  OA22X1 U25933 ( .IN1(n22964), .IN2(n22889), .IN3(n22933), .IN4(n22888), .Q(
        n22907) );
  OA22X1 U25934 ( .IN1(n22909), .IN2(n22891), .IN3(n22917), .IN4(n22890), .Q(
        n22906) );
  AO22X1 U25935 ( .IN1(n29277), .IN2(m0s12_data_i[24]), .IN3(n29286), .IN4(
        m0s3_data_i[24]), .Q(n22903) );
  AO22X1 U25936 ( .IN1(n29280), .IN2(m0s9_data_i[24]), .IN3(n29281), .IN4(
        m0s8_data_i[24]), .Q(n22902) );
  AO22X1 U25937 ( .IN1(n29285), .IN2(m0s4_data_i[24]), .IN3(n29278), .IN4(
        m0s11_data_i[24]), .Q(n22901) );
  OA22X1 U25938 ( .IN1(n22894), .IN2(n22893), .IN3(n22962), .IN4(n22892), .Q(
        n22899) );
  OA22X1 U25939 ( .IN1(n22960), .IN2(n22896), .IN3(n22937), .IN4(n22895), .Q(
        n22898) );
  NAND2X0 U25940 ( .IN1(n29290), .IN2(m0s0_data_i[24]), .QN(n22897) );
  NAND3X0 U25941 ( .IN1(n22899), .IN2(n22898), .IN3(n22897), .QN(n22900) );
  NOR4X0 U25942 ( .IN1(n22903), .IN2(n22902), .IN3(n22901), .IN4(n22900), .QN(
        n22905) );
  NAND2X0 U25943 ( .IN1(s15_data_i[24]), .IN2(n22973), .QN(n22904) );
  NAND4X0 U25944 ( .IN1(n22907), .IN2(n22906), .IN3(n22905), .IN4(n22904), 
        .QN(m2_data_o[24]) );
  OA22X1 U25945 ( .IN1(n22960), .IN2(n22910), .IN3(n22909), .IN4(n22908), .Q(
        n22929) );
  OA22X1 U25946 ( .IN1(n22954), .IN2(n22912), .IN3(n22962), .IN4(n22911), .Q(
        n22928) );
  AO22X1 U25947 ( .IN1(n29284), .IN2(m0s5_data_i[27]), .IN3(n29275), .IN4(
        m0s14_data_i[27]), .Q(n22925) );
  AO22X1 U25948 ( .IN1(n29283), .IN2(m0s6_data_i[27]), .IN3(n29280), .IN4(
        m0s9_data_i[27]), .Q(n22924) );
  AO22X1 U25949 ( .IN1(n29285), .IN2(m0s4_data_i[27]), .IN3(n29278), .IN4(
        m0s11_data_i[27]), .Q(n22923) );
  OA22X1 U25950 ( .IN1(n22958), .IN2(n22915), .IN3(n22914), .IN4(n22913), .Q(
        n22921) );
  OA22X1 U25951 ( .IN1(n22933), .IN2(n22918), .IN3(n22917), .IN4(n22916), .Q(
        n22920) );
  NAND2X0 U25952 ( .IN1(n29290), .IN2(m0s0_data_i[27]), .QN(n22919) );
  NAND3X0 U25953 ( .IN1(n22921), .IN2(n22920), .IN3(n22919), .QN(n22922) );
  NOR4X0 U25954 ( .IN1(n22925), .IN2(n22924), .IN3(n22923), .IN4(n22922), .QN(
        n22927) );
  NAND2X0 U25955 ( .IN1(s15_data_i[27]), .IN2(n22973), .QN(n22926) );
  NAND4X0 U25956 ( .IN1(n22929), .IN2(n22928), .IN3(n22927), .IN4(n22926), 
        .QN(m2_data_o[27]) );
  OA22X1 U25957 ( .IN1(n22933), .IN2(n22932), .IN3(n22931), .IN4(n22930), .Q(
        n22952) );
  OA22X1 U25958 ( .IN1(n22958), .IN2(n22935), .IN3(n22956), .IN4(n22934), .Q(
        n22951) );
  AO22X1 U25959 ( .IN1(n29281), .IN2(m0s8_data_i[28]), .IN3(n29286), .IN4(
        m0s3_data_i[28]), .Q(n22948) );
  AO22X1 U25960 ( .IN1(n29282), .IN2(m0s7_data_i[28]), .IN3(n29287), .IN4(
        m0s2_data_i[28]), .Q(n22947) );
  AO22X1 U25961 ( .IN1(n29275), .IN2(m0s14_data_i[28]), .IN3(n29279), .IN4(
        m0s10_data_i[28]), .Q(n22946) );
  OA22X1 U25962 ( .IN1(n22939), .IN2(n22938), .IN3(n22937), .IN4(n22936), .Q(
        n22944) );
  OA22X1 U25963 ( .IN1(n22960), .IN2(n22941), .IN3(n22964), .IN4(n22940), .Q(
        n22943) );
  NAND2X0 U25964 ( .IN1(n29290), .IN2(m0s0_data_i[28]), .QN(n22942) );
  NAND3X0 U25965 ( .IN1(n22944), .IN2(n22943), .IN3(n22942), .QN(n22945) );
  NOR4X0 U25966 ( .IN1(n22948), .IN2(n22947), .IN3(n22946), .IN4(n22945), .QN(
        n22950) );
  NAND2X0 U25967 ( .IN1(s15_data_i[28]), .IN2(n22973), .QN(n22949) );
  NAND4X0 U25968 ( .IN1(n22952), .IN2(n22951), .IN3(n22950), .IN4(n22949), 
        .QN(m2_data_o[28]) );
  OA22X1 U25969 ( .IN1(n22956), .IN2(n22955), .IN3(n22954), .IN4(n22953), .Q(
        n22977) );
  OA22X1 U25970 ( .IN1(n22960), .IN2(n22959), .IN3(n22958), .IN4(n22957), .Q(
        n22976) );
  AO22X1 U25971 ( .IN1(n29285), .IN2(m0s4_data_i[29]), .IN3(n29275), .IN4(
        m0s14_data_i[29]), .Q(n22972) );
  AO22X1 U25972 ( .IN1(n29282), .IN2(m0s7_data_i[29]), .IN3(n29281), .IN4(
        m0s8_data_i[29]), .Q(n22971) );
  AO22X1 U25973 ( .IN1(n29278), .IN2(m0s11_data_i[29]), .IN3(n29290), .IN4(
        m0s0_data_i[29]), .Q(n22970) );
  OA22X1 U25974 ( .IN1(n22964), .IN2(n22963), .IN3(n22962), .IN4(n22961), .Q(
        n22968) );
  NAND2X0 U25975 ( .IN1(n29284), .IN2(m0s5_data_i[29]), .QN(n22967) );
  NAND2X0 U25976 ( .IN1(n29287), .IN2(m0s2_data_i[29]), .QN(n22966) );
  NAND2X0 U25977 ( .IN1(n29276), .IN2(m0s13_data_i[29]), .QN(n22965) );
  NAND4X0 U25978 ( .IN1(n22968), .IN2(n22967), .IN3(n22966), .IN4(n22965), 
        .QN(n22969) );
  NOR4X0 U25979 ( .IN1(n22972), .IN2(n22971), .IN3(n22970), .IN4(n22969), .QN(
        n22975) );
  NAND2X0 U25980 ( .IN1(s15_data_i[29]), .IN2(n22973), .QN(n22974) );
  NAND4X0 U25981 ( .IN1(n22977), .IN2(n22976), .IN3(n22975), .IN4(n22974), 
        .QN(m2_data_o[29]) );
  OA22X1 U25982 ( .IN1(n22979), .IN2(n23087), .IN3(n22978), .IN4(n23091), .Q(
        n22997) );
  OA22X1 U25983 ( .IN1(n22981), .IN2(n23089), .IN3(n22980), .IN4(n23063), .Q(
        n22996) );
  AO22X1 U25984 ( .IN1(m0s10_data_i[9]), .IN2(n29298), .IN3(m0s14_data_i[9]), 
        .IN4(n29294), .Q(n22992) );
  AO22X1 U25985 ( .IN1(m0s2_data_i[9]), .IN2(n29306), .IN3(m0s1_data_i[9]), 
        .IN4(n29307), .Q(n22991) );
  AO22X1 U25986 ( .IN1(m0s13_data_i[9]), .IN2(n29295), .IN3(m0s11_data_i[9]), 
        .IN4(n29297), .Q(n22990) );
  OA22X1 U25987 ( .IN1(n22984), .IN2(n23021), .IN3(n22983), .IN4(n22982), .Q(
        n22988) );
  NAND2X0 U25988 ( .IN1(m0s7_data_i[9]), .IN2(n29301), .QN(n22987) );
  NAND2X0 U25989 ( .IN1(m0s6_data_i[9]), .IN2(n29302), .QN(n22986) );
  NAND2X0 U25990 ( .IN1(m0s0_data_i[9]), .IN2(n29309), .QN(n22985) );
  NAND4X0 U25991 ( .IN1(n22988), .IN2(n22987), .IN3(n22986), .IN4(n22985), 
        .QN(n22989) );
  NOR4X0 U25992 ( .IN1(n22992), .IN2(n22991), .IN3(n22990), .IN4(n22989), .QN(
        n22995) );
  NAND2X0 U25993 ( .IN1(n29293), .IN2(n22993), .QN(n22994) );
  NAND4X0 U25994 ( .IN1(n22997), .IN2(n22996), .IN3(n22995), .IN4(n22994), 
        .QN(m3_data_o[9]) );
  OA22X1 U25995 ( .IN1(n22999), .IN2(n23069), .IN3(n22998), .IN4(n23063), .Q(
        n23017) );
  OA22X1 U25996 ( .IN1(n23001), .IN2(n23067), .IN3(n23000), .IN4(n23091), .Q(
        n23016) );
  AO22X1 U25997 ( .IN1(m0s9_data_i[11]), .IN2(n29299), .IN3(m0s5_data_i[11]), 
        .IN4(n29303), .Q(n23012) );
  AO22X1 U25998 ( .IN1(m0s2_data_i[11]), .IN2(n29306), .IN3(m0s0_data_i[11]), 
        .IN4(n29309), .Q(n23011) );
  AO22X1 U25999 ( .IN1(m0s12_data_i[11]), .IN2(n29296), .IN3(m0s1_data_i[11]), 
        .IN4(n29307), .Q(n23010) );
  OA22X1 U26000 ( .IN1(n23004), .IN2(n23003), .IN3(n23002), .IN4(n23089), .Q(
        n23008) );
  NAND2X0 U26001 ( .IN1(m0s13_data_i[11]), .IN2(n29295), .QN(n23007) );
  NAND2X0 U26002 ( .IN1(m0s7_data_i[11]), .IN2(n29301), .QN(n23006) );
  NAND2X0 U26003 ( .IN1(m0s10_data_i[11]), .IN2(n29298), .QN(n23005) );
  NAND4X0 U26004 ( .IN1(n23008), .IN2(n23007), .IN3(n23006), .IN4(n23005), 
        .QN(n23009) );
  NOR4X0 U26005 ( .IN1(n23012), .IN2(n23011), .IN3(n23010), .IN4(n23009), .QN(
        n23015) );
  NAND2X0 U26006 ( .IN1(n29293), .IN2(n23013), .QN(n23014) );
  NAND4X0 U26007 ( .IN1(n23017), .IN2(n23016), .IN3(n23015), .IN4(n23014), 
        .QN(m3_data_o[11]) );
  OA22X1 U26008 ( .IN1(n23019), .IN2(n23065), .IN3(n23018), .IN4(n23067), .Q(
        n23038) );
  OA22X1 U26009 ( .IN1(n23022), .IN2(n23021), .IN3(n23020), .IN4(n23085), .Q(
        n23037) );
  AO22X1 U26010 ( .IN1(m0s8_data_i[12]), .IN2(n29300), .IN3(m0s10_data_i[12]), 
        .IN4(n29298), .Q(n23033) );
  AO22X1 U26011 ( .IN1(m0s4_data_i[12]), .IN2(n29304), .IN3(m0s5_data_i[12]), 
        .IN4(n29303), .Q(n23032) );
  AO22X1 U26012 ( .IN1(m0s7_data_i[12]), .IN2(n29301), .IN3(m0s6_data_i[12]), 
        .IN4(n29302), .Q(n23031) );
  OA22X1 U26013 ( .IN1(n23024), .IN2(n23069), .IN3(n23023), .IN4(n23089), .Q(
        n23029) );
  OA22X1 U26014 ( .IN1(n23026), .IN2(n23059), .IN3(n23025), .IN4(n23087), .Q(
        n23028) );
  NAND2X0 U26015 ( .IN1(m0s13_data_i[12]), .IN2(n29295), .QN(n23027) );
  NAND3X0 U26016 ( .IN1(n23029), .IN2(n23028), .IN3(n23027), .QN(n23030) );
  NOR4X0 U26017 ( .IN1(n23033), .IN2(n23032), .IN3(n23031), .IN4(n23030), .QN(
        n23036) );
  NAND2X0 U26018 ( .IN1(n29293), .IN2(n23034), .QN(n23035) );
  NAND4X0 U26019 ( .IN1(n23038), .IN2(n23037), .IN3(n23036), .IN4(n23035), 
        .QN(m3_data_o[12]) );
  OA22X1 U26020 ( .IN1(n23040), .IN2(n23059), .IN3(n23039), .IN4(n23069), .Q(
        n23057) );
  OA22X1 U26021 ( .IN1(n23042), .IN2(n23065), .IN3(n23041), .IN4(n23067), .Q(
        n23056) );
  AO22X1 U26022 ( .IN1(m0s4_data_i[13]), .IN2(n29304), .IN3(m0s3_data_i[13]), 
        .IN4(n29305), .Q(n23052) );
  AO22X1 U26023 ( .IN1(m0s6_data_i[13]), .IN2(n29302), .IN3(m0s1_data_i[13]), 
        .IN4(n29307), .Q(n23051) );
  AO22X1 U26024 ( .IN1(m0s7_data_i[13]), .IN2(n29301), .IN3(m0s12_data_i[13]), 
        .IN4(n29296), .Q(n23050) );
  OA22X1 U26025 ( .IN1(n23044), .IN2(n23083), .IN3(n23043), .IN4(n23021), .Q(
        n23048) );
  NAND2X0 U26026 ( .IN1(m0s5_data_i[13]), .IN2(n29303), .QN(n23047) );
  NAND2X0 U26027 ( .IN1(m0s13_data_i[13]), .IN2(n29295), .QN(n23046) );
  NAND2X0 U26028 ( .IN1(m0s8_data_i[13]), .IN2(n29300), .QN(n23045) );
  NAND4X0 U26029 ( .IN1(n23048), .IN2(n23047), .IN3(n23046), .IN4(n23045), 
        .QN(n23049) );
  NOR4X0 U26030 ( .IN1(n23052), .IN2(n23051), .IN3(n23050), .IN4(n23049), .QN(
        n23055) );
  NAND2X0 U26031 ( .IN1(n29293), .IN2(n23053), .QN(n23054) );
  NAND4X0 U26032 ( .IN1(n23057), .IN2(n23056), .IN3(n23055), .IN4(n23054), 
        .QN(m3_data_o[13]) );
  OA22X1 U26033 ( .IN1(n23060), .IN2(n23059), .IN3(n23058), .IN4(n23021), .Q(
        n23082) );
  OA22X1 U26034 ( .IN1(n23062), .IN2(n23091), .IN3(n23061), .IN4(n23085), .Q(
        n23081) );
  AO22X1 U26035 ( .IN1(m0s3_data_i[14]), .IN2(n29305), .IN3(m0s13_data_i[14]), 
        .IN4(n29295), .Q(n23077) );
  AO22X1 U26036 ( .IN1(m0s6_data_i[14]), .IN2(n29302), .IN3(m0s5_data_i[14]), 
        .IN4(n29303), .Q(n23076) );
  AO22X1 U26037 ( .IN1(m0s7_data_i[14]), .IN2(n29301), .IN3(m0s12_data_i[14]), 
        .IN4(n29296), .Q(n23075) );
  OA22X1 U26038 ( .IN1(n23066), .IN2(n23065), .IN3(n23064), .IN4(n23063), .Q(
        n23073) );
  OA22X1 U26039 ( .IN1(n23070), .IN2(n23069), .IN3(n23068), .IN4(n23067), .Q(
        n23072) );
  NAND2X0 U26040 ( .IN1(m0s10_data_i[14]), .IN2(n29298), .QN(n23071) );
  NAND3X0 U26041 ( .IN1(n23073), .IN2(n23072), .IN3(n23071), .QN(n23074) );
  NOR4X0 U26042 ( .IN1(n23077), .IN2(n23076), .IN3(n23075), .IN4(n23074), .QN(
        n23080) );
  NAND2X0 U26043 ( .IN1(n29293), .IN2(n23078), .QN(n23079) );
  NAND4X0 U26044 ( .IN1(n23082), .IN2(n23081), .IN3(n23080), .IN4(n23079), 
        .QN(m3_data_o[14]) );
  OA22X1 U26045 ( .IN1(n23086), .IN2(n23085), .IN3(n23084), .IN4(n23083), .Q(
        n23107) );
  OA22X1 U26046 ( .IN1(n23090), .IN2(n23089), .IN3(n23088), .IN4(n23087), .Q(
        n23106) );
  AO22X1 U26047 ( .IN1(m0s2_data_i[15]), .IN2(n29306), .IN3(m0s11_data_i[15]), 
        .IN4(n29297), .Q(n23102) );
  AO22X1 U26048 ( .IN1(m0s6_data_i[15]), .IN2(n29302), .IN3(m0s0_data_i[15]), 
        .IN4(n29309), .Q(n23101) );
  AO22X1 U26049 ( .IN1(m0s9_data_i[15]), .IN2(n29299), .IN3(m0s13_data_i[15]), 
        .IN4(n29295), .Q(n23100) );
  OA22X1 U26050 ( .IN1(n23094), .IN2(n23093), .IN3(n23092), .IN4(n23091), .Q(
        n23098) );
  NAND2X0 U26051 ( .IN1(m0s4_data_i[15]), .IN2(n29304), .QN(n23097) );
  NAND2X0 U26052 ( .IN1(m0s5_data_i[15]), .IN2(n29303), .QN(n23096) );
  NAND2X0 U26053 ( .IN1(m0s14_data_i[15]), .IN2(n29294), .QN(n23095) );
  NAND4X0 U26054 ( .IN1(n23098), .IN2(n23097), .IN3(n23096), .IN4(n23095), 
        .QN(n23099) );
  NOR4X0 U26055 ( .IN1(n23102), .IN2(n23101), .IN3(n23100), .IN4(n23099), .QN(
        n23105) );
  NAND2X0 U26056 ( .IN1(n29293), .IN2(n23103), .QN(n23104) );
  NAND4X0 U26057 ( .IN1(n23107), .IN2(n23106), .IN3(n23105), .IN4(n23104), 
        .QN(m3_data_o[15]) );
  NOR2X0 U26058 ( .IN1(\rf/rf_ack ), .IN2(n23445), .QN(\rf/N19 ) );
  INVX0 U26059 ( .INP(m4s0_we), .ZN(n28122) );
  INVX0 U26060 ( .INP(m6s0_we), .ZN(n28127) );
  OA22X1 U26061 ( .IN1(n23836), .IN2(n28122), .IN3(n23833), .IN4(n28127), .Q(
        n23111) );
  INVX0 U26062 ( .INP(m0s0_we), .ZN(n28124) );
  INVX0 U26063 ( .INP(m5s0_we), .ZN(n28125) );
  OA22X1 U26064 ( .IN1(n23823), .IN2(n28124), .IN3(n23832), .IN4(n28125), .Q(
        n23110) );
  INVX0 U26065 ( .INP(m1s0_we), .ZN(n28128) );
  INVX0 U26066 ( .INP(m2s0_we), .ZN(n28123) );
  OA22X1 U26067 ( .IN1(n23818), .IN2(n28128), .IN3(n23817), .IN4(n28123), .Q(
        n23109) );
  INVX0 U26068 ( .INP(m3s0_we), .ZN(n28126) );
  INVX0 U26069 ( .INP(m7s0_we), .ZN(n28121) );
  OA22X1 U26070 ( .IN1(n23835), .IN2(n28126), .IN3(n23824), .IN4(n28121), .Q(
        n23108) );
  NAND4X0 U26071 ( .IN1(n23111), .IN2(n23110), .IN3(n23109), .IN4(n23108), 
        .QN(s15_we_o) );
  AND3X1 U26072 ( .IN1(n23501), .IN2(n34379), .IN3(s15_we_o), .Q(\rf/N18 ) );
  OR2X1 U26073 ( .IN1(n23113), .IN2(n23112), .Q(n23209) );
  NOR2X0 U26074 ( .IN1(n23114), .IN2(n23209), .QN(n29002) );
  NAND2X0 U26075 ( .IN1(n29249), .IN2(n29002), .QN(n27498) );
  OR2X1 U26076 ( .IN1(n23116), .IN2(n23115), .Q(n23248) );
  NOR2X0 U26077 ( .IN1(n23117), .IN2(n23248), .QN(n29130) );
  NAND2X0 U26078 ( .IN1(n29242), .IN2(n29130), .QN(n25373) );
  OA22X1 U26079 ( .IN1(n27498), .IN2(n23214), .IN3(n25373), .IN4(n23253), .Q(
        n23177) );
  OR2X1 U26080 ( .IN1(n23119), .IN2(n23118), .Q(n23242) );
  NOR2X0 U26081 ( .IN1(n23120), .IN2(n23242), .QN(n29038) );
  NAND2X0 U26082 ( .IN1(n29247), .IN2(n29038), .QN(n26892) );
  OR2X1 U26083 ( .IN1(n23122), .IN2(n23121), .Q(n23244) );
  NOR2X0 U26084 ( .IN1(n23123), .IN2(n23244), .QN(n29120) );
  NAND2X0 U26085 ( .IN1(n29243), .IN2(n29120), .QN(n25672) );
  OA22X1 U26086 ( .IN1(n26892), .IN2(n23247), .IN3(n25672), .IN4(n23246), .Q(
        n23176) );
  NOR2X0 U26087 ( .IN1(n23125), .IN2(n23124), .QN(n23239) );
  AND2X1 U26088 ( .IN1(n23239), .IN2(n23126), .Q(n29218) );
  INVX0 U26089 ( .INP(n29218), .ZN(n24131) );
  NOR2X0 U26090 ( .IN1(n23127), .IN2(n24131), .QN(n23847) );
  NOR2X0 U26091 ( .IN1(n23129), .IN2(n23128), .QN(n23211) );
  AND2X1 U26092 ( .IN1(n23211), .IN2(n23130), .Q(n29202) );
  INVX0 U26093 ( .INP(n29202), .ZN(n24392) );
  NOR2X0 U26094 ( .IN1(n23131), .IN2(n24392), .QN(n23191) );
  AO22X1 U26095 ( .IN1(n23847), .IN2(s14_ack_i), .IN3(n23191), .IN4(s13_ack_i), 
        .Q(n23173) );
  NOR2X0 U26096 ( .IN1(n23133), .IN2(n23132), .QN(n23228) );
  AND2X1 U26097 ( .IN1(n23134), .IN2(n23228), .Q(n29066) );
  INVX0 U26098 ( .INP(n29066), .ZN(n26879) );
  NOR2X0 U26099 ( .IN1(n23135), .IN2(n26879), .QN(n26588) );
  NOR2X0 U26100 ( .IN1(n23137), .IN2(n23136), .QN(n23231) );
  AND2X1 U26101 ( .IN1(n23138), .IN2(n23231), .Q(n29081) );
  INVX0 U26102 ( .INP(n29081), .ZN(n26559) );
  NOR2X0 U26103 ( .IN1(n23139), .IN2(n26559), .QN(n23204) );
  AO22X1 U26104 ( .IN1(n26588), .IN2(s5_ack_i), .IN3(n23204), .IN4(s6_ack_i), 
        .Q(n23172) );
  NOR2X0 U26105 ( .IN1(n23141), .IN2(n23140), .QN(n23237) );
  AND2X1 U26106 ( .IN1(n23142), .IN2(n23237), .Q(n28984) );
  INVX0 U26107 ( .INP(n28984), .ZN(n28098) );
  NOR2X0 U26108 ( .IN1(n22178), .IN2(n28098), .QN(n27807) );
  NOR2X0 U26109 ( .IN1(n23144), .IN2(n23143), .QN(n23216) );
  AND2X1 U26110 ( .IN1(n23145), .IN2(n23216), .Q(n29099) );
  NAND2X0 U26111 ( .IN1(n29244), .IN2(n29099), .QN(n25978) );
  INVX0 U26112 ( .INP(n25978), .ZN(n23196) );
  AO22X1 U26113 ( .IN1(n27807), .IN2(s1_ack_i), .IN3(n23196), .IN4(s7_ack_i), 
        .Q(n23171) );
  NOR2X0 U26114 ( .IN1(n23147), .IN2(n23146), .QN(n23222) );
  AND2X1 U26115 ( .IN1(n23148), .IN2(n23222), .Q(n29165) );
  INVX0 U26116 ( .INP(n29165), .ZN(n25053) );
  NOR2X0 U26117 ( .IN1(n23149), .IN2(n25053), .QN(n24759) );
  NOR2X0 U26118 ( .IN1(n23151), .IN2(n23150), .QN(n23225) );
  AND2X1 U26119 ( .IN1(n23152), .IN2(n23225), .Q(n29191) );
  INVX0 U26120 ( .INP(n29191), .ZN(n24737) );
  NOR2X0 U26121 ( .IN1(n23153), .IN2(n24737), .QN(n23198) );
  AO22X1 U26122 ( .IN1(n24759), .IN2(s11_ack_i), .IN3(n23198), .IN4(s12_ack_i), 
        .Q(n23163) );
  NOR2X0 U26123 ( .IN1(n23155), .IN2(n23154), .QN(n23250) );
  AND2X1 U26124 ( .IN1(n23250), .IN2(n23156), .Q(n28974) );
  INVX0 U26125 ( .INP(n28974), .ZN(n28949) );
  NOR2X0 U26126 ( .IN1(n23157), .IN2(n28949), .QN(n28112) );
  NOR2X0 U26127 ( .IN1(n23159), .IN2(n23158), .QN(n23218) );
  AND2X1 U26128 ( .IN1(n23160), .IN2(n23218), .Q(n29155) );
  INVX0 U26129 ( .INP(n29155), .ZN(n25348) );
  NOR2X0 U26130 ( .IN1(n23161), .IN2(n25348), .QN(n25064) );
  AO22X1 U26131 ( .IN1(n28112), .IN2(s0_ack_i), .IN3(n25064), .IN4(s10_ack_i), 
        .Q(n23162) );
  NOR2X0 U26132 ( .IN1(n23163), .IN2(n23162), .QN(n23169) );
  NOR2X0 U26133 ( .IN1(n23165), .IN2(n23164), .QN(n23234) );
  AND2X1 U26134 ( .IN1(n23166), .IN2(n23234), .Q(n29030) );
  INVX0 U26135 ( .INP(n29030), .ZN(n27438) );
  NOR2X0 U26136 ( .IN1(n23167), .IN2(n27438), .QN(n23197) );
  NAND2X0 U26137 ( .IN1(n23197), .IN2(s3_ack_i), .QN(n23168) );
  NAND2X0 U26138 ( .IN1(n23169), .IN2(n23168), .QN(n23170) );
  NOR4X0 U26139 ( .IN1(n23173), .IN2(n23172), .IN3(n23171), .IN4(n23170), .QN(
        n23175) );
  NAND2X0 U26140 ( .IN1(n23203), .IN2(n23261), .QN(n23174) );
  NAND4X0 U26141 ( .IN1(n23177), .IN2(n23176), .IN3(n23175), .IN4(n23174), 
        .QN(m0_ack_o) );
  INVX0 U26142 ( .INP(n23204), .ZN(n26281) );
  INVX0 U26143 ( .INP(n23198), .ZN(n24459) );
  OA22X1 U26144 ( .IN1(n26281), .IN2(n23400), .IN3(n24459), .IN4(n23407), .Q(
        n23189) );
  OA22X1 U26145 ( .IN1(n27498), .IN2(n23396), .IN3(n25373), .IN4(n23401), .Q(
        n23188) );
  AO22X1 U26146 ( .IN1(n23191), .IN2(s13_err_i), .IN3(n28112), .IN4(s0_err_i), 
        .Q(n23185) );
  INVX0 U26147 ( .INP(n25672), .ZN(n23195) );
  AO22X1 U26148 ( .IN1(n23195), .IN2(s8_err_i), .IN3(n26588), .IN4(s5_err_i), 
        .Q(n23184) );
  INVX0 U26149 ( .INP(n26892), .ZN(n23190) );
  AO22X1 U26150 ( .IN1(n23190), .IN2(s4_err_i), .IN3(n23196), .IN4(s7_err_i), 
        .Q(n23183) );
  AO22X1 U26151 ( .IN1(n23197), .IN2(s3_err_i), .IN3(n27807), .IN4(s1_err_i), 
        .Q(n23179) );
  AO22X1 U26152 ( .IN1(n24759), .IN2(s11_err_i), .IN3(n25064), .IN4(s10_err_i), 
        .Q(n23178) );
  NOR2X0 U26153 ( .IN1(n23179), .IN2(n23178), .QN(n23181) );
  NAND2X0 U26154 ( .IN1(n23847), .IN2(s14_err_i), .QN(n23180) );
  NAND2X0 U26155 ( .IN1(n23181), .IN2(n23180), .QN(n23182) );
  NOR4X0 U26156 ( .IN1(n23185), .IN2(n23184), .IN3(n23183), .IN4(n23182), .QN(
        n23187) );
  NAND3X0 U26157 ( .IN1(n23203), .IN2(s15_err_i), .IN3(n23445), .QN(n23186) );
  NAND4X0 U26158 ( .IN1(n23189), .IN2(n23188), .IN3(n23187), .IN4(n23186), 
        .QN(m0_err_o) );
  AO22X1 U26159 ( .IN1(n23190), .IN2(s4_rty_i), .IN3(n28112), .IN4(s0_rty_i), 
        .Q(n23194) );
  INVX0 U26160 ( .INP(n23191), .ZN(n24155) );
  OAI22X1 U26161 ( .IN1(n25373), .IN2(n23431), .IN3(n24155), .IN4(n23430), 
        .QN(n23193) );
  AO22X1 U26162 ( .IN1(n26588), .IN2(s5_rty_i), .IN3(n23847), .IN4(s14_rty_i), 
        .Q(n23192) );
  NOR3X0 U26163 ( .IN1(n23194), .IN2(n23193), .IN3(n23192), .QN(n23208) );
  AO22X1 U26164 ( .IN1(n23195), .IN2(s8_rty_i), .IN3(n25064), .IN4(s10_rty_i), 
        .Q(n23202) );
  AO22X1 U26165 ( .IN1(n23196), .IN2(s7_rty_i), .IN3(n24759), .IN4(s11_rty_i), 
        .Q(n23201) );
  INVX0 U26166 ( .INP(n23197), .ZN(n27196) );
  OAI22X1 U26167 ( .IN1(n27498), .IN2(n23435), .IN3(n27196), .IN4(n23427), 
        .QN(n23200) );
  AO22X1 U26168 ( .IN1(n27807), .IN2(s1_rty_i), .IN3(n23198), .IN4(s12_rty_i), 
        .Q(n23199) );
  NOR4X0 U26169 ( .IN1(n23202), .IN2(n23201), .IN3(n23200), .IN4(n23199), .QN(
        n23207) );
  NAND3X0 U26170 ( .IN1(n23203), .IN2(s15_rty_i), .IN3(n23445), .QN(n23206) );
  NAND2X0 U26171 ( .IN1(n23204), .IN2(s6_rty_i), .QN(n23205) );
  NAND4X0 U26172 ( .IN1(n23208), .IN2(n23207), .IN3(n23206), .IN4(n23205), 
        .QN(m0_rty_o) );
  NOR2X0 U26173 ( .IN1(n23210), .IN2(n23209), .QN(n29009) );
  NAND2X0 U26174 ( .IN1(n29268), .IN2(n29009), .QN(n27501) );
  AND2X1 U26175 ( .IN1(n23212), .IN2(n23211), .Q(n29200) );
  NAND2X0 U26176 ( .IN1(n29257), .IN2(n29200), .QN(n24153) );
  OA22X1 U26177 ( .IN1(n23214), .IN2(n27501), .IN3(n23213), .IN4(n24153), .Q(
        n23265) );
  AND2X1 U26178 ( .IN1(n23216), .IN2(n23215), .Q(n29093) );
  NAND2X0 U26179 ( .IN1(n29263), .IN2(n29093), .QN(n25979) );
  AND2X1 U26180 ( .IN1(n23218), .IN2(n23217), .Q(n29153) );
  NAND2X0 U26181 ( .IN1(n29260), .IN2(n29153), .QN(n25062) );
  OA22X1 U26182 ( .IN1(n23220), .IN2(n25979), .IN3(n23219), .IN4(n25062), .Q(
        n23264) );
  AND2X1 U26183 ( .IN1(n23222), .IN2(n23221), .Q(n29163) );
  INVX0 U26184 ( .INP(n29163), .ZN(n25044) );
  NOR2X0 U26185 ( .IN1(n23223), .IN2(n25044), .QN(n23278) );
  AND2X1 U26186 ( .IN1(n23225), .IN2(n23224), .Q(n29181) );
  INVX0 U26187 ( .INP(n29181), .ZN(n24747) );
  NOR2X0 U26188 ( .IN1(n23226), .IN2(n24747), .QN(n24454) );
  AO22X1 U26189 ( .IN1(s11_ack_i), .IN2(n23278), .IN3(s12_ack_i), .IN4(n24454), 
        .Q(n23260) );
  AND2X1 U26190 ( .IN1(n23228), .IN2(n23227), .Q(n29058) );
  INVX0 U26191 ( .INP(n29058), .ZN(n26878) );
  NOR2X0 U26192 ( .IN1(n23229), .IN2(n26878), .QN(n26583) );
  AND2X1 U26193 ( .IN1(n23231), .IN2(n23230), .Q(n29076) );
  INVX0 U26194 ( .INP(n29076), .ZN(n26560) );
  NOR2X0 U26195 ( .IN1(n23232), .IN2(n26560), .QN(n23280) );
  AO22X1 U26196 ( .IN1(s5_ack_i), .IN2(n26583), .IN3(s6_ack_i), .IN4(n23280), 
        .Q(n23259) );
  AND2X1 U26197 ( .IN1(n23234), .IN2(n23233), .Q(n29027) );
  INVX0 U26198 ( .INP(n29027), .ZN(n27480) );
  NOR2X0 U26199 ( .IN1(n23235), .IN2(n27480), .QN(n27197) );
  AND2X1 U26200 ( .IN1(n23237), .IN2(n23236), .Q(n28993) );
  INVX0 U26201 ( .INP(n28993), .ZN(n28103) );
  NOR2X0 U26202 ( .IN1(n23238), .IN2(n28103), .QN(n27804) );
  AO22X1 U26203 ( .IN1(s3_ack_i), .IN2(n27197), .IN3(s1_ack_i), .IN4(n27804), 
        .Q(n23258) );
  AND2X1 U26204 ( .IN1(n23240), .IN2(n23239), .Q(n29227) );
  INVX0 U26205 ( .INP(n29227), .ZN(n24139) );
  NOR2X0 U26206 ( .IN1(n23241), .IN2(n24139), .QN(n23846) );
  NAND2X0 U26207 ( .IN1(n23846), .IN2(s14_ack_i), .QN(n23256) );
  NOR2X0 U26208 ( .IN1(n23243), .IN2(n23242), .QN(n29040) );
  NAND2X0 U26209 ( .IN1(n29266), .IN2(n29040), .QN(n26895) );
  NOR2X0 U26210 ( .IN1(n23245), .IN2(n23244), .QN(n29117) );
  NAND2X0 U26211 ( .IN1(n29262), .IN2(n29117), .QN(n25678) );
  OA22X1 U26212 ( .IN1(n23247), .IN2(n26895), .IN3(n23246), .IN4(n25678), .Q(
        n23255) );
  NOR2X0 U26213 ( .IN1(n23249), .IN2(n23248), .QN(n29137) );
  NAND2X0 U26214 ( .IN1(n29261), .IN2(n29137), .QN(n25371) );
  AND2X1 U26215 ( .IN1(n23251), .IN2(n23250), .Q(n28968) );
  NAND2X0 U26216 ( .IN1(n29271), .IN2(n28968), .QN(n28116) );
  OA22X1 U26217 ( .IN1(n23253), .IN2(n25371), .IN3(n23252), .IN4(n28116), .Q(
        n23254) );
  NAND3X0 U26218 ( .IN1(n23256), .IN2(n23255), .IN3(n23254), .QN(n23257) );
  NOR4X0 U26219 ( .IN1(n23260), .IN2(n23259), .IN3(n23258), .IN4(n23257), .QN(
        n23263) );
  NAND2X0 U26220 ( .IN1(n23289), .IN2(n23261), .QN(n23262) );
  NAND4X0 U26221 ( .IN1(n23265), .IN2(n23264), .IN3(n23263), .IN4(n23262), 
        .QN(m1_ack_o) );
  AOI22X1 U26222 ( .IN1(n23846), .IN2(s14_err_i), .IN3(n27197), .IN4(s3_err_i), 
        .QN(n23277) );
  OA22X1 U26223 ( .IN1(n25979), .IN2(n23406), .IN3(n28116), .IN4(n23405), .Q(
        n23276) );
  NOR2X0 U26224 ( .IN1(n25371), .IN2(n23401), .QN(n23273) );
  AO22X1 U26225 ( .IN1(n26583), .IN2(s5_err_i), .IN3(n27804), .IN4(s1_err_i), 
        .Q(n23272) );
  INVX0 U26226 ( .INP(n24153), .ZN(n23279) );
  AO22X1 U26227 ( .IN1(n23278), .IN2(s11_err_i), .IN3(n23279), .IN4(s13_err_i), 
        .Q(n23271) );
  OA22X1 U26228 ( .IN1(n27501), .IN2(n23396), .IN3(n26895), .IN4(n23395), .Q(
        n23269) );
  OA22X1 U26229 ( .IN1(n25062), .IN2(n23408), .IN3(n25678), .IN4(n23394), .Q(
        n23268) );
  NAND2X0 U26230 ( .IN1(n23280), .IN2(s6_err_i), .QN(n23267) );
  NAND2X0 U26231 ( .IN1(n24454), .IN2(s12_err_i), .QN(n23266) );
  NAND4X0 U26232 ( .IN1(n23269), .IN2(n23268), .IN3(n23267), .IN4(n23266), 
        .QN(n23270) );
  NOR4X0 U26233 ( .IN1(n23273), .IN2(n23272), .IN3(n23271), .IN4(n23270), .QN(
        n23275) );
  NAND3X0 U26234 ( .IN1(n23289), .IN2(s15_err_i), .IN3(n23445), .QN(n23274) );
  NAND4X0 U26235 ( .IN1(n23277), .IN2(n23276), .IN3(n23275), .IN4(n23274), 
        .QN(m1_err_o) );
  AOI22X1 U26236 ( .IN1(n26583), .IN2(s5_rty_i), .IN3(n23846), .IN4(s14_rty_i), 
        .QN(n23293) );
  OA22X1 U26237 ( .IN1(n25979), .IN2(n23421), .IN3(n25371), .IN4(n23431), .Q(
        n23292) );
  INVX0 U26238 ( .INP(n23278), .ZN(n24757) );
  OAI22X1 U26239 ( .IN1(n24757), .IN2(n23426), .IN3(n27501), .IN4(n23435), 
        .QN(n23288) );
  AO22X1 U26240 ( .IN1(n24454), .IN2(s12_rty_i), .IN3(n23279), .IN4(s13_rty_i), 
        .Q(n23287) );
  INVX0 U26241 ( .INP(n23280), .ZN(n26280) );
  OAI22X1 U26242 ( .IN1(n26280), .IN2(n23429), .IN3(n25678), .IN4(n23428), 
        .QN(n23286) );
  OA22X1 U26243 ( .IN1(n28116), .IN2(n23432), .IN3(n26895), .IN4(n23436), .Q(
        n23284) );
  NAND2X0 U26244 ( .IN1(n27804), .IN2(s1_rty_i), .QN(n23283) );
  NAND2X0 U26245 ( .IN1(n27197), .IN2(s3_rty_i), .QN(n23282) );
  OR2X1 U26246 ( .IN1(n25062), .IN2(n23422), .Q(n23281) );
  NAND4X0 U26247 ( .IN1(n23284), .IN2(n23283), .IN3(n23282), .IN4(n23281), 
        .QN(n23285) );
  NOR4X0 U26248 ( .IN1(n23288), .IN2(n23287), .IN3(n23286), .IN4(n23285), .QN(
        n23291) );
  NAND3X0 U26249 ( .IN1(n23289), .IN2(s15_rty_i), .IN3(n23445), .QN(n23290) );
  NAND4X0 U26250 ( .IN1(n23293), .IN2(n23292), .IN3(n23291), .IN4(n23290), 
        .QN(m1_rty_o) );
  OA22X1 U26251 ( .IN1(n26589), .IN2(n23404), .IN3(n27500), .IN4(n23396), .Q(
        n23305) );
  OA22X1 U26252 ( .IN1(n23850), .IN2(n23398), .IN3(n25369), .IN4(n23401), .Q(
        n23304) );
  OA22X1 U26253 ( .IN1(n26279), .IN2(n23400), .IN3(n24152), .IN4(n23402), .Q(
        n23301) );
  OA22X1 U26254 ( .IN1(n25671), .IN2(n23394), .IN3(n24762), .IN4(n23397), .Q(
        n23300) );
  OA22X1 U26255 ( .IN1(n25977), .IN2(n23406), .IN3(n27198), .IN4(n23399), .Q(
        n23299) );
  NOR2X0 U26256 ( .IN1(n23408), .IN2(n25065), .QN(n23297) );
  OA22X1 U26257 ( .IN1(n26893), .IN2(n23395), .IN3(n24455), .IN4(n23407), .Q(
        n23295) );
  INVX0 U26258 ( .INP(s1_err_i), .ZN(n23403) );
  OA22X1 U26259 ( .IN1(n27802), .IN2(n23403), .IN3(n28110), .IN4(n23405), .Q(
        n23294) );
  NAND2X0 U26260 ( .IN1(n23295), .IN2(n23294), .QN(n23296) );
  NOR2X0 U26261 ( .IN1(n23297), .IN2(n23296), .QN(n23298) );
  AND4X1 U26262 ( .IN1(n23301), .IN2(n23300), .IN3(n23299), .IN4(n23298), .Q(
        n23303) );
  NAND3X0 U26263 ( .IN1(n23314), .IN2(s15_err_i), .IN3(n23445), .QN(n23302) );
  NAND4X0 U26264 ( .IN1(n23305), .IN2(n23304), .IN3(n23303), .IN4(n23302), 
        .QN(m3_err_o) );
  OA22X1 U26265 ( .IN1(n25369), .IN2(n23431), .IN3(n28110), .IN4(n23432), .Q(
        n23318) );
  OA22X1 U26266 ( .IN1(n24762), .IN2(n23426), .IN3(n26589), .IN4(n23423), .Q(
        n23317) );
  OA22X1 U26267 ( .IN1(n24152), .IN2(n23430), .IN3(n24455), .IN4(n23425), .Q(
        n23313) );
  OA22X1 U26268 ( .IN1(n26279), .IN2(n23429), .IN3(n27198), .IN4(n23427), .Q(
        n23312) );
  OA22X1 U26269 ( .IN1(n23850), .IN2(n23433), .IN3(n25671), .IN4(n23428), .Q(
        n23311) );
  NOR2X0 U26270 ( .IN1(n23422), .IN2(n25065), .QN(n23309) );
  OA22X1 U26271 ( .IN1(n26893), .IN2(n23436), .IN3(n25977), .IN4(n23421), .Q(
        n23307) );
  OA22X1 U26272 ( .IN1(n27802), .IN2(n23424), .IN3(n27500), .IN4(n23435), .Q(
        n23306) );
  NAND2X0 U26273 ( .IN1(n23307), .IN2(n23306), .QN(n23308) );
  NOR2X0 U26274 ( .IN1(n23309), .IN2(n23308), .QN(n23310) );
  AND4X1 U26275 ( .IN1(n23313), .IN2(n23312), .IN3(n23311), .IN4(n23310), .Q(
        n23316) );
  NAND3X0 U26276 ( .IN1(n23314), .IN2(s15_rty_i), .IN3(n23445), .QN(n23315) );
  NAND4X0 U26277 ( .IN1(n23318), .IN2(n23317), .IN3(n23316), .IN4(n23315), 
        .QN(m3_rty_o) );
  OA22X1 U26278 ( .IN1(n25067), .IN2(n23408), .IN3(n26891), .IN4(n23395), .Q(
        n23330) );
  OA22X1 U26279 ( .IN1(n23848), .IN2(n23398), .IN3(n27805), .IN4(n23403), .Q(
        n23329) );
  OA22X1 U26280 ( .IN1(n24154), .IN2(n23402), .IN3(n24452), .IN4(n23407), .Q(
        n23326) );
  OA22X1 U26281 ( .IN1(n25975), .IN2(n23406), .IN3(n27504), .IN4(n23396), .Q(
        n23325) );
  OA22X1 U26282 ( .IN1(n25367), .IN2(n23401), .IN3(n25673), .IN4(n23394), .Q(
        n23324) );
  NOR2X0 U26283 ( .IN1(n23397), .IN2(n24760), .QN(n23322) );
  OA22X1 U26284 ( .IN1(n26584), .IN2(n23404), .IN3(n26283), .IN4(n23400), .Q(
        n23320) );
  OA22X1 U26285 ( .IN1(n28115), .IN2(n23405), .IN3(n27195), .IN4(n23399), .Q(
        n23319) );
  NAND2X0 U26286 ( .IN1(n23320), .IN2(n23319), .QN(n23321) );
  NOR2X0 U26287 ( .IN1(n23322), .IN2(n23321), .QN(n23323) );
  AND4X1 U26288 ( .IN1(n23326), .IN2(n23325), .IN3(n23324), .IN4(n23323), .Q(
        n23328) );
  NAND3X0 U26289 ( .IN1(n23339), .IN2(s15_err_i), .IN3(n23445), .QN(n23327) );
  NAND4X0 U26290 ( .IN1(n23330), .IN2(n23329), .IN3(n23328), .IN4(n23327), 
        .QN(m4_err_o) );
  OA22X1 U26291 ( .IN1(n24760), .IN2(n23426), .IN3(n24452), .IN4(n23425), .Q(
        n23343) );
  OA22X1 U26292 ( .IN1(n25367), .IN2(n23431), .IN3(n26891), .IN4(n23436), .Q(
        n23342) );
  OA22X1 U26293 ( .IN1(n25975), .IN2(n23421), .IN3(n23848), .IN4(n23433), .Q(
        n23338) );
  OA22X1 U26294 ( .IN1(n28115), .IN2(n23432), .IN3(n26283), .IN4(n23429), .Q(
        n23337) );
  OA22X1 U26295 ( .IN1(n26584), .IN2(n23423), .IN3(n27504), .IN4(n23435), .Q(
        n23336) );
  NOR2X0 U26296 ( .IN1(n23430), .IN2(n24154), .QN(n23334) );
  OA22X1 U26297 ( .IN1(n25067), .IN2(n23422), .IN3(n27805), .IN4(n23424), .Q(
        n23332) );
  OA22X1 U26298 ( .IN1(n25673), .IN2(n23428), .IN3(n27195), .IN4(n23427), .Q(
        n23331) );
  NAND2X0 U26299 ( .IN1(n23332), .IN2(n23331), .QN(n23333) );
  NOR2X0 U26300 ( .IN1(n23334), .IN2(n23333), .QN(n23335) );
  AND4X1 U26301 ( .IN1(n23338), .IN2(n23337), .IN3(n23336), .IN4(n23335), .Q(
        n23341) );
  NAND3X0 U26302 ( .IN1(n23339), .IN2(s15_rty_i), .IN3(n23445), .QN(n23340) );
  NAND4X0 U26303 ( .IN1(n23343), .IN2(n23342), .IN3(n23341), .IN4(n23340), 
        .QN(m4_rty_o) );
  OA22X1 U26304 ( .IN1(n27803), .IN2(n23403), .IN3(n26889), .IN4(n23395), .Q(
        n23355) );
  OA22X1 U26305 ( .IN1(n25069), .IN2(n23408), .IN3(n27200), .IN4(n23399), .Q(
        n23354) );
  OA22X1 U26306 ( .IN1(n24148), .IN2(n23402), .IN3(n25677), .IN4(n23394), .Q(
        n23351) );
  OA22X1 U26307 ( .IN1(n28108), .IN2(n23405), .IN3(n26285), .IN4(n23400), .Q(
        n23350) );
  OA22X1 U26308 ( .IN1(n27502), .IN2(n23396), .IN3(n26586), .IN4(n23404), .Q(
        n23349) );
  NOR2X0 U26309 ( .IN1(n23407), .IN2(n24457), .QN(n23347) );
  OA22X1 U26310 ( .IN1(n24764), .IN2(n23397), .IN3(n25976), .IN4(n23406), .Q(
        n23345) );
  OA22X1 U26311 ( .IN1(n25370), .IN2(n23401), .IN3(n23843), .IN4(n23398), .Q(
        n23344) );
  NAND2X0 U26312 ( .IN1(n23345), .IN2(n23344), .QN(n23346) );
  NOR2X0 U26313 ( .IN1(n23347), .IN2(n23346), .QN(n23348) );
  AND4X1 U26314 ( .IN1(n23351), .IN2(n23350), .IN3(n23349), .IN4(n23348), .Q(
        n23353) );
  NAND3X0 U26315 ( .IN1(n23364), .IN2(s15_err_i), .IN3(n23445), .QN(n23352) );
  NAND4X0 U26316 ( .IN1(n23355), .IN2(n23354), .IN3(n23353), .IN4(n23352), 
        .QN(m5_err_o) );
  OA22X1 U26317 ( .IN1(n27502), .IN2(n23435), .IN3(n27200), .IN4(n23427), .Q(
        n23368) );
  OA22X1 U26318 ( .IN1(n28108), .IN2(n23432), .IN3(n23843), .IN4(n23433), .Q(
        n23367) );
  OA22X1 U26319 ( .IN1(n24148), .IN2(n23430), .IN3(n26889), .IN4(n23436), .Q(
        n23363) );
  OA22X1 U26320 ( .IN1(n25370), .IN2(n23431), .IN3(n26285), .IN4(n23429), .Q(
        n23362) );
  OA22X1 U26321 ( .IN1(n25069), .IN2(n23422), .IN3(n26586), .IN4(n23423), .Q(
        n23361) );
  NOR2X0 U26322 ( .IN1(n23426), .IN2(n24764), .QN(n23359) );
  OA22X1 U26323 ( .IN1(n24457), .IN2(n23425), .IN3(n25976), .IN4(n23421), .Q(
        n23357) );
  OA22X1 U26324 ( .IN1(n27803), .IN2(n23424), .IN3(n25677), .IN4(n23428), .Q(
        n23356) );
  NAND2X0 U26325 ( .IN1(n23357), .IN2(n23356), .QN(n23358) );
  NOR2X0 U26326 ( .IN1(n23359), .IN2(n23358), .QN(n23360) );
  AND4X1 U26327 ( .IN1(n23363), .IN2(n23362), .IN3(n23361), .IN4(n23360), .Q(
        n23366) );
  NAND3X0 U26328 ( .IN1(n23364), .IN2(s15_rty_i), .IN3(n23445), .QN(n23365) );
  NAND4X0 U26329 ( .IN1(n23368), .IN2(n23367), .IN3(n23366), .IN4(n23365), 
        .QN(m5_rty_o) );
  OA22X1 U26330 ( .IN1(n23851), .IN2(n23398), .IN3(n24758), .IN4(n23397), .Q(
        n23380) );
  OA22X1 U26331 ( .IN1(n25980), .IN2(n23406), .IN3(n27810), .IN4(n23403), .Q(
        n23379) );
  OA22X1 U26332 ( .IN1(n26591), .IN2(n23404), .IN3(n24453), .IN4(n23407), .Q(
        n23376) );
  OA22X1 U26333 ( .IN1(n26896), .IN2(n23395), .IN3(n24150), .IN4(n23402), .Q(
        n23375) );
  OA22X1 U26334 ( .IN1(n26284), .IN2(n23400), .IN3(n25068), .IN4(n23408), .Q(
        n23374) );
  NOR2X0 U26335 ( .IN1(n23396), .IN2(n27499), .QN(n23372) );
  OA22X1 U26336 ( .IN1(n27193), .IN2(n23399), .IN3(n28114), .IN4(n23405), .Q(
        n23370) );
  OA22X1 U26337 ( .IN1(n25675), .IN2(n23394), .IN3(n25374), .IN4(n23401), .Q(
        n23369) );
  NAND2X0 U26338 ( .IN1(n23370), .IN2(n23369), .QN(n23371) );
  NOR2X0 U26339 ( .IN1(n23372), .IN2(n23371), .QN(n23373) );
  AND4X1 U26340 ( .IN1(n23376), .IN2(n23375), .IN3(n23374), .IN4(n23373), .Q(
        n23378) );
  NAND3X0 U26341 ( .IN1(n23389), .IN2(s15_err_i), .IN3(n23445), .QN(n23377) );
  NAND4X0 U26342 ( .IN1(n23380), .IN2(n23379), .IN3(n23378), .IN4(n23377), 
        .QN(m6_err_o) );
  OA22X1 U26343 ( .IN1(n24758), .IN2(n23426), .IN3(n25068), .IN4(n23422), .Q(
        n23393) );
  OA22X1 U26344 ( .IN1(n26591), .IN2(n23423), .IN3(n28114), .IN4(n23432), .Q(
        n23392) );
  OA22X1 U26345 ( .IN1(n27810), .IN2(n23424), .IN3(n25675), .IN4(n23428), .Q(
        n23388) );
  OA22X1 U26346 ( .IN1(n23851), .IN2(n23433), .IN3(n24453), .IN4(n23425), .Q(
        n23387) );
  OA22X1 U26347 ( .IN1(n27193), .IN2(n23427), .IN3(n26284), .IN4(n23429), .Q(
        n23386) );
  NOR2X0 U26348 ( .IN1(n23435), .IN2(n27499), .QN(n23384) );
  OA22X1 U26349 ( .IN1(n26896), .IN2(n23436), .IN3(n24150), .IN4(n23430), .Q(
        n23382) );
  OA22X1 U26350 ( .IN1(n25980), .IN2(n23421), .IN3(n25374), .IN4(n23431), .Q(
        n23381) );
  NAND2X0 U26351 ( .IN1(n23382), .IN2(n23381), .QN(n23383) );
  NOR2X0 U26352 ( .IN1(n23384), .IN2(n23383), .QN(n23385) );
  AND4X1 U26353 ( .IN1(n23388), .IN2(n23387), .IN3(n23386), .IN4(n23385), .Q(
        n23391) );
  NAND3X0 U26354 ( .IN1(n23389), .IN2(s15_rty_i), .IN3(n23445), .QN(n23390) );
  NAND4X0 U26355 ( .IN1(n23393), .IN2(n23392), .IN3(n23391), .IN4(n23390), 
        .QN(m6_rty_o) );
  OA22X1 U26356 ( .IN1(n26890), .IN2(n23395), .IN3(n25674), .IN4(n23394), .Q(
        n23420) );
  OA22X1 U26357 ( .IN1(n24763), .IN2(n23397), .IN3(n27505), .IN4(n23396), .Q(
        n23419) );
  INVX0 U26358 ( .INP(n23845), .ZN(n23434) );
  OA22X1 U26359 ( .IN1(n27201), .IN2(n23399), .IN3(n23434), .IN4(n23398), .Q(
        n23416) );
  OA22X1 U26360 ( .IN1(n25368), .IN2(n23401), .IN3(n26286), .IN4(n23400), .Q(
        n23415) );
  OA22X1 U26361 ( .IN1(n27809), .IN2(n23403), .IN3(n24149), .IN4(n23402), .Q(
        n23414) );
  NOR2X0 U26362 ( .IN1(n23404), .IN2(n26587), .QN(n23412) );
  OA22X1 U26363 ( .IN1(n25981), .IN2(n23406), .IN3(n28111), .IN4(n23405), .Q(
        n23410) );
  OA22X1 U26364 ( .IN1(n25070), .IN2(n23408), .IN3(n24460), .IN4(n23407), .Q(
        n23409) );
  NAND2X0 U26365 ( .IN1(n23410), .IN2(n23409), .QN(n23411) );
  NOR2X0 U26366 ( .IN1(n23412), .IN2(n23411), .QN(n23413) );
  AND4X1 U26367 ( .IN1(n23416), .IN2(n23415), .IN3(n23414), .IN4(n23413), .Q(
        n23418) );
  NAND3X0 U26368 ( .IN1(n23446), .IN2(s15_err_i), .IN3(n23445), .QN(n23417) );
  NAND4X0 U26369 ( .IN1(n23420), .IN2(n23419), .IN3(n23418), .IN4(n23417), 
        .QN(m7_err_o) );
  OA22X1 U26370 ( .IN1(n25070), .IN2(n23422), .IN3(n25981), .IN4(n23421), .Q(
        n23450) );
  OA22X1 U26371 ( .IN1(n27809), .IN2(n23424), .IN3(n26587), .IN4(n23423), .Q(
        n23449) );
  OA22X1 U26372 ( .IN1(n24763), .IN2(n23426), .IN3(n24460), .IN4(n23425), .Q(
        n23444) );
  OA22X1 U26373 ( .IN1(n25674), .IN2(n23428), .IN3(n27201), .IN4(n23427), .Q(
        n23443) );
  OA22X1 U26374 ( .IN1(n24149), .IN2(n23430), .IN3(n26286), .IN4(n23429), .Q(
        n23442) );
  NOR2X0 U26375 ( .IN1(n23431), .IN2(n25368), .QN(n23440) );
  OA22X1 U26376 ( .IN1(n23434), .IN2(n23433), .IN3(n28111), .IN4(n23432), .Q(
        n23438) );
  OA22X1 U26377 ( .IN1(n26890), .IN2(n23436), .IN3(n27505), .IN4(n23435), .Q(
        n23437) );
  NAND2X0 U26378 ( .IN1(n23438), .IN2(n23437), .QN(n23439) );
  NOR2X0 U26379 ( .IN1(n23440), .IN2(n23439), .QN(n23441) );
  AND4X1 U26380 ( .IN1(n23444), .IN2(n23443), .IN3(n23442), .IN4(n23441), .Q(
        n23448) );
  NAND3X0 U26381 ( .IN1(n23446), .IN2(s15_rty_i), .IN3(n23445), .QN(n23447) );
  NAND4X0 U26382 ( .IN1(n23450), .IN2(n23449), .IN3(n23448), .IN4(n23447), 
        .QN(m7_rty_o) );
  NOR2X0 U26383 ( .IN1(n18178), .IN2(n23451), .QN(s15_cyc_o) );
  NOR2X0 U26384 ( .IN1(s15_addr_o[2]), .IN2(s15_addr_o[3]), .QN(n23459) );
  INVX0 U26385 ( .INP(s15_addr_o[5]), .ZN(n23458) );
  NOR2X0 U26386 ( .IN1(n23458), .IN2(s15_addr_o[4]), .QN(n23461) );
  NAND2X0 U26387 ( .IN1(n23459), .IN2(n23461), .QN(n31938) );
  INVX0 U26388 ( .INP(s15_addr_o[4]), .ZN(n23457) );
  NOR2X0 U26389 ( .IN1(n23457), .IN2(s15_addr_o[5]), .QN(n23462) );
  NAND2X0 U26390 ( .IN1(n23459), .IN2(n23462), .QN(n30624) );
  OA22X1 U26391 ( .IN1(n13916), .IN2(n31938), .IN3(n13888), .IN4(n30624), .Q(
        n23456) );
  INVX0 U26392 ( .INP(s15_addr_o[2]), .ZN(n23452) );
  AND2X1 U26393 ( .IN1(s15_addr_o[3]), .IN2(n23452), .Q(n23460) );
  NAND2X0 U26394 ( .IN1(n23460), .IN2(n23461), .QN(n32456) );
  NOR2X0 U26395 ( .IN1(n23452), .IN2(s15_addr_o[3]), .QN(n23465) );
  NAND2X0 U26396 ( .IN1(n23465), .IN2(n23462), .QN(n30975) );
  OA22X1 U26397 ( .IN1(n13920), .IN2(n32456), .IN3(n13890), .IN4(n30975), .Q(
        n23455) );
  NAND4X0 U26398 ( .IN1(s15_addr_o[5]), .IN2(s15_addr_o[4]), .IN3(
        s15_addr_o[2]), .IN4(s15_addr_o[3]), .QN(n33762) );
  NOR2X0 U26399 ( .IN1(s15_addr_o[5]), .IN2(s15_addr_o[4]), .QN(n23464) );
  NAND2X0 U26400 ( .IN1(n23464), .IN2(n23459), .QN(n29387) );
  OA22X1 U26401 ( .IN1(n13914), .IN2(n33762), .IN3(n13896), .IN4(n29387), .Q(
        n23454) );
  AND2X1 U26402 ( .IN1(s15_addr_o[2]), .IN2(s15_addr_o[3]), .Q(n23463) );
  NAND2X0 U26403 ( .IN1(n23464), .IN2(n23463), .QN(n30329) );
  NAND2X0 U26404 ( .IN1(n23460), .IN2(n23462), .QN(n31332) );
  OA22X1 U26405 ( .IN1(n13902), .IN2(n30329), .IN3(n13892), .IN4(n31332), .Q(
        n23453) );
  NAND4X0 U26406 ( .IN1(n23456), .IN2(n23455), .IN3(n23454), .IN4(n23453), 
        .QN(n23472) );
  NAND2X0 U26407 ( .IN1(n23463), .IN2(n23461), .QN(n32714) );
  NOR2X0 U26408 ( .IN1(n23458), .IN2(n23457), .QN(n23466) );
  NAND2X0 U26409 ( .IN1(n23466), .IN2(n23459), .QN(n32944) );
  OA22X1 U26410 ( .IN1(n13922), .IN2(n32714), .IN3(n13908), .IN4(n32944), .Q(
        n23470) );
  NAND2X0 U26411 ( .IN1(n23460), .IN2(n23464), .QN(n30008) );
  NAND2X0 U26412 ( .IN1(n23466), .IN2(n23460), .QN(n33536) );
  OA22X1 U26413 ( .IN1(n13900), .IN2(n30008), .IN3(n13912), .IN4(n33536), .Q(
        n23469) );
  NAND2X0 U26414 ( .IN1(n23461), .IN2(n23465), .QN(n32138) );
  NAND2X0 U26415 ( .IN1(n23463), .IN2(n23462), .QN(n31627) );
  OA22X1 U26416 ( .IN1(n13918), .IN2(n32138), .IN3(n13894), .IN4(n31627), .Q(
        n23468) );
  NAND2X0 U26417 ( .IN1(n23464), .IN2(n23465), .QN(n29729) );
  NAND2X0 U26418 ( .IN1(n23466), .IN2(n23465), .QN(n33238) );
  OA22X1 U26419 ( .IN1(n13898), .IN2(n29729), .IN3(n13910), .IN4(n33238), .Q(
        n23467) );
  NAND4X0 U26420 ( .IN1(n23470), .IN2(n23469), .IN3(n23468), .IN4(n23467), 
        .QN(n23471) );
  OA21X1 U26421 ( .IN1(n23472), .IN2(n23471), .IN3(n23501), .Q(\rf/N115 ) );
  OA22X1 U26422 ( .IN1(n13862), .IN2(n30975), .IN3(n13874), .IN4(n33238), .Q(
        n23476) );
  OA22X1 U26423 ( .IN1(n13878), .IN2(n32138), .IN3(n13867), .IN4(n30008), .Q(
        n23475) );
  OA22X1 U26424 ( .IN1(n13873), .IN2(n32944), .IN3(n13865), .IN4(n29387), .Q(
        n23474) );
  OA22X1 U26425 ( .IN1(n13868), .IN2(n30329), .IN3(n13880), .IN4(n32714), .Q(
        n23473) );
  NAND4X0 U26426 ( .IN1(n23476), .IN2(n23475), .IN3(n23474), .IN4(n23473), 
        .QN(n23482) );
  OA22X1 U26427 ( .IN1(n13864), .IN2(n31627), .IN3(n13879), .IN4(n32456), .Q(
        n23480) );
  OA22X1 U26428 ( .IN1(n13876), .IN2(n33762), .IN3(n13875), .IN4(n33536), .Q(
        n23479) );
  OA22X1 U26429 ( .IN1(n13861), .IN2(n30624), .IN3(n13866), .IN4(n29729), .Q(
        n23478) );
  OA22X1 U26430 ( .IN1(n13877), .IN2(n31938), .IN3(n13863), .IN4(n31332), .Q(
        n23477) );
  NAND4X0 U26431 ( .IN1(n23480), .IN2(n23479), .IN3(n23478), .IN4(n23477), 
        .QN(n23481) );
  OA21X1 U26432 ( .IN1(n23482), .IN2(n23481), .IN3(n23501), .Q(\rf/N116 ) );
  OA22X1 U26433 ( .IN1(n13852), .IN2(n32138), .IN3(n13850), .IN4(n33762), .Q(
        n23486) );
  OA22X1 U26434 ( .IN1(n13848), .IN2(n33238), .IN3(n13841), .IN4(n30008), .Q(
        n23485) );
  OA22X1 U26435 ( .IN1(n13851), .IN2(n31938), .IN3(n13838), .IN4(n31627), .Q(
        n23484) );
  OA22X1 U26436 ( .IN1(n13854), .IN2(n32714), .IN3(n13837), .IN4(n31332), .Q(
        n23483) );
  NAND4X0 U26437 ( .IN1(n23486), .IN2(n23485), .IN3(n23484), .IN4(n23483), 
        .QN(n23492) );
  OA22X1 U26438 ( .IN1(n13849), .IN2(n33536), .IN3(n13836), .IN4(n30975), .Q(
        n23490) );
  OA22X1 U26439 ( .IN1(n13840), .IN2(n29729), .IN3(n13839), .IN4(n29387), .Q(
        n23489) );
  OA22X1 U26440 ( .IN1(n13842), .IN2(n30329), .IN3(n13847), .IN4(n32944), .Q(
        n23488) );
  OA22X1 U26441 ( .IN1(n13835), .IN2(n30624), .IN3(n13853), .IN4(n32456), .Q(
        n23487) );
  NAND4X0 U26442 ( .IN1(n23490), .IN2(n23489), .IN3(n23488), .IN4(n23487), 
        .QN(n23491) );
  OA21X1 U26443 ( .IN1(n23492), .IN2(n23491), .IN3(n23501), .Q(\rf/N117 ) );
  OA22X1 U26444 ( .IN1(n13814), .IN2(n29729), .IN3(n13811), .IN4(n31332), .Q(
        n23496) );
  OA22X1 U26445 ( .IN1(n13827), .IN2(n32456), .IN3(n13815), .IN4(n30008), .Q(
        n23495) );
  OA22X1 U26446 ( .IN1(n13816), .IN2(n30329), .IN3(n13826), .IN4(n32138), .Q(
        n23494) );
  OA22X1 U26447 ( .IN1(n13809), .IN2(n30624), .IN3(n13825), .IN4(n31938), .Q(
        n23493) );
  NAND4X0 U26448 ( .IN1(n23496), .IN2(n23495), .IN3(n23494), .IN4(n23493), 
        .QN(n23503) );
  OA22X1 U26449 ( .IN1(n13822), .IN2(n33238), .IN3(n13824), .IN4(n33762), .Q(
        n23500) );
  OA22X1 U26450 ( .IN1(n13823), .IN2(n33536), .IN3(n13828), .IN4(n32714), .Q(
        n23499) );
  OA22X1 U26451 ( .IN1(n13810), .IN2(n30975), .IN3(n13813), .IN4(n29387), .Q(
        n23498) );
  OA22X1 U26452 ( .IN1(n13821), .IN2(n32944), .IN3(n13812), .IN4(n31627), .Q(
        n23497) );
  NAND4X0 U26453 ( .IN1(n23500), .IN2(n23499), .IN3(n23498), .IN4(n23497), 
        .QN(n23502) );
  OA21X1 U26454 ( .IN1(n23503), .IN2(n23502), .IN3(n23501), .Q(\rf/N118 ) );
  OA22X1 U26455 ( .IN1(n13795), .IN2(n32944), .IN3(n13788), .IN4(n29729), .Q(
        n23507) );
  OA22X1 U26456 ( .IN1(n13801), .IN2(n32456), .IN3(n13783), .IN4(n30624), .Q(
        n23506) );
  OA22X1 U26457 ( .IN1(n13785), .IN2(n31332), .IN3(n13784), .IN4(n30975), .Q(
        n23505) );
  OA22X1 U26458 ( .IN1(n13786), .IN2(n31627), .IN3(n13789), .IN4(n30008), .Q(
        n23504) );
  NAND4X0 U26459 ( .IN1(n23507), .IN2(n23506), .IN3(n23505), .IN4(n23504), 
        .QN(n23513) );
  OA22X1 U26460 ( .IN1(n13798), .IN2(n33762), .IN3(n13796), .IN4(n33238), .Q(
        n23511) );
  OA22X1 U26461 ( .IN1(n13802), .IN2(n32714), .IN3(n13800), .IN4(n32138), .Q(
        n23510) );
  OA22X1 U26462 ( .IN1(n13787), .IN2(n29387), .IN3(n13790), .IN4(n30329), .Q(
        n23509) );
  OA22X1 U26463 ( .IN1(n13797), .IN2(n33536), .IN3(n13799), .IN4(n31938), .Q(
        n23508) );
  NAND4X0 U26464 ( .IN1(n23511), .IN2(n23510), .IN3(n23509), .IN4(n23508), 
        .QN(n23512) );
  OA21X1 U26465 ( .IN1(n23513), .IN2(n23512), .IN3(n23622), .Q(\rf/N119 ) );
  OA22X1 U26466 ( .IN1(n13771), .IN2(n33536), .IN3(n13764), .IN4(n30329), .Q(
        n23517) );
  OA22X1 U26467 ( .IN1(n13773), .IN2(n31938), .IN3(n13757), .IN4(n30624), .Q(
        n23516) );
  OA22X1 U26468 ( .IN1(n13770), .IN2(n33238), .IN3(n13774), .IN4(n32138), .Q(
        n23515) );
  OA22X1 U26469 ( .IN1(n13775), .IN2(n32456), .IN3(n13772), .IN4(n33762), .Q(
        n23514) );
  NAND4X0 U26470 ( .IN1(n23517), .IN2(n23516), .IN3(n23515), .IN4(n23514), 
        .QN(n23523) );
  OA22X1 U26471 ( .IN1(n13760), .IN2(n31627), .IN3(n13761), .IN4(n29387), .Q(
        n23521) );
  OA22X1 U26472 ( .IN1(n13758), .IN2(n30975), .IN3(n13769), .IN4(n32944), .Q(
        n23520) );
  OA22X1 U26473 ( .IN1(n13759), .IN2(n31332), .IN3(n13762), .IN4(n29729), .Q(
        n23519) );
  OA22X1 U26474 ( .IN1(n13763), .IN2(n30008), .IN3(n13776), .IN4(n32714), .Q(
        n23518) );
  NAND4X0 U26475 ( .IN1(n23521), .IN2(n23520), .IN3(n23519), .IN4(n23518), 
        .QN(n23522) );
  OA21X1 U26476 ( .IN1(n23523), .IN2(n23522), .IN3(n23622), .Q(\rf/N120 ) );
  OA22X1 U26477 ( .IN1(n13732), .IN2(n30975), .IN3(n13737), .IN4(n30008), .Q(
        n23527) );
  OA22X1 U26478 ( .IN1(n13731), .IN2(n30624), .IN3(n13749), .IN4(n32456), .Q(
        n23526) );
  OA22X1 U26479 ( .IN1(n13748), .IN2(n32138), .IN3(n13746), .IN4(n33762), .Q(
        n23525) );
  OA22X1 U26480 ( .IN1(n13743), .IN2(n32944), .IN3(n13745), .IN4(n33536), .Q(
        n23524) );
  NAND4X0 U26481 ( .IN1(n23527), .IN2(n23526), .IN3(n23525), .IN4(n23524), 
        .QN(n23533) );
  OA22X1 U26482 ( .IN1(n13738), .IN2(n30329), .IN3(n13744), .IN4(n33238), .Q(
        n23531) );
  OA22X1 U26483 ( .IN1(n13735), .IN2(n29387), .IN3(n13747), .IN4(n31938), .Q(
        n23530) );
  OA22X1 U26484 ( .IN1(n13750), .IN2(n32714), .IN3(n13733), .IN4(n31332), .Q(
        n23529) );
  OA22X1 U26485 ( .IN1(n13734), .IN2(n31627), .IN3(n13736), .IN4(n29729), .Q(
        n23528) );
  NAND4X0 U26486 ( .IN1(n23531), .IN2(n23530), .IN3(n23529), .IN4(n23528), 
        .QN(n23532) );
  OA21X1 U26487 ( .IN1(n23533), .IN2(n23532), .IN3(n23622), .Q(\rf/N121 ) );
  OA22X1 U26488 ( .IN1(n13721), .IN2(n31938), .IN3(n13707), .IN4(n31332), .Q(
        n23537) );
  OA22X1 U26489 ( .IN1(n13708), .IN2(n31627), .IN3(n13720), .IN4(n33762), .Q(
        n23536) );
  OA22X1 U26490 ( .IN1(n13712), .IN2(n30329), .IN3(n13722), .IN4(n32138), .Q(
        n23535) );
  OA22X1 U26491 ( .IN1(n13706), .IN2(n30975), .IN3(n13718), .IN4(n33238), .Q(
        n23534) );
  NAND4X0 U26492 ( .IN1(n23537), .IN2(n23536), .IN3(n23535), .IN4(n23534), 
        .QN(n23543) );
  OA22X1 U26493 ( .IN1(n13723), .IN2(n32456), .IN3(n13719), .IN4(n33536), .Q(
        n23541) );
  OA22X1 U26494 ( .IN1(n13724), .IN2(n32714), .IN3(n13711), .IN4(n30008), .Q(
        n23540) );
  OA22X1 U26495 ( .IN1(n13717), .IN2(n32944), .IN3(n13705), .IN4(n30624), .Q(
        n23539) );
  OA22X1 U26496 ( .IN1(n13709), .IN2(n29387), .IN3(n13710), .IN4(n29729), .Q(
        n23538) );
  NAND4X0 U26497 ( .IN1(n23541), .IN2(n23540), .IN3(n23539), .IN4(n23538), 
        .QN(n23542) );
  OA21X1 U26498 ( .IN1(n23543), .IN2(n23542), .IN3(n23622), .Q(\rf/N122 ) );
  OA22X1 U26499 ( .IN1(n13683), .IN2(n29387), .IN3(n13686), .IN4(n30329), .Q(
        n23547) );
  OA22X1 U26500 ( .IN1(n13697), .IN2(n32456), .IN3(n13695), .IN4(n31938), .Q(
        n23546) );
  OA22X1 U26501 ( .IN1(n13680), .IN2(n30975), .IN3(n13679), .IN4(n30624), .Q(
        n23545) );
  OA22X1 U26502 ( .IN1(n13694), .IN2(n33762), .IN3(n13682), .IN4(n31627), .Q(
        n23544) );
  NAND4X0 U26503 ( .IN1(n23547), .IN2(n23546), .IN3(n23545), .IN4(n23544), 
        .QN(n23553) );
  OA22X1 U26504 ( .IN1(n13698), .IN2(n32714), .IN3(n13693), .IN4(n33536), .Q(
        n23551) );
  OA22X1 U26505 ( .IN1(n13691), .IN2(n32944), .IN3(n13685), .IN4(n30008), .Q(
        n23550) );
  OA22X1 U26506 ( .IN1(n13696), .IN2(n32138), .IN3(n13681), .IN4(n31332), .Q(
        n23549) );
  OA22X1 U26507 ( .IN1(n13692), .IN2(n33238), .IN3(n13684), .IN4(n29729), .Q(
        n23548) );
  NAND4X0 U26508 ( .IN1(n23551), .IN2(n23550), .IN3(n23549), .IN4(n23548), 
        .QN(n23552) );
  OA21X1 U26509 ( .IN1(n23553), .IN2(n23552), .IN3(n23622), .Q(\rf/N123 ) );
  OA22X1 U26510 ( .IN1(n13655), .IN2(n31332), .IN3(n13666), .IN4(n33238), .Q(
        n23557) );
  OA22X1 U26511 ( .IN1(n13658), .IN2(n29729), .IN3(n13653), .IN4(n30624), .Q(
        n23556) );
  OA22X1 U26512 ( .IN1(n13660), .IN2(n30329), .IN3(n13657), .IN4(n29387), .Q(
        n23555) );
  OA22X1 U26513 ( .IN1(n13665), .IN2(n32944), .IN3(n13668), .IN4(n33762), .Q(
        n23554) );
  NAND4X0 U26514 ( .IN1(n23557), .IN2(n23556), .IN3(n23555), .IN4(n23554), 
        .QN(n23563) );
  OA22X1 U26515 ( .IN1(n13672), .IN2(n32714), .IN3(n13669), .IN4(n31938), .Q(
        n23561) );
  OA22X1 U26516 ( .IN1(n13654), .IN2(n30975), .IN3(n13659), .IN4(n30008), .Q(
        n23560) );
  OA22X1 U26517 ( .IN1(n13656), .IN2(n31627), .IN3(n13670), .IN4(n32138), .Q(
        n23559) );
  OA22X1 U26518 ( .IN1(n13667), .IN2(n33536), .IN3(n13671), .IN4(n32456), .Q(
        n23558) );
  NAND4X0 U26519 ( .IN1(n23561), .IN2(n23560), .IN3(n23559), .IN4(n23558), 
        .QN(n23562) );
  OA21X1 U26520 ( .IN1(n23563), .IN2(n23562), .IN3(n23622), .Q(\rf/N124 ) );
  OA22X1 U26521 ( .IN1(n13639), .IN2(n32944), .IN3(n13646), .IN4(n32714), .Q(
        n23567) );
  OA22X1 U26522 ( .IN1(n13640), .IN2(n33238), .IN3(n13643), .IN4(n31938), .Q(
        n23566) );
  OA22X1 U26523 ( .IN1(n13645), .IN2(n32456), .IN3(n13641), .IN4(n33536), .Q(
        n23565) );
  OA22X1 U26524 ( .IN1(n13627), .IN2(n30624), .IN3(n13632), .IN4(n29729), .Q(
        n23564) );
  NAND4X0 U26525 ( .IN1(n23567), .IN2(n23566), .IN3(n23565), .IN4(n23564), 
        .QN(n23573) );
  OA22X1 U26526 ( .IN1(n13642), .IN2(n33762), .IN3(n13628), .IN4(n30975), .Q(
        n23571) );
  OA22X1 U26527 ( .IN1(n13631), .IN2(n29387), .IN3(n13630), .IN4(n31627), .Q(
        n23570) );
  OA22X1 U26528 ( .IN1(n13634), .IN2(n30329), .IN3(n13629), .IN4(n31332), .Q(
        n23569) );
  OA22X1 U26529 ( .IN1(n13633), .IN2(n30008), .IN3(n13644), .IN4(n32138), .Q(
        n23568) );
  NAND4X0 U26530 ( .IN1(n23571), .IN2(n23570), .IN3(n23569), .IN4(n23568), 
        .QN(n23572) );
  OA21X1 U26531 ( .IN1(n23573), .IN2(n23572), .IN3(n23622), .Q(\rf/N125 ) );
  OA22X1 U26532 ( .IN1(n13619), .IN2(n32456), .IN3(n13605), .IN4(n29387), .Q(
        n23577) );
  OA22X1 U26533 ( .IN1(n13614), .IN2(n33238), .IN3(n13602), .IN4(n30975), .Q(
        n23576) );
  OA22X1 U26534 ( .IN1(n13618), .IN2(n32138), .IN3(n13616), .IN4(n33762), .Q(
        n23575) );
  OA22X1 U26535 ( .IN1(n13606), .IN2(n29729), .IN3(n13620), .IN4(n32714), .Q(
        n23574) );
  NAND4X0 U26536 ( .IN1(n23577), .IN2(n23576), .IN3(n23575), .IN4(n23574), 
        .QN(n23583) );
  OA22X1 U26537 ( .IN1(n13608), .IN2(n30329), .IN3(n13604), .IN4(n31627), .Q(
        n23581) );
  OA22X1 U26538 ( .IN1(n13601), .IN2(n30624), .IN3(n13617), .IN4(n31938), .Q(
        n23580) );
  OA22X1 U26539 ( .IN1(n13607), .IN2(n30008), .IN3(n13603), .IN4(n31332), .Q(
        n23579) );
  OA22X1 U26540 ( .IN1(n13613), .IN2(n32944), .IN3(n13615), .IN4(n33536), .Q(
        n23578) );
  NAND4X0 U26541 ( .IN1(n23581), .IN2(n23580), .IN3(n23579), .IN4(n23578), 
        .QN(n23582) );
  OA21X1 U26542 ( .IN1(n23583), .IN2(n23582), .IN3(n23622), .Q(\rf/N126 ) );
  OA22X1 U26543 ( .IN1(n13592), .IN2(n32138), .IN3(n13575), .IN4(n30624), .Q(
        n23587) );
  OA22X1 U26544 ( .IN1(n13579), .IN2(n29387), .IN3(n13594), .IN4(n32714), .Q(
        n23586) );
  OA22X1 U26545 ( .IN1(n13578), .IN2(n31627), .IN3(n13591), .IN4(n31938), .Q(
        n23585) );
  OA22X1 U26546 ( .IN1(n13587), .IN2(n32944), .IN3(n13589), .IN4(n33536), .Q(
        n23584) );
  NAND4X0 U26547 ( .IN1(n23587), .IN2(n23586), .IN3(n23585), .IN4(n23584), 
        .QN(n23593) );
  OA22X1 U26548 ( .IN1(n13582), .IN2(n30329), .IN3(n13593), .IN4(n32456), .Q(
        n23591) );
  OA22X1 U26549 ( .IN1(n13580), .IN2(n29729), .IN3(n13576), .IN4(n30975), .Q(
        n23590) );
  OA22X1 U26550 ( .IN1(n13588), .IN2(n33238), .IN3(n13590), .IN4(n33762), .Q(
        n23589) );
  OA22X1 U26551 ( .IN1(n13581), .IN2(n30008), .IN3(n13577), .IN4(n31332), .Q(
        n23588) );
  NAND4X0 U26552 ( .IN1(n23591), .IN2(n23590), .IN3(n23589), .IN4(n23588), 
        .QN(n23592) );
  OA21X1 U26553 ( .IN1(n23593), .IN2(n23592), .IN3(n23622), .Q(\rf/N127 ) );
  OA22X1 U26554 ( .IN1(n13551), .IN2(n31332), .IN3(n13550), .IN4(n30975), .Q(
        n23597) );
  OA22X1 U26555 ( .IN1(n13568), .IN2(n32714), .IN3(n13563), .IN4(n33536), .Q(
        n23596) );
  OA22X1 U26556 ( .IN1(n13567), .IN2(n32456), .IN3(n13549), .IN4(n30624), .Q(
        n23595) );
  OA22X1 U26557 ( .IN1(n13566), .IN2(n32138), .IN3(n13555), .IN4(n30008), .Q(
        n23594) );
  NAND4X0 U26558 ( .IN1(n23597), .IN2(n23596), .IN3(n23595), .IN4(n23594), 
        .QN(n23603) );
  OA22X1 U26559 ( .IN1(n13564), .IN2(n33762), .IN3(n13565), .IN4(n31938), .Q(
        n23601) );
  OA22X1 U26560 ( .IN1(n13552), .IN2(n31627), .IN3(n13553), .IN4(n29387), .Q(
        n23600) );
  OA22X1 U26561 ( .IN1(n13556), .IN2(n30329), .IN3(n13554), .IN4(n29729), .Q(
        n23599) );
  OA22X1 U26562 ( .IN1(n13562), .IN2(n33238), .IN3(n13561), .IN4(n32944), .Q(
        n23598) );
  NAND4X0 U26563 ( .IN1(n23601), .IN2(n23600), .IN3(n23599), .IN4(n23598), 
        .QN(n23602) );
  OA21X1 U26564 ( .IN1(n23603), .IN2(n23602), .IN3(n23622), .Q(\rf/N128 ) );
  OA22X1 U26565 ( .IN1(n13538), .IN2(n33762), .IN3(n13526), .IN4(n31627), .Q(
        n23607) );
  OA22X1 U26566 ( .IN1(n13523), .IN2(n30624), .IN3(n13528), .IN4(n29729), .Q(
        n23606) );
  OA22X1 U26567 ( .IN1(n13539), .IN2(n31938), .IN3(n13541), .IN4(n32456), .Q(
        n23605) );
  OA22X1 U26568 ( .IN1(n13542), .IN2(n32714), .IN3(n13529), .IN4(n30008), .Q(
        n23604) );
  NAND4X0 U26569 ( .IN1(n23607), .IN2(n23606), .IN3(n23605), .IN4(n23604), 
        .QN(n23613) );
  OA22X1 U26570 ( .IN1(n13530), .IN2(n30329), .IN3(n13527), .IN4(n29387), .Q(
        n23611) );
  OA22X1 U26571 ( .IN1(n13535), .IN2(n32944), .IN3(n13537), .IN4(n33536), .Q(
        n23610) );
  OA22X1 U26572 ( .IN1(n13540), .IN2(n32138), .IN3(n13525), .IN4(n31332), .Q(
        n23609) );
  OA22X1 U26573 ( .IN1(n13524), .IN2(n30975), .IN3(n13536), .IN4(n33238), .Q(
        n23608) );
  NAND4X0 U26574 ( .IN1(n23611), .IN2(n23610), .IN3(n23609), .IN4(n23608), 
        .QN(n23612) );
  OA21X1 U26575 ( .IN1(n23613), .IN2(n23612), .IN3(n23622), .Q(\rf/N129 ) );
  OA22X1 U26576 ( .IN1(n13469), .IN2(n31332), .IN3(n13464), .IN4(n30624), .Q(
        n23617) );
  OA22X1 U26577 ( .IN1(n13494), .IN2(n32456), .IN3(n13482), .IN4(n33238), .Q(
        n23616) );
  OA22X1 U26578 ( .IN1(n13484), .IN2(n33536), .IN3(n13465), .IN4(n30975), .Q(
        n23615) );
  OA22X1 U26579 ( .IN1(n13471), .IN2(n29387), .IN3(n13495), .IN4(n32714), .Q(
        n23614) );
  NAND4X0 U26580 ( .IN1(n23617), .IN2(n23616), .IN3(n23615), .IN4(n23614), 
        .QN(n23624) );
  OA22X1 U26581 ( .IN1(n13475), .IN2(n30329), .IN3(n13489), .IN4(n31938), .Q(
        n23621) );
  OA22X1 U26582 ( .IN1(n13470), .IN2(n31627), .IN3(n13485), .IN4(n33762), .Q(
        n23620) );
  OA22X1 U26583 ( .IN1(n13474), .IN2(n30008), .IN3(n13490), .IN4(n32138), .Q(
        n23619) );
  OA22X1 U26584 ( .IN1(n13481), .IN2(n32944), .IN3(n13472), .IN4(n29729), .Q(
        n23618) );
  NAND4X0 U26585 ( .IN1(n23621), .IN2(n23620), .IN3(n23619), .IN4(n23618), 
        .QN(n23623) );
  OA21X1 U26586 ( .IN1(n23624), .IN2(n23623), .IN3(n23622), .Q(\rf/N130 ) );
  NAND4X0 U26587 ( .IN1(n23628), .IN2(n23627), .IN3(n23626), .IN4(n23625), 
        .QN(n23634) );
  NAND4X0 U26588 ( .IN1(n23632), .IN2(n23631), .IN3(n23630), .IN4(n23629), 
        .QN(n23633) );
  OR2X1 U26589 ( .IN1(n23634), .IN2(n23633), .Q(s15_stb_o) );
  INVX0 U26590 ( .INP(m4s0_data_o[16]), .ZN(n28329) );
  INVX0 U26591 ( .INP(m7s0_data_o[16]), .ZN(n28327) );
  OA22X1 U26592 ( .IN1(n23825), .IN2(n28329), .IN3(n23824), .IN4(n28327), .Q(
        n23638) );
  INVX0 U26593 ( .INP(m5s0_data_o[16]), .ZN(n28325) );
  INVX0 U26594 ( .INP(m2s0_data_o[16]), .ZN(n28331) );
  OA22X1 U26595 ( .IN1(n23832), .IN2(n28325), .IN3(n23837), .IN4(n28331), .Q(
        n23637) );
  INVX0 U26596 ( .INP(m3s0_data_o[16]), .ZN(n28326) );
  INVX0 U26597 ( .INP(m1s0_data_o[16]), .ZN(n28332) );
  OA22X1 U26598 ( .IN1(n23812), .IN2(n28326), .IN3(n23831), .IN4(n28332), .Q(
        n23636) );
  INVX0 U26599 ( .INP(m0s0_data_o[16]), .ZN(n28330) );
  INVX0 U26600 ( .INP(m6s0_data_o[16]), .ZN(n28328) );
  OA22X1 U26601 ( .IN1(n23838), .IN2(n28330), .IN3(n23833), .IN4(n28328), .Q(
        n23635) );
  NAND4X0 U26602 ( .IN1(n23638), .IN2(n23637), .IN3(n23636), .IN4(n23635), 
        .QN(s15_data_o[16]) );
  INVX0 U26603 ( .INP(m6s0_data_o[17]), .ZN(n28343) );
  INVX0 U26604 ( .INP(m1s0_data_o[17]), .ZN(n28344) );
  OA22X1 U26605 ( .IN1(n23799), .IN2(n28343), .IN3(n23831), .IN4(n28344), .Q(
        n23642) );
  INVX0 U26606 ( .INP(m3s0_data_o[17]), .ZN(n28338) );
  INVX0 U26607 ( .INP(m7s0_data_o[17]), .ZN(n28341) );
  OA22X1 U26608 ( .IN1(n23812), .IN2(n28338), .IN3(n23824), .IN4(n28341), .Q(
        n23641) );
  INVX0 U26609 ( .INP(m0s0_data_o[17]), .ZN(n28340) );
  INVX0 U26610 ( .INP(m5s0_data_o[17]), .ZN(n28339) );
  OA22X1 U26611 ( .IN1(n23823), .IN2(n28340), .IN3(n23832), .IN4(n28339), .Q(
        n23640) );
  INVX0 U26612 ( .INP(m4s0_data_o[17]), .ZN(n28337) );
  INVX0 U26613 ( .INP(m2s0_data_o[17]), .ZN(n28342) );
  OA22X1 U26614 ( .IN1(n23836), .IN2(n28337), .IN3(n23817), .IN4(n28342), .Q(
        n23639) );
  NAND4X0 U26615 ( .IN1(n23642), .IN2(n23641), .IN3(n23640), .IN4(n23639), 
        .QN(s15_data_o[17]) );
  INVX0 U26616 ( .INP(m4s0_data_o[18]), .ZN(n28354) );
  INVX0 U26617 ( .INP(m5s0_data_o[18]), .ZN(n28349) );
  OA22X1 U26618 ( .IN1(n23825), .IN2(n28354), .IN3(n23826), .IN4(n28349), .Q(
        n23646) );
  INVX0 U26619 ( .INP(m6s0_data_o[18]), .ZN(n28351) );
  INVX0 U26620 ( .INP(m1s0_data_o[18]), .ZN(n28356) );
  OA22X1 U26621 ( .IN1(n23799), .IN2(n28351), .IN3(n23831), .IN4(n28356), .Q(
        n23645) );
  INVX0 U26622 ( .INP(m0s0_data_o[18]), .ZN(n28352) );
  INVX0 U26623 ( .INP(m3s0_data_o[18]), .ZN(n28355) );
  OA22X1 U26624 ( .IN1(n23838), .IN2(n28352), .IN3(n23835), .IN4(n28355), .Q(
        n23644) );
  INVX0 U26625 ( .INP(m7s0_data_o[18]), .ZN(n28353) );
  INVX0 U26626 ( .INP(m2s0_data_o[18]), .ZN(n28350) );
  OA22X1 U26627 ( .IN1(n23824), .IN2(n28353), .IN3(n23837), .IN4(n28350), .Q(
        n23643) );
  NAND4X0 U26628 ( .IN1(n23646), .IN2(n23645), .IN3(n23644), .IN4(n23643), 
        .QN(s15_data_o[18]) );
  INVX0 U26629 ( .INP(m0s0_data_o[19]), .ZN(n28366) );
  INVX0 U26630 ( .INP(m2s0_data_o[19]), .ZN(n28362) );
  OA22X1 U26631 ( .IN1(n23823), .IN2(n28366), .IN3(n23837), .IN4(n28362), .Q(
        n23650) );
  INVX0 U26632 ( .INP(m5s0_data_o[19]), .ZN(n28361) );
  INVX0 U26633 ( .INP(m7s0_data_o[19]), .ZN(n28367) );
  OA22X1 U26634 ( .IN1(n23832), .IN2(n28361), .IN3(n23824), .IN4(n28367), .Q(
        n23649) );
  INVX0 U26635 ( .INP(m4s0_data_o[19]), .ZN(n28365) );
  INVX0 U26636 ( .INP(m1s0_data_o[19]), .ZN(n28364) );
  OA22X1 U26637 ( .IN1(n23825), .IN2(n28365), .IN3(n23831), .IN4(n28364), .Q(
        n23648) );
  INVX0 U26638 ( .INP(m3s0_data_o[19]), .ZN(n28363) );
  INVX0 U26639 ( .INP(m6s0_data_o[19]), .ZN(n28368) );
  OA22X1 U26640 ( .IN1(n23835), .IN2(n28363), .IN3(n23833), .IN4(n28368), .Q(
        n23647) );
  NAND4X0 U26641 ( .IN1(n23650), .IN2(n23649), .IN3(n23648), .IN4(n23647), 
        .QN(s15_data_o[19]) );
  INVX0 U26642 ( .INP(m0s0_data_o[20]), .ZN(n28378) );
  INVX0 U26643 ( .INP(m3s0_data_o[20]), .ZN(n28373) );
  OA22X1 U26644 ( .IN1(n23838), .IN2(n28378), .IN3(n23835), .IN4(n28373), .Q(
        n23654) );
  INVX0 U26645 ( .INP(m6s0_data_o[20]), .ZN(n28379) );
  INVX0 U26646 ( .INP(m2s0_data_o[20]), .ZN(n28374) );
  OA22X1 U26647 ( .IN1(n23799), .IN2(n28379), .IN3(n23817), .IN4(n28374), .Q(
        n23653) );
  INVX0 U26648 ( .INP(m7s0_data_o[20]), .ZN(n28375) );
  INVX0 U26649 ( .INP(m1s0_data_o[20]), .ZN(n28377) );
  OA22X1 U26650 ( .IN1(n23834), .IN2(n28375), .IN3(n23831), .IN4(n28377), .Q(
        n23652) );
  INVX0 U26651 ( .INP(m4s0_data_o[20]), .ZN(n28376) );
  INVX0 U26652 ( .INP(m5s0_data_o[20]), .ZN(n28380) );
  OA22X1 U26653 ( .IN1(n23836), .IN2(n28376), .IN3(n23826), .IN4(n28380), .Q(
        n23651) );
  NAND4X0 U26654 ( .IN1(n23654), .IN2(n23653), .IN3(n23652), .IN4(n23651), 
        .QN(s15_data_o[20]) );
  INVX0 U26655 ( .INP(m6s0_data_o[21]), .ZN(n28389) );
  INVX0 U26656 ( .INP(m1s0_data_o[21]), .ZN(n28386) );
  OA22X1 U26657 ( .IN1(n23799), .IN2(n28389), .IN3(n23831), .IN4(n28386), .Q(
        n23658) );
  INVX0 U26658 ( .INP(m0s0_data_o[21]), .ZN(n28392) );
  INVX0 U26659 ( .INP(m2s0_data_o[21]), .ZN(n28390) );
  OA22X1 U26660 ( .IN1(n23823), .IN2(n28392), .IN3(n23817), .IN4(n28390), .Q(
        n23657) );
  INVX0 U26661 ( .INP(m5s0_data_o[21]), .ZN(n28385) );
  INVX0 U26662 ( .INP(m3s0_data_o[21]), .ZN(n28388) );
  OA22X1 U26663 ( .IN1(n23832), .IN2(n28385), .IN3(n23835), .IN4(n28388), .Q(
        n23656) );
  INVX0 U26664 ( .INP(m4s0_data_o[21]), .ZN(n28387) );
  INVX0 U26665 ( .INP(m7s0_data_o[21]), .ZN(n28391) );
  OA22X1 U26666 ( .IN1(n23836), .IN2(n28387), .IN3(n23824), .IN4(n28391), .Q(
        n23655) );
  NAND4X0 U26667 ( .IN1(n23658), .IN2(n23657), .IN3(n23656), .IN4(n23655), 
        .QN(s15_data_o[21]) );
  INVX0 U26668 ( .INP(m4s0_data_o[22]), .ZN(n28398) );
  INVX0 U26669 ( .INP(m3s0_data_o[22]), .ZN(n28403) );
  OA22X1 U26670 ( .IN1(n23825), .IN2(n28398), .IN3(n23835), .IN4(n28403), .Q(
        n23662) );
  INVX0 U26671 ( .INP(m1s0_data_o[22]), .ZN(n28402) );
  INVX0 U26672 ( .INP(m2s0_data_o[22]), .ZN(n28404) );
  OA22X1 U26673 ( .IN1(n23818), .IN2(n28402), .IN3(n23837), .IN4(n28404), .Q(
        n23661) );
  INVX0 U26674 ( .INP(m5s0_data_o[22]), .ZN(n28399) );
  INVX0 U26675 ( .INP(m7s0_data_o[22]), .ZN(n28397) );
  OA22X1 U26676 ( .IN1(n23832), .IN2(n28399), .IN3(n23824), .IN4(n28397), .Q(
        n23660) );
  INVX0 U26677 ( .INP(m0s0_data_o[22]), .ZN(n28400) );
  INVX0 U26678 ( .INP(m6s0_data_o[22]), .ZN(n28401) );
  OA22X1 U26679 ( .IN1(n23838), .IN2(n28400), .IN3(n23799), .IN4(n28401), .Q(
        n23659) );
  NAND4X0 U26680 ( .IN1(n23662), .IN2(n23661), .IN3(n23660), .IN4(n23659), 
        .QN(s15_data_o[22]) );
  INVX0 U26681 ( .INP(m7s0_data_o[23]), .ZN(n28411) );
  INVX0 U26682 ( .INP(m2s0_data_o[23]), .ZN(n28414) );
  OA22X1 U26683 ( .IN1(n23834), .IN2(n28411), .IN3(n23817), .IN4(n28414), .Q(
        n23666) );
  INVX0 U26684 ( .INP(m0s0_data_o[23]), .ZN(n28416) );
  INVX0 U26685 ( .INP(m3s0_data_o[23]), .ZN(n28413) );
  OA22X1 U26686 ( .IN1(n23823), .IN2(n28416), .IN3(n23835), .IN4(n28413), .Q(
        n23665) );
  INVX0 U26687 ( .INP(m4s0_data_o[23]), .ZN(n28410) );
  INVX0 U26688 ( .INP(m5s0_data_o[23]), .ZN(n28412) );
  OA22X1 U26689 ( .IN1(n23825), .IN2(n28410), .IN3(n23832), .IN4(n28412), .Q(
        n23664) );
  INVX0 U26690 ( .INP(m6s0_data_o[23]), .ZN(n28409) );
  INVX0 U26691 ( .INP(m1s0_data_o[23]), .ZN(n28415) );
  OA22X1 U26692 ( .IN1(n23799), .IN2(n28409), .IN3(n23831), .IN4(n28415), .Q(
        n23663) );
  NAND4X0 U26693 ( .IN1(n23666), .IN2(n23665), .IN3(n23664), .IN4(n23663), 
        .QN(s15_data_o[23]) );
  INVX0 U26694 ( .INP(m0s0_data_o[24]), .ZN(n28426) );
  INVX0 U26695 ( .INP(m2s0_data_o[24]), .ZN(n28422) );
  OA22X1 U26696 ( .IN1(n23838), .IN2(n28426), .IN3(n23837), .IN4(n28422), .Q(
        n23670) );
  INVX0 U26697 ( .INP(m7s0_data_o[24]), .ZN(n28423) );
  INVX0 U26698 ( .INP(m1s0_data_o[24]), .ZN(n28424) );
  OA22X1 U26699 ( .IN1(n23824), .IN2(n28423), .IN3(n23831), .IN4(n28424), .Q(
        n23669) );
  INVX0 U26700 ( .INP(m4s0_data_o[24]), .ZN(n28425) );
  INVX0 U26701 ( .INP(m5s0_data_o[24]), .ZN(n28428) );
  OA22X1 U26702 ( .IN1(n23836), .IN2(n28425), .IN3(n23826), .IN4(n28428), .Q(
        n23668) );
  INVX0 U26703 ( .INP(m3s0_data_o[24]), .ZN(n28421) );
  INVX0 U26704 ( .INP(m6s0_data_o[24]), .ZN(n28427) );
  OA22X1 U26705 ( .IN1(n23812), .IN2(n28421), .IN3(n23799), .IN4(n28427), .Q(
        n23667) );
  NAND4X0 U26706 ( .IN1(n23670), .IN2(n23669), .IN3(n23668), .IN4(n23667), 
        .QN(s15_data_o[24]) );
  INVX0 U26707 ( .INP(m6s0_data_o[25]), .ZN(n28436) );
  INVX0 U26708 ( .INP(m1s0_data_o[25]), .ZN(n28440) );
  OA22X1 U26709 ( .IN1(n23799), .IN2(n28436), .IN3(n23831), .IN4(n28440), .Q(
        n23674) );
  INVX0 U26710 ( .INP(m4s0_data_o[25]), .ZN(n28433) );
  INVX0 U26711 ( .INP(m5s0_data_o[25]), .ZN(n28437) );
  OA22X1 U26712 ( .IN1(n23825), .IN2(n28433), .IN3(n23832), .IN4(n28437), .Q(
        n23673) );
  INVX0 U26713 ( .INP(m0s0_data_o[25]), .ZN(n28438) );
  INVX0 U26714 ( .INP(m2s0_data_o[25]), .ZN(n28434) );
  OA22X1 U26715 ( .IN1(n23838), .IN2(n28438), .IN3(n23837), .IN4(n28434), .Q(
        n23672) );
  INVX0 U26716 ( .INP(m3s0_data_o[25]), .ZN(n28439) );
  INVX0 U26717 ( .INP(m7s0_data_o[25]), .ZN(n28435) );
  OA22X1 U26718 ( .IN1(n23835), .IN2(n28439), .IN3(n23824), .IN4(n28435), .Q(
        n23671) );
  NAND4X0 U26719 ( .IN1(n23674), .IN2(n23673), .IN3(n23672), .IN4(n23671), 
        .QN(s15_data_o[25]) );
  INVX0 U26720 ( .INP(m3s0_data_o[26]), .ZN(n28446) );
  INVX0 U26721 ( .INP(m6s0_data_o[26]), .ZN(n28447) );
  OA22X1 U26722 ( .IN1(n23812), .IN2(n28446), .IN3(n23799), .IN4(n28447), .Q(
        n23678) );
  INVX0 U26723 ( .INP(m4s0_data_o[26]), .ZN(n28449) );
  INVX0 U26724 ( .INP(m1s0_data_o[26]), .ZN(n28451) );
  OA22X1 U26725 ( .IN1(n23825), .IN2(n28449), .IN3(n23831), .IN4(n28451), .Q(
        n23677) );
  INVX0 U26726 ( .INP(m5s0_data_o[26]), .ZN(n28448) );
  INVX0 U26727 ( .INP(m2s0_data_o[26]), .ZN(n28450) );
  OA22X1 U26728 ( .IN1(n23832), .IN2(n28448), .IN3(n23817), .IN4(n28450), .Q(
        n23676) );
  INVX0 U26729 ( .INP(m0s0_data_o[26]), .ZN(n28452) );
  INVX0 U26730 ( .INP(m7s0_data_o[26]), .ZN(n28445) );
  OA22X1 U26731 ( .IN1(n23838), .IN2(n28452), .IN3(n23824), .IN4(n28445), .Q(
        n23675) );
  NAND4X0 U26732 ( .IN1(n23678), .IN2(n23677), .IN3(n23676), .IN4(n23675), 
        .QN(s15_data_o[26]) );
  INVX0 U26733 ( .INP(m4s0_data_o[27]), .ZN(n28457) );
  INVX0 U26734 ( .INP(m5s0_data_o[27]), .ZN(n28463) );
  OA22X1 U26735 ( .IN1(n23825), .IN2(n28457), .IN3(n23832), .IN4(n28463), .Q(
        n23682) );
  INVX0 U26736 ( .INP(m0s0_data_o[27]), .ZN(n28462) );
  INVX0 U26737 ( .INP(m6s0_data_o[27]), .ZN(n28460) );
  OA22X1 U26738 ( .IN1(n23838), .IN2(n28462), .IN3(n23799), .IN4(n28460), .Q(
        n23681) );
  INVX0 U26739 ( .INP(m7s0_data_o[27]), .ZN(n28459) );
  INVX0 U26740 ( .INP(m1s0_data_o[27]), .ZN(n28461) );
  OA22X1 U26741 ( .IN1(n23834), .IN2(n28459), .IN3(n23831), .IN4(n28461), .Q(
        n23680) );
  INVX0 U26742 ( .INP(m3s0_data_o[27]), .ZN(n28458) );
  INVX0 U26743 ( .INP(m2s0_data_o[27]), .ZN(n28464) );
  OA22X1 U26744 ( .IN1(n23835), .IN2(n28458), .IN3(n23817), .IN4(n28464), .Q(
        n23679) );
  NAND4X0 U26745 ( .IN1(n23682), .IN2(n23681), .IN3(n23680), .IN4(n23679), 
        .QN(s15_data_o[27]) );
  INVX0 U26746 ( .INP(m4s0_data_o[28]), .ZN(n28471) );
  INVX0 U26747 ( .INP(m3s0_data_o[28]), .ZN(n28470) );
  OA22X1 U26748 ( .IN1(n23825), .IN2(n28471), .IN3(n23835), .IN4(n28470), .Q(
        n23686) );
  INVX0 U26749 ( .INP(m6s0_data_o[28]), .ZN(n28469) );
  INVX0 U26750 ( .INP(m1s0_data_o[28]), .ZN(n28476) );
  OA22X1 U26751 ( .IN1(n23799), .IN2(n28469), .IN3(n23831), .IN4(n28476), .Q(
        n23685) );
  INVX0 U26752 ( .INP(m0s0_data_o[28]), .ZN(n28474) );
  INVX0 U26753 ( .INP(m5s0_data_o[28]), .ZN(n28475) );
  OA22X1 U26754 ( .IN1(n23838), .IN2(n28474), .IN3(n23832), .IN4(n28475), .Q(
        n23684) );
  INVX0 U26755 ( .INP(m7s0_data_o[28]), .ZN(n28473) );
  INVX0 U26756 ( .INP(m2s0_data_o[28]), .ZN(n28472) );
  OA22X1 U26757 ( .IN1(n23824), .IN2(n28473), .IN3(n23817), .IN4(n28472), .Q(
        n23683) );
  NAND4X0 U26758 ( .IN1(n23686), .IN2(n23685), .IN3(n23684), .IN4(n23683), 
        .QN(s15_data_o[28]) );
  INVX0 U26759 ( .INP(m7s0_data_o[29]), .ZN(n28481) );
  INVX0 U26760 ( .INP(m1s0_data_o[29]), .ZN(n28482) );
  OA22X1 U26761 ( .IN1(n23834), .IN2(n28481), .IN3(n23831), .IN4(n28482), .Q(
        n23690) );
  INVX0 U26762 ( .INP(m3s0_data_o[29]), .ZN(n28486) );
  INVX0 U26763 ( .INP(m2s0_data_o[29]), .ZN(n28488) );
  OA22X1 U26764 ( .IN1(n23812), .IN2(n28486), .IN3(n23817), .IN4(n28488), .Q(
        n23689) );
  INVX0 U26765 ( .INP(m4s0_data_o[29]), .ZN(n28487) );
  INVX0 U26766 ( .INP(m6s0_data_o[29]), .ZN(n28485) );
  OA22X1 U26767 ( .IN1(n23825), .IN2(n28487), .IN3(n23799), .IN4(n28485), .Q(
        n23688) );
  INVX0 U26768 ( .INP(m0s0_data_o[29]), .ZN(n28484) );
  INVX0 U26769 ( .INP(m5s0_data_o[29]), .ZN(n28483) );
  OA22X1 U26770 ( .IN1(n23838), .IN2(n28484), .IN3(n23826), .IN4(n28483), .Q(
        n23687) );
  NAND4X0 U26771 ( .IN1(n23690), .IN2(n23689), .IN3(n23688), .IN4(n23687), 
        .QN(s15_data_o[29]) );
  INVX0 U26772 ( .INP(m5s0_data_o[30]), .ZN(n28495) );
  INVX0 U26773 ( .INP(m6s0_data_o[30]), .ZN(n28500) );
  OA22X1 U26774 ( .IN1(n23832), .IN2(n28495), .IN3(n23799), .IN4(n28500), .Q(
        n23694) );
  INVX0 U26775 ( .INP(m1s0_data_o[30]), .ZN(n28498) );
  INVX0 U26776 ( .INP(m2s0_data_o[30]), .ZN(n28497) );
  OA22X1 U26777 ( .IN1(n23818), .IN2(n28498), .IN3(n23817), .IN4(n28497), .Q(
        n23693) );
  INVX0 U26778 ( .INP(m0s0_data_o[30]), .ZN(n28494) );
  INVX0 U26779 ( .INP(m3s0_data_o[30]), .ZN(n28496) );
  OA22X1 U26780 ( .IN1(n23838), .IN2(n28494), .IN3(n23835), .IN4(n28496), .Q(
        n23692) );
  INVX0 U26781 ( .INP(m4s0_data_o[30]), .ZN(n28493) );
  INVX0 U26782 ( .INP(m7s0_data_o[30]), .ZN(n28499) );
  OA22X1 U26783 ( .IN1(n23825), .IN2(n28493), .IN3(n23834), .IN4(n28499), .Q(
        n23691) );
  NAND4X0 U26784 ( .IN1(n23694), .IN2(n23693), .IN3(n23692), .IN4(n23691), 
        .QN(s15_data_o[30]) );
  INVX0 U26785 ( .INP(m0s0_data_o[31]), .ZN(n28510) );
  INVX0 U26786 ( .INP(m3s0_data_o[31]), .ZN(n28505) );
  OA22X1 U26787 ( .IN1(n23838), .IN2(n28510), .IN3(n23835), .IN4(n28505), .Q(
        n23698) );
  INVX0 U26788 ( .INP(m5s0_data_o[31]), .ZN(n28508) );
  INVX0 U26789 ( .INP(m6s0_data_o[31]), .ZN(n28511) );
  OA22X1 U26790 ( .IN1(n23832), .IN2(n28508), .IN3(n23799), .IN4(n28511), .Q(
        n23697) );
  INVX0 U26791 ( .INP(m7s0_data_o[31]), .ZN(n28507) );
  INVX0 U26792 ( .INP(m2s0_data_o[31]), .ZN(n28506) );
  OA22X1 U26793 ( .IN1(n23824), .IN2(n28507), .IN3(n23817), .IN4(n28506), .Q(
        n23696) );
  INVX0 U26794 ( .INP(m4s0_data_o[31]), .ZN(n28512) );
  INVX0 U26795 ( .INP(m1s0_data_o[31]), .ZN(n28509) );
  OA22X1 U26796 ( .IN1(n23825), .IN2(n28512), .IN3(n23831), .IN4(n28509), .Q(
        n23695) );
  NAND4X0 U26797 ( .IN1(n23698), .IN2(n23697), .IN3(n23696), .IN4(n23695), 
        .QN(s15_data_o[31]) );
  INVX0 U26798 ( .INP(m3s0_sel[0]), .ZN(n28524) );
  INVX0 U26799 ( .INP(m6s0_sel[0]), .ZN(n28521) );
  OA22X1 U26800 ( .IN1(n23812), .IN2(n28524), .IN3(n23799), .IN4(n28521), .Q(
        n23702) );
  INVX0 U26801 ( .INP(m5s0_sel[0]), .ZN(n28520) );
  INVX0 U26802 ( .INP(m1s0_sel[0]), .ZN(n28517) );
  OA22X1 U26803 ( .IN1(n23832), .IN2(n28520), .IN3(n23831), .IN4(n28517), .Q(
        n23701) );
  INVX0 U26804 ( .INP(m0s0_sel[0]), .ZN(n28518) );
  INVX0 U26805 ( .INP(m7s0_sel[0]), .ZN(n28519) );
  OA22X1 U26806 ( .IN1(n23838), .IN2(n28518), .IN3(n23824), .IN4(n28519), .Q(
        n23700) );
  INVX0 U26807 ( .INP(m4s0_sel[0]), .ZN(n28523) );
  INVX0 U26808 ( .INP(m2s0_sel[0]), .ZN(n28522) );
  OA22X1 U26809 ( .IN1(n23825), .IN2(n28523), .IN3(n23817), .IN4(n28522), .Q(
        n23699) );
  NAND4X0 U26810 ( .IN1(n23702), .IN2(n23701), .IN3(n23700), .IN4(n23699), 
        .QN(s15_sel_o[0]) );
  INVX0 U26811 ( .INP(m4s0_sel[1]), .ZN(n28535) );
  INVX0 U26812 ( .INP(m1s0_sel[1]), .ZN(n28532) );
  OA22X1 U26813 ( .IN1(n23836), .IN2(n28535), .IN3(n23818), .IN4(n28532), .Q(
        n23706) );
  INVX0 U26814 ( .INP(m0s0_sel[1]), .ZN(n28534) );
  INVX0 U26815 ( .INP(m5s0_sel[1]), .ZN(n28533) );
  OA22X1 U26816 ( .IN1(n23838), .IN2(n28534), .IN3(n23826), .IN4(n28533), .Q(
        n23705) );
  INVX0 U26817 ( .INP(m7s0_sel[1]), .ZN(n28529) );
  INVX0 U26818 ( .INP(m2s0_sel[1]), .ZN(n28530) );
  OA22X1 U26819 ( .IN1(n23834), .IN2(n28529), .IN3(n23817), .IN4(n28530), .Q(
        n23704) );
  INVX0 U26820 ( .INP(m3s0_sel[1]), .ZN(n28536) );
  INVX0 U26821 ( .INP(m6s0_sel[1]), .ZN(n28531) );
  OA22X1 U26822 ( .IN1(n23812), .IN2(n28536), .IN3(n23799), .IN4(n28531), .Q(
        n23703) );
  NAND4X0 U26823 ( .IN1(n23706), .IN2(n23705), .IN3(n23704), .IN4(n23703), 
        .QN(s15_sel_o[1]) );
  INVX0 U26824 ( .INP(m0s0_sel[2]), .ZN(n28544) );
  INVX0 U26825 ( .INP(m1s0_sel[2]), .ZN(n28546) );
  OA22X1 U26826 ( .IN1(n23838), .IN2(n28544), .IN3(n23831), .IN4(n28546), .Q(
        n23710) );
  INVX0 U26827 ( .INP(m5s0_sel[2]), .ZN(n28542) );
  INVX0 U26828 ( .INP(m6s0_sel[2]), .ZN(n28545) );
  OA22X1 U26829 ( .IN1(n23826), .IN2(n28542), .IN3(n23799), .IN4(n28545), .Q(
        n23709) );
  INVX0 U26830 ( .INP(m4s0_sel[2]), .ZN(n28547) );
  INVX0 U26831 ( .INP(m7s0_sel[2]), .ZN(n28541) );
  OA22X1 U26832 ( .IN1(n23836), .IN2(n28547), .IN3(n23834), .IN4(n28541), .Q(
        n23708) );
  INVX0 U26833 ( .INP(m3s0_sel[2]), .ZN(n28548) );
  INVX0 U26834 ( .INP(m2s0_sel[2]), .ZN(n28543) );
  OA22X1 U26835 ( .IN1(n23812), .IN2(n28548), .IN3(n23817), .IN4(n28543), .Q(
        n23707) );
  NAND4X0 U26836 ( .IN1(n23710), .IN2(n23709), .IN3(n23708), .IN4(n23707), 
        .QN(s15_sel_o[2]) );
  INVX0 U26837 ( .INP(m0s0_sel[3]), .ZN(n28558) );
  INVX0 U26838 ( .INP(m3s0_sel[3]), .ZN(n28557) );
  OA22X1 U26839 ( .IN1(n23838), .IN2(n28558), .IN3(n23835), .IN4(n28557), .Q(
        n23714) );
  INVX0 U26840 ( .INP(m4s0_sel[3]), .ZN(n28556) );
  INVX0 U26841 ( .INP(m5s0_sel[3]), .ZN(n28560) );
  OA22X1 U26842 ( .IN1(n23825), .IN2(n28556), .IN3(n23832), .IN4(n28560), .Q(
        n23713) );
  INVX0 U26843 ( .INP(m7s0_sel[3]), .ZN(n28555) );
  INVX0 U26844 ( .INP(m2s0_sel[3]), .ZN(n28553) );
  OA22X1 U26845 ( .IN1(n23834), .IN2(n28555), .IN3(n23817), .IN4(n28553), .Q(
        n23712) );
  INVX0 U26846 ( .INP(m6s0_sel[3]), .ZN(n28559) );
  INVX0 U26847 ( .INP(m1s0_sel[3]), .ZN(n28554) );
  OA22X1 U26848 ( .IN1(n23799), .IN2(n28559), .IN3(n23818), .IN4(n28554), .Q(
        n23711) );
  NAND4X0 U26849 ( .IN1(n23714), .IN2(n23713), .IN3(n23712), .IN4(n23711), 
        .QN(s15_sel_o[3]) );
  INVX0 U26850 ( .INP(m5s0_addr[0]), .ZN(n28567) );
  INVX0 U26851 ( .INP(m7s0_addr[0]), .ZN(n28569) );
  OA22X1 U26852 ( .IN1(n23826), .IN2(n28567), .IN3(n23824), .IN4(n28569), .Q(
        n23718) );
  INVX0 U26853 ( .INP(m0s0_addr[0]), .ZN(n28572) );
  INVX0 U26854 ( .INP(m4s0_addr[0]), .ZN(n28568) );
  OA22X1 U26855 ( .IN1(n23838), .IN2(n28572), .IN3(n23825), .IN4(n28568), .Q(
        n23717) );
  INVX0 U26856 ( .INP(m3s0_addr[0]), .ZN(n28566) );
  INVX0 U26857 ( .INP(m2s0_addr[0]), .ZN(n28571) );
  OA22X1 U26858 ( .IN1(n23812), .IN2(n28566), .IN3(n23817), .IN4(n28571), .Q(
        n23716) );
  INVX0 U26859 ( .INP(m6s0_addr[0]), .ZN(n28565) );
  INVX0 U26860 ( .INP(m1s0_addr[0]), .ZN(n28570) );
  OA22X1 U26861 ( .IN1(n23799), .IN2(n28565), .IN3(n23831), .IN4(n28570), .Q(
        n23715) );
  NAND4X0 U26862 ( .IN1(n23718), .IN2(n23717), .IN3(n23716), .IN4(n23715), 
        .QN(s15_addr_o[0]) );
  INVX0 U26863 ( .INP(m0s0_addr[1]), .ZN(n28580) );
  INVX0 U26864 ( .INP(m4s0_addr[1]), .ZN(n28579) );
  OA22X1 U26865 ( .IN1(n23838), .IN2(n28580), .IN3(n23836), .IN4(n28579), .Q(
        n23722) );
  INVX0 U26866 ( .INP(m7s0_addr[1]), .ZN(n28583) );
  INVX0 U26867 ( .INP(m1s0_addr[1]), .ZN(n28578) );
  OA22X1 U26868 ( .IN1(n23834), .IN2(n28583), .IN3(n23818), .IN4(n28578), .Q(
        n23721) );
  INVX0 U26869 ( .INP(m5s0_addr[1]), .ZN(n28584) );
  INVX0 U26870 ( .INP(m6s0_addr[1]), .ZN(n28577) );
  OA22X1 U26871 ( .IN1(n23826), .IN2(n28584), .IN3(n23799), .IN4(n28577), .Q(
        n23720) );
  INVX0 U26872 ( .INP(m3s0_addr[1]), .ZN(n28581) );
  INVX0 U26873 ( .INP(m2s0_addr[1]), .ZN(n28582) );
  OA22X1 U26874 ( .IN1(n23812), .IN2(n28581), .IN3(n23817), .IN4(n28582), .Q(
        n23719) );
  NAND4X0 U26875 ( .IN1(n23722), .IN2(n23721), .IN3(n23720), .IN4(n23719), 
        .QN(s15_addr_o[1]) );
  INVX0 U26876 ( .INP(m5s0_addr[6]), .ZN(n28637) );
  INVX0 U26877 ( .INP(m6s0_addr[6]), .ZN(n28641) );
  OA22X1 U26878 ( .IN1(n23832), .IN2(n28637), .IN3(n23833), .IN4(n28641), .Q(
        n23726) );
  INVX0 U26879 ( .INP(m0s0_addr[6]), .ZN(n28642) );
  INVX0 U26880 ( .INP(m4s0_addr[6]), .ZN(n28638) );
  OA22X1 U26881 ( .IN1(n23838), .IN2(n28642), .IN3(n23825), .IN4(n28638), .Q(
        n23725) );
  INVX0 U26882 ( .INP(m7s0_addr[6]), .ZN(n28639) );
  INVX0 U26883 ( .INP(m1s0_addr[6]), .ZN(n28640) );
  OA22X1 U26884 ( .IN1(n23834), .IN2(n28639), .IN3(n23831), .IN4(n28640), .Q(
        n23724) );
  INVX0 U26885 ( .INP(m3s0_addr[6]), .ZN(n28643) );
  INVX0 U26886 ( .INP(m2s0_addr[6]), .ZN(n28644) );
  OA22X1 U26887 ( .IN1(n23812), .IN2(n28643), .IN3(n23817), .IN4(n28644), .Q(
        n23723) );
  NAND4X0 U26888 ( .IN1(n23726), .IN2(n23725), .IN3(n23724), .IN4(n23723), 
        .QN(s15_addr_o[6]) );
  INVX0 U26889 ( .INP(m7s0_addr[7]), .ZN(n28655) );
  INVX0 U26890 ( .INP(m6s0_addr[7]), .ZN(n28651) );
  OA22X1 U26891 ( .IN1(n23834), .IN2(n28655), .IN3(n23833), .IN4(n28651), .Q(
        n23730) );
  INVX0 U26892 ( .INP(m4s0_addr[7]), .ZN(n28650) );
  INVX0 U26893 ( .INP(m2s0_addr[7]), .ZN(n28656) );
  OA22X1 U26894 ( .IN1(n23825), .IN2(n28650), .IN3(n23817), .IN4(n28656), .Q(
        n23729) );
  INVX0 U26895 ( .INP(m5s0_addr[7]), .ZN(n28649) );
  INVX0 U26896 ( .INP(m1s0_addr[7]), .ZN(n28652) );
  OA22X1 U26897 ( .IN1(n23826), .IN2(n28649), .IN3(n23818), .IN4(n28652), .Q(
        n23728) );
  INVX0 U26898 ( .INP(m0s0_addr[7]), .ZN(n28654) );
  INVX0 U26899 ( .INP(m3s0_addr[7]), .ZN(n28653) );
  OA22X1 U26900 ( .IN1(n23838), .IN2(n28654), .IN3(n23835), .IN4(n28653), .Q(
        n23727) );
  NAND4X0 U26901 ( .IN1(n23730), .IN2(n23729), .IN3(n23728), .IN4(n23727), 
        .QN(s15_addr_o[7]) );
  INVX0 U26902 ( .INP(m5s0_addr[8]), .ZN(n28662) );
  INVX0 U26903 ( .INP(m2s0_addr[8]), .ZN(n28666) );
  OA22X1 U26904 ( .IN1(n23826), .IN2(n28662), .IN3(n23817), .IN4(n28666), .Q(
        n23734) );
  INVX0 U26905 ( .INP(m4s0_addr[8]), .ZN(n28668) );
  INVX0 U26906 ( .INP(m3s0_addr[8]), .ZN(n28665) );
  OA22X1 U26907 ( .IN1(n23836), .IN2(n28668), .IN3(n23812), .IN4(n28665), .Q(
        n23733) );
  INVX0 U26908 ( .INP(m0s0_addr[8]), .ZN(n28664) );
  INVX0 U26909 ( .INP(m1s0_addr[8]), .ZN(n28663) );
  OA22X1 U26910 ( .IN1(n23838), .IN2(n28664), .IN3(n23831), .IN4(n28663), .Q(
        n23732) );
  INVX0 U26911 ( .INP(m7s0_addr[8]), .ZN(n28667) );
  INVX0 U26912 ( .INP(m6s0_addr[8]), .ZN(n28661) );
  OA22X1 U26913 ( .IN1(n23834), .IN2(n28667), .IN3(n23833), .IN4(n28661), .Q(
        n23731) );
  NAND4X0 U26914 ( .IN1(n23734), .IN2(n23733), .IN3(n23732), .IN4(n23731), 
        .QN(s15_addr_o[8]) );
  INVX0 U26915 ( .INP(m0s0_addr[9]), .ZN(n28680) );
  INVX0 U26916 ( .INP(m4s0_addr[9]), .ZN(n28673) );
  OA22X1 U26917 ( .IN1(n23838), .IN2(n28680), .IN3(n23836), .IN4(n28673), .Q(
        n23738) );
  INVX0 U26918 ( .INP(m6s0_addr[9]), .ZN(n28675) );
  INVX0 U26919 ( .INP(m1s0_addr[9]), .ZN(n28679) );
  OA22X1 U26920 ( .IN1(n23799), .IN2(n28675), .IN3(n23818), .IN4(n28679), .Q(
        n23737) );
  INVX0 U26921 ( .INP(m3s0_addr[9]), .ZN(n28676) );
  INVX0 U26922 ( .INP(m7s0_addr[9]), .ZN(n28677) );
  OA22X1 U26923 ( .IN1(n23812), .IN2(n28676), .IN3(n23824), .IN4(n28677), .Q(
        n23736) );
  INVX0 U26924 ( .INP(m5s0_addr[9]), .ZN(n28678) );
  INVX0 U26925 ( .INP(m2s0_addr[9]), .ZN(n28674) );
  OA22X1 U26926 ( .IN1(n23826), .IN2(n28678), .IN3(n23817), .IN4(n28674), .Q(
        n23735) );
  NAND4X0 U26927 ( .IN1(n23738), .IN2(n23737), .IN3(n23736), .IN4(n23735), 
        .QN(s15_addr_o[9]) );
  INVX0 U26928 ( .INP(m0s0_addr[10]), .ZN(n28692) );
  INVX0 U26929 ( .INP(m3s0_addr[10]), .ZN(n28687) );
  OA22X1 U26930 ( .IN1(n23823), .IN2(n28692), .IN3(n23812), .IN4(n28687), .Q(
        n23742) );
  INVX0 U26931 ( .INP(m1s0_addr[10]), .ZN(n28686) );
  INVX0 U26932 ( .INP(m2s0_addr[10]), .ZN(n28688) );
  OA22X1 U26933 ( .IN1(n23818), .IN2(n28686), .IN3(n23817), .IN4(n28688), .Q(
        n23741) );
  INVX0 U26934 ( .INP(m7s0_addr[10]), .ZN(n28689) );
  INVX0 U26935 ( .INP(m6s0_addr[10]), .ZN(n28690) );
  OA22X1 U26936 ( .IN1(n23834), .IN2(n28689), .IN3(n23833), .IN4(n28690), .Q(
        n23740) );
  INVX0 U26937 ( .INP(m4s0_addr[10]), .ZN(n28685) );
  INVX0 U26938 ( .INP(m5s0_addr[10]), .ZN(n28691) );
  OA22X1 U26939 ( .IN1(n23836), .IN2(n28685), .IN3(n23826), .IN4(n28691), .Q(
        n23739) );
  NAND4X0 U26940 ( .IN1(n23742), .IN2(n23741), .IN3(n23740), .IN4(n23739), 
        .QN(s15_addr_o[10]) );
  INVX0 U26941 ( .INP(m5s0_addr[11]), .ZN(n28703) );
  INVX0 U26942 ( .INP(m1s0_addr[11]), .ZN(n28698) );
  OA22X1 U26943 ( .IN1(n23826), .IN2(n28703), .IN3(n23831), .IN4(n28698), .Q(
        n23746) );
  INVX0 U26944 ( .INP(m0s0_addr[11]), .ZN(n28702) );
  INVX0 U26945 ( .INP(m2s0_addr[11]), .ZN(n28697) );
  OA22X1 U26946 ( .IN1(n23838), .IN2(n28702), .IN3(n23817), .IN4(n28697), .Q(
        n23745) );
  INVX0 U26947 ( .INP(m7s0_addr[11]), .ZN(n28699) );
  INVX0 U26948 ( .INP(m6s0_addr[11]), .ZN(n28700) );
  OA22X1 U26949 ( .IN1(n23834), .IN2(n28699), .IN3(n23833), .IN4(n28700), .Q(
        n23744) );
  INVX0 U26950 ( .INP(m4s0_addr[11]), .ZN(n28701) );
  INVX0 U26951 ( .INP(m3s0_addr[11]), .ZN(n28704) );
  OA22X1 U26952 ( .IN1(n23836), .IN2(n28701), .IN3(n23835), .IN4(n28704), .Q(
        n23743) );
  NAND4X0 U26953 ( .IN1(n23746), .IN2(n23745), .IN3(n23744), .IN4(n23743), 
        .QN(s15_addr_o[11]) );
  INVX0 U26954 ( .INP(m4s0_addr[12]), .ZN(n28709) );
  INVX0 U26955 ( .INP(m6s0_addr[12]), .ZN(n28711) );
  OA22X1 U26956 ( .IN1(n23836), .IN2(n28709), .IN3(n23833), .IN4(n28711), .Q(
        n23750) );
  INVX0 U26957 ( .INP(m0s0_addr[12]), .ZN(n28714) );
  INVX0 U26958 ( .INP(m2s0_addr[12]), .ZN(n28712) );
  OA22X1 U26959 ( .IN1(n23823), .IN2(n28714), .IN3(n23817), .IN4(n28712), .Q(
        n23749) );
  INVX0 U26960 ( .INP(m5s0_addr[12]), .ZN(n28715) );
  INVX0 U26961 ( .INP(m3s0_addr[12]), .ZN(n28716) );
  OA22X1 U26962 ( .IN1(n23826), .IN2(n28715), .IN3(n23835), .IN4(n28716), .Q(
        n23748) );
  INVX0 U26963 ( .INP(m7s0_addr[12]), .ZN(n28713) );
  INVX0 U26964 ( .INP(m1s0_addr[12]), .ZN(n28710) );
  OA22X1 U26965 ( .IN1(n23834), .IN2(n28713), .IN3(n23818), .IN4(n28710), .Q(
        n23747) );
  NAND4X0 U26966 ( .IN1(n23750), .IN2(n23749), .IN3(n23748), .IN4(n23747), 
        .QN(s15_addr_o[12]) );
  INVX0 U26967 ( .INP(m0s0_addr[13]), .ZN(n28722) );
  INVX0 U26968 ( .INP(m4s0_addr[13]), .ZN(n28723) );
  OA22X1 U26969 ( .IN1(n23823), .IN2(n28722), .IN3(n23825), .IN4(n28723), .Q(
        n23754) );
  INVX0 U26970 ( .INP(m6s0_addr[13]), .ZN(n28725) );
  INVX0 U26971 ( .INP(m1s0_addr[13]), .ZN(n28728) );
  OA22X1 U26972 ( .IN1(n23799), .IN2(n28725), .IN3(n23831), .IN4(n28728), .Q(
        n23753) );
  INVX0 U26973 ( .INP(m7s0_addr[13]), .ZN(n28727) );
  INVX0 U26974 ( .INP(m2s0_addr[13]), .ZN(n28726) );
  OA22X1 U26975 ( .IN1(n23834), .IN2(n28727), .IN3(n23817), .IN4(n28726), .Q(
        n23752) );
  INVX0 U26976 ( .INP(m5s0_addr[13]), .ZN(n28721) );
  INVX0 U26977 ( .INP(m3s0_addr[13]), .ZN(n28724) );
  OA22X1 U26978 ( .IN1(n23826), .IN2(n28721), .IN3(n23812), .IN4(n28724), .Q(
        n23751) );
  NAND4X0 U26979 ( .IN1(n23754), .IN2(n23753), .IN3(n23752), .IN4(n23751), 
        .QN(s15_addr_o[13]) );
  INVX0 U26980 ( .INP(m7s0_addr[14]), .ZN(n28739) );
  INVX0 U26981 ( .INP(m2s0_addr[14]), .ZN(n28736) );
  OA22X1 U26982 ( .IN1(n23834), .IN2(n28739), .IN3(n23837), .IN4(n28736), .Q(
        n23758) );
  INVX0 U26983 ( .INP(m4s0_addr[14]), .ZN(n28740) );
  INVX0 U26984 ( .INP(m1s0_addr[14]), .ZN(n28738) );
  OA22X1 U26985 ( .IN1(n23836), .IN2(n28740), .IN3(n23818), .IN4(n28738), .Q(
        n23757) );
  INVX0 U26986 ( .INP(m0s0_addr[14]), .ZN(n28734) );
  INVX0 U26987 ( .INP(m6s0_addr[14]), .ZN(n28733) );
  OA22X1 U26988 ( .IN1(n23838), .IN2(n28734), .IN3(n23833), .IN4(n28733), .Q(
        n23756) );
  INVX0 U26989 ( .INP(m5s0_addr[14]), .ZN(n28737) );
  INVX0 U26990 ( .INP(m3s0_addr[14]), .ZN(n28735) );
  OA22X1 U26991 ( .IN1(n23826), .IN2(n28737), .IN3(n23835), .IN4(n28735), .Q(
        n23755) );
  NAND4X0 U26992 ( .IN1(n23758), .IN2(n23757), .IN3(n23756), .IN4(n23755), 
        .QN(s15_addr_o[14]) );
  INVX0 U26993 ( .INP(m0s0_addr[15]), .ZN(n28746) );
  INVX0 U26994 ( .INP(m1s0_addr[15]), .ZN(n28748) );
  OA22X1 U26995 ( .IN1(n23838), .IN2(n28746), .IN3(n23831), .IN4(n28748), .Q(
        n23762) );
  INVX0 U26996 ( .INP(m4s0_addr[15]), .ZN(n28747) );
  INVX0 U26997 ( .INP(m2s0_addr[15]), .ZN(n28750) );
  OA22X1 U26998 ( .IN1(n23836), .IN2(n28747), .IN3(n23817), .IN4(n28750), .Q(
        n23761) );
  INVX0 U26999 ( .INP(m3s0_addr[15]), .ZN(n28752) );
  INVX0 U27000 ( .INP(m7s0_addr[15]), .ZN(n28745) );
  OA22X1 U27001 ( .IN1(n23812), .IN2(n28752), .IN3(n23834), .IN4(n28745), .Q(
        n23760) );
  INVX0 U27002 ( .INP(m5s0_addr[15]), .ZN(n28751) );
  INVX0 U27003 ( .INP(m6s0_addr[15]), .ZN(n28749) );
  OA22X1 U27004 ( .IN1(n23826), .IN2(n28751), .IN3(n23833), .IN4(n28749), .Q(
        n23759) );
  NAND4X0 U27005 ( .IN1(n23762), .IN2(n23761), .IN3(n23760), .IN4(n23759), 
        .QN(s15_addr_o[15]) );
  INVX0 U27006 ( .INP(m5s0_addr[16]), .ZN(n28757) );
  INVX0 U27007 ( .INP(m7s0_addr[16]), .ZN(n28763) );
  OA22X1 U27008 ( .IN1(n23826), .IN2(n28757), .IN3(n23824), .IN4(n28763), .Q(
        n23766) );
  INVX0 U27009 ( .INP(m4s0_addr[16]), .ZN(n28759) );
  INVX0 U27010 ( .INP(m1s0_addr[16]), .ZN(n28762) );
  OA22X1 U27011 ( .IN1(n23836), .IN2(n28759), .IN3(n23818), .IN4(n28762), .Q(
        n23765) );
  INVX0 U27012 ( .INP(m0s0_addr[16]), .ZN(n28758) );
  INVX0 U27013 ( .INP(m2s0_addr[16]), .ZN(n28760) );
  OA22X1 U27014 ( .IN1(n23823), .IN2(n28758), .IN3(n23837), .IN4(n28760), .Q(
        n23764) );
  INVX0 U27015 ( .INP(m3s0_addr[16]), .ZN(n28761) );
  INVX0 U27016 ( .INP(m6s0_addr[16]), .ZN(n28764) );
  OA22X1 U27017 ( .IN1(n23812), .IN2(n28761), .IN3(n23833), .IN4(n28764), .Q(
        n23763) );
  NAND4X0 U27018 ( .IN1(n23766), .IN2(n23765), .IN3(n23764), .IN4(n23763), 
        .QN(s15_addr_o[16]) );
  INVX0 U27019 ( .INP(m5s0_addr[17]), .ZN(n28771) );
  INVX0 U27020 ( .INP(m7s0_addr[17]), .ZN(n28769) );
  OA22X1 U27021 ( .IN1(n23826), .IN2(n28771), .IN3(n23824), .IN4(n28769), .Q(
        n23770) );
  INVX0 U27022 ( .INP(m4s0_addr[17]), .ZN(n28775) );
  INVX0 U27023 ( .INP(m3s0_addr[17]), .ZN(n28773) );
  OA22X1 U27024 ( .IN1(n23836), .IN2(n28775), .IN3(n23835), .IN4(n28773), .Q(
        n23769) );
  INVX0 U27025 ( .INP(m0s0_addr[17]), .ZN(n28772) );
  INVX0 U27026 ( .INP(m2s0_addr[17]), .ZN(n28774) );
  OA22X1 U27027 ( .IN1(n23838), .IN2(n28772), .IN3(n23817), .IN4(n28774), .Q(
        n23768) );
  INVX0 U27028 ( .INP(m6s0_addr[17]), .ZN(n28770) );
  INVX0 U27029 ( .INP(m1s0_addr[17]), .ZN(n28776) );
  OA22X1 U27030 ( .IN1(n23799), .IN2(n28770), .IN3(n23831), .IN4(n28776), .Q(
        n23767) );
  NAND4X0 U27031 ( .IN1(n23770), .IN2(n23769), .IN3(n23768), .IN4(n23767), 
        .QN(s15_addr_o[17]) );
  INVX0 U27032 ( .INP(m6s0_addr[18]), .ZN(n28785) );
  INVX0 U27033 ( .INP(m1s0_addr[18]), .ZN(n28788) );
  OA22X1 U27034 ( .IN1(n23799), .IN2(n28785), .IN3(n23818), .IN4(n28788), .Q(
        n23774) );
  INVX0 U27035 ( .INP(m0s0_addr[18]), .ZN(n28786) );
  INVX0 U27036 ( .INP(m4s0_addr[18]), .ZN(n28784) );
  OA22X1 U27037 ( .IN1(n23823), .IN2(n28786), .IN3(n23825), .IN4(n28784), .Q(
        n23773) );
  INVX0 U27038 ( .INP(m5s0_addr[18]), .ZN(n28783) );
  INVX0 U27039 ( .INP(m2s0_addr[18]), .ZN(n28787) );
  OA22X1 U27040 ( .IN1(n23826), .IN2(n28783), .IN3(n23837), .IN4(n28787), .Q(
        n23772) );
  INVX0 U27041 ( .INP(m3s0_addr[18]), .ZN(n28782) );
  INVX0 U27042 ( .INP(m7s0_addr[18]), .ZN(n28781) );
  OA22X1 U27043 ( .IN1(n23812), .IN2(n28782), .IN3(n23824), .IN4(n28781), .Q(
        n23771) );
  NAND4X0 U27044 ( .IN1(n23774), .IN2(n23773), .IN3(n23772), .IN4(n23771), 
        .QN(s15_addr_o[18]) );
  INVX0 U27045 ( .INP(m3s0_addr[19]), .ZN(n28794) );
  INVX0 U27046 ( .INP(m1s0_addr[19]), .ZN(n28800) );
  OA22X1 U27047 ( .IN1(n23812), .IN2(n28794), .IN3(n23818), .IN4(n28800), .Q(
        n23778) );
  INVX0 U27048 ( .INP(m0s0_addr[19]), .ZN(n28796) );
  INVX0 U27049 ( .INP(m2s0_addr[19]), .ZN(n28798) );
  OA22X1 U27050 ( .IN1(n23823), .IN2(n28796), .IN3(n23817), .IN4(n28798), .Q(
        n23777) );
  INVX0 U27051 ( .INP(m7s0_addr[19]), .ZN(n28799) );
  INVX0 U27052 ( .INP(m6s0_addr[19]), .ZN(n28793) );
  OA22X1 U27053 ( .IN1(n23834), .IN2(n28799), .IN3(n23833), .IN4(n28793), .Q(
        n23776) );
  INVX0 U27054 ( .INP(m4s0_addr[19]), .ZN(n28797) );
  INVX0 U27055 ( .INP(m5s0_addr[19]), .ZN(n28795) );
  OA22X1 U27056 ( .IN1(n23836), .IN2(n28797), .IN3(n23832), .IN4(n28795), .Q(
        n23775) );
  NAND4X0 U27057 ( .IN1(n23778), .IN2(n23777), .IN3(n23776), .IN4(n23775), 
        .QN(s15_addr_o[19]) );
  INVX0 U27058 ( .INP(m0s0_addr[20]), .ZN(n28812) );
  INVX0 U27059 ( .INP(m1s0_addr[20]), .ZN(n28808) );
  OA22X1 U27060 ( .IN1(n23838), .IN2(n28812), .IN3(n23831), .IN4(n28808), .Q(
        n23782) );
  INVX0 U27061 ( .INP(m3s0_addr[20]), .ZN(n28810) );
  INVX0 U27062 ( .INP(m7s0_addr[20]), .ZN(n28805) );
  OA22X1 U27063 ( .IN1(n23812), .IN2(n28810), .IN3(n23824), .IN4(n28805), .Q(
        n23781) );
  INVX0 U27064 ( .INP(m6s0_addr[20]), .ZN(n28809) );
  INVX0 U27065 ( .INP(m2s0_addr[20]), .ZN(n28807) );
  OA22X1 U27066 ( .IN1(n23799), .IN2(n28809), .IN3(n23837), .IN4(n28807), .Q(
        n23780) );
  INVX0 U27067 ( .INP(m4s0_addr[20]), .ZN(n28806) );
  INVX0 U27068 ( .INP(m5s0_addr[20]), .ZN(n28811) );
  OA22X1 U27069 ( .IN1(n23836), .IN2(n28806), .IN3(n23832), .IN4(n28811), .Q(
        n23779) );
  NAND4X0 U27070 ( .IN1(n23782), .IN2(n23781), .IN3(n23780), .IN4(n23779), 
        .QN(s15_addr_o[20]) );
  INVX0 U27071 ( .INP(m4s0_addr[21]), .ZN(n28821) );
  INVX0 U27072 ( .INP(m3s0_addr[21]), .ZN(n28819) );
  OA22X1 U27073 ( .IN1(n23836), .IN2(n28821), .IN3(n23835), .IN4(n28819), .Q(
        n23786) );
  INVX0 U27074 ( .INP(m7s0_addr[21]), .ZN(n28817) );
  INVX0 U27075 ( .INP(m6s0_addr[21]), .ZN(n28818) );
  OA22X1 U27076 ( .IN1(n23834), .IN2(n28817), .IN3(n23833), .IN4(n28818), .Q(
        n23785) );
  INVX0 U27077 ( .INP(m0s0_addr[21]), .ZN(n28822) );
  INVX0 U27078 ( .INP(m1s0_addr[21]), .ZN(n28824) );
  OA22X1 U27079 ( .IN1(n23838), .IN2(n28822), .IN3(n23818), .IN4(n28824), .Q(
        n23784) );
  INVX0 U27080 ( .INP(m5s0_addr[21]), .ZN(n28823) );
  INVX0 U27081 ( .INP(m2s0_addr[21]), .ZN(n28820) );
  OA22X1 U27082 ( .IN1(n23826), .IN2(n28823), .IN3(n23817), .IN4(n28820), .Q(
        n23783) );
  NAND4X0 U27083 ( .IN1(n23786), .IN2(n23785), .IN3(n23784), .IN4(n23783), 
        .QN(s15_addr_o[21]) );
  INVX0 U27084 ( .INP(m4s0_addr[22]), .ZN(n28836) );
  INVX0 U27085 ( .INP(m7s0_addr[22]), .ZN(n28829) );
  OA22X1 U27086 ( .IN1(n23836), .IN2(n28836), .IN3(n23834), .IN4(n28829), .Q(
        n23790) );
  INVX0 U27087 ( .INP(m6s0_addr[22]), .ZN(n28837) );
  INVX0 U27088 ( .INP(m2s0_addr[22]), .ZN(n28831) );
  OA22X1 U27089 ( .IN1(n23799), .IN2(n28837), .IN3(n23837), .IN4(n28831), .Q(
        n23789) );
  INVX0 U27090 ( .INP(m5s0_addr[22]), .ZN(n28834) );
  INVX0 U27091 ( .INP(m1s0_addr[22]), .ZN(n28832) );
  OA22X1 U27092 ( .IN1(n23826), .IN2(n28834), .IN3(n23818), .IN4(n28832), .Q(
        n23788) );
  INVX0 U27093 ( .INP(m0s0_addr[22]), .ZN(n28833) );
  INVX0 U27094 ( .INP(m3s0_addr[22]), .ZN(n28838) );
  OA22X1 U27095 ( .IN1(n23823), .IN2(n28833), .IN3(n23835), .IN4(n28838), .Q(
        n23787) );
  NAND4X0 U27096 ( .IN1(n23790), .IN2(n23789), .IN3(n23788), .IN4(n23787), 
        .QN(s15_addr_o[22]) );
  INVX0 U27097 ( .INP(m3s0_addr[23]), .ZN(n28850) );
  INVX0 U27098 ( .INP(m6s0_addr[23]), .ZN(n28846) );
  OA22X1 U27099 ( .IN1(n23812), .IN2(n28850), .IN3(n23833), .IN4(n28846), .Q(
        n23794) );
  INVX0 U27100 ( .INP(m7s0_addr[23]), .ZN(n28851) );
  INVX0 U27101 ( .INP(m2s0_addr[23]), .ZN(n28843) );
  OA22X1 U27102 ( .IN1(n23834), .IN2(n28851), .IN3(n23817), .IN4(n28843), .Q(
        n23793) );
  INVX0 U27103 ( .INP(m5s0_addr[23]), .ZN(n28849) );
  INVX0 U27104 ( .INP(m1s0_addr[23]), .ZN(n28845) );
  OA22X1 U27105 ( .IN1(n23826), .IN2(n28849), .IN3(n23831), .IN4(n28845), .Q(
        n23792) );
  INVX0 U27106 ( .INP(m0s0_addr[23]), .ZN(n28848) );
  INVX0 U27107 ( .INP(m4s0_addr[23]), .ZN(n28852) );
  OA22X1 U27108 ( .IN1(n23823), .IN2(n28848), .IN3(n23825), .IN4(n28852), .Q(
        n23791) );
  NAND4X0 U27109 ( .IN1(n23794), .IN2(n23793), .IN3(n23792), .IN4(n23791), 
        .QN(s15_addr_o[23]) );
  INVX0 U27110 ( .INP(m5s0_addr[24]), .ZN(n28859) );
  INVX0 U27111 ( .INP(m3s0_addr[24]), .ZN(n28857) );
  OA22X1 U27112 ( .IN1(n23826), .IN2(n28859), .IN3(n23812), .IN4(n28857), .Q(
        n23798) );
  INVX0 U27113 ( .INP(m0s0_addr[24]), .ZN(n28863) );
  INVX0 U27114 ( .INP(m7s0_addr[24]), .ZN(n28860) );
  OA22X1 U27115 ( .IN1(n23823), .IN2(n28863), .IN3(n23824), .IN4(n28860), .Q(
        n23797) );
  INVX0 U27116 ( .INP(m6s0_addr[24]), .ZN(n28865) );
  INVX0 U27117 ( .INP(m1s0_addr[24]), .ZN(n28864) );
  OA22X1 U27118 ( .IN1(n23799), .IN2(n28865), .IN3(n23831), .IN4(n28864), .Q(
        n23796) );
  INVX0 U27119 ( .INP(m4s0_addr[24]), .ZN(n28861) );
  INVX0 U27120 ( .INP(m2s0_addr[24]), .ZN(n28858) );
  OA22X1 U27121 ( .IN1(n23836), .IN2(n28861), .IN3(n23837), .IN4(n28858), .Q(
        n23795) );
  NAND4X0 U27122 ( .IN1(n23798), .IN2(n23797), .IN3(n23796), .IN4(n23795), 
        .QN(s15_addr_o[24]) );
  INVX0 U27123 ( .INP(m5s0_addr[25]), .ZN(n28876) );
  INVX0 U27124 ( .INP(m3s0_addr[25]), .ZN(n28874) );
  OA22X1 U27125 ( .IN1(n23826), .IN2(n28876), .IN3(n23835), .IN4(n28874), .Q(
        n23803) );
  INVX0 U27126 ( .INP(m0s0_addr[25]), .ZN(n28870) );
  INVX0 U27127 ( .INP(m4s0_addr[25]), .ZN(n28872) );
  OA22X1 U27128 ( .IN1(n23823), .IN2(n28870), .IN3(n23825), .IN4(n28872), .Q(
        n23802) );
  INVX0 U27129 ( .INP(m6s0_addr[25]), .ZN(n28871) );
  INVX0 U27130 ( .INP(m1s0_addr[25]), .ZN(n28877) );
  OA22X1 U27131 ( .IN1(n23799), .IN2(n28871), .IN3(n23818), .IN4(n28877), .Q(
        n23801) );
  INVX0 U27132 ( .INP(m7s0_addr[25]), .ZN(n28875) );
  INVX0 U27133 ( .INP(m2s0_addr[25]), .ZN(n28873) );
  OA22X1 U27134 ( .IN1(n23834), .IN2(n28875), .IN3(n23817), .IN4(n28873), .Q(
        n23800) );
  NAND4X0 U27135 ( .IN1(n23803), .IN2(n23802), .IN3(n23801), .IN4(n23800), 
        .QN(s15_addr_o[25]) );
  INVX0 U27136 ( .INP(m0s0_addr[26]), .ZN(n28884) );
  INVX0 U27137 ( .INP(m7s0_addr[26]), .ZN(n28889) );
  OA22X1 U27138 ( .IN1(n23823), .IN2(n28884), .IN3(n23834), .IN4(n28889), .Q(
        n23807) );
  INVX0 U27139 ( .INP(m1s0_addr[26]), .ZN(n28887) );
  INVX0 U27140 ( .INP(m2s0_addr[26]), .ZN(n28885) );
  OA22X1 U27141 ( .IN1(n23818), .IN2(n28887), .IN3(n23837), .IN4(n28885), .Q(
        n23806) );
  INVX0 U27142 ( .INP(m4s0_addr[26]), .ZN(n28886) );
  INVX0 U27143 ( .INP(m6s0_addr[26]), .ZN(n28883) );
  OA22X1 U27144 ( .IN1(n23836), .IN2(n28886), .IN3(n23833), .IN4(n28883), .Q(
        n23805) );
  INVX0 U27145 ( .INP(m5s0_addr[26]), .ZN(n28888) );
  INVX0 U27146 ( .INP(m3s0_addr[26]), .ZN(n28882) );
  OA22X1 U27147 ( .IN1(n23826), .IN2(n28888), .IN3(n23835), .IN4(n28882), .Q(
        n23804) );
  NAND4X0 U27148 ( .IN1(n23807), .IN2(n23806), .IN3(n23805), .IN4(n23804), 
        .QN(s15_addr_o[26]) );
  INVX0 U27149 ( .INP(m3s0_addr[27]), .ZN(n28901) );
  INVX0 U27150 ( .INP(m6s0_addr[27]), .ZN(n28897) );
  OA22X1 U27151 ( .IN1(n23812), .IN2(n28901), .IN3(n23833), .IN4(n28897), .Q(
        n23811) );
  INVX0 U27152 ( .INP(m4s0_addr[27]), .ZN(n28900) );
  INVX0 U27153 ( .INP(m2s0_addr[27]), .ZN(n28899) );
  OA22X1 U27154 ( .IN1(n23836), .IN2(n28900), .IN3(n23817), .IN4(n28899), .Q(
        n23810) );
  INVX0 U27155 ( .INP(m5s0_addr[27]), .ZN(n28896) );
  INVX0 U27156 ( .INP(m1s0_addr[27]), .ZN(n28895) );
  OA22X1 U27157 ( .IN1(n23832), .IN2(n28896), .IN3(n23831), .IN4(n28895), .Q(
        n23809) );
  INVX0 U27158 ( .INP(m0s0_addr[27]), .ZN(n28894) );
  INVX0 U27159 ( .INP(m7s0_addr[27]), .ZN(n28898) );
  OA22X1 U27160 ( .IN1(n23823), .IN2(n28894), .IN3(n23834), .IN4(n28898), .Q(
        n23808) );
  NAND4X0 U27161 ( .IN1(n23811), .IN2(n23810), .IN3(n23809), .IN4(n23808), 
        .QN(s15_addr_o[27]) );
  OA22X1 U27162 ( .IN1(n23812), .IN2(n28908), .IN3(n23818), .IN4(n28911), .Q(
        n23816) );
  OA22X1 U27163 ( .IN1(n23824), .IN2(n28913), .IN3(n23837), .IN4(n28909), .Q(
        n23815) );
  OA22X1 U27164 ( .IN1(n23823), .IN2(n28912), .IN3(n23826), .IN4(n28910), .Q(
        n23814) );
  OA22X1 U27165 ( .IN1(n23836), .IN2(n28906), .IN3(n23833), .IN4(n28907), .Q(
        n23813) );
  NAND4X0 U27166 ( .IN1(n23816), .IN2(n23815), .IN3(n23814), .IN4(n23813), 
        .QN(s15_addr_o[28]) );
  OA22X1 U27167 ( .IN1(n23835), .IN2(n28919), .IN3(n23817), .IN4(n28926), .Q(
        n23822) );
  OA22X1 U27168 ( .IN1(n23838), .IN2(n28925), .IN3(n23833), .IN4(n28922), .Q(
        n23821) );
  OA22X1 U27169 ( .IN1(n23834), .IN2(n28921), .IN3(n23818), .IN4(n28924), .Q(
        n23820) );
  OA22X1 U27170 ( .IN1(n23836), .IN2(n28923), .IN3(n23832), .IN4(n28920), .Q(
        n23819) );
  NAND4X0 U27171 ( .IN1(n23822), .IN2(n23821), .IN3(n23820), .IN4(n23819), 
        .QN(s15_addr_o[29]) );
  OA22X1 U27172 ( .IN1(n23823), .IN2(n28931), .IN3(n23833), .IN4(n28937), .Q(
        n23830) );
  OA22X1 U27173 ( .IN1(n23824), .IN2(n28933), .IN3(n23831), .IN4(n28935), .Q(
        n23829) );
  OA22X1 U27174 ( .IN1(n23825), .IN2(n28939), .IN3(n23837), .IN4(n28932), .Q(
        n23828) );
  OA22X1 U27175 ( .IN1(n23826), .IN2(n28936), .IN3(n23835), .IN4(n28940), .Q(
        n23827) );
  NAND4X0 U27176 ( .IN1(n23830), .IN2(n23829), .IN3(n23828), .IN4(n23827), 
        .QN(s15_addr_o[30]) );
  OA22X1 U27177 ( .IN1(n23832), .IN2(n28954), .IN3(n23831), .IN4(n28952), .Q(
        n23842) );
  OA22X1 U27178 ( .IN1(n23834), .IN2(n28960), .IN3(n23833), .IN4(n28956), .Q(
        n23841) );
  OA22X1 U27179 ( .IN1(n23836), .IN2(n28946), .IN3(n23835), .IN4(n28958), .Q(
        n23840) );
  OA22X1 U27180 ( .IN1(n23838), .IN2(n28950), .IN3(n23837), .IN4(n28948), .Q(
        n23839) );
  NAND4X0 U27181 ( .IN1(n23842), .IN2(n23841), .IN3(n23840), .IN4(n23839), 
        .QN(s15_addr_o[31]) );
  INVX0 U27182 ( .INP(m2_stb_i), .ZN(n29273) );
  INVX0 U27183 ( .INP(m5_stb_i), .ZN(n29330) );
  OA22X1 U27184 ( .IN1(n29273), .IN2(n23844), .IN3(n29330), .IN4(n23843), .Q(
        n23855) );
  AOI22X1 U27185 ( .IN1(m1_stb_i), .IN2(n23846), .IN3(m7_stb_i), .IN4(n23845), 
        .QN(n23854) );
  INVX0 U27186 ( .INP(m0_stb_i), .ZN(n29235) );
  INVX0 U27187 ( .INP(n23847), .ZN(n23849) );
  INVX0 U27188 ( .INP(m4_stb_i), .ZN(n29311) );
  OA22X1 U27189 ( .IN1(n29235), .IN2(n23849), .IN3(n29311), .IN4(n23848), .Q(
        n23853) );
  INVX0 U27190 ( .INP(m6_stb_i), .ZN(n29349) );
  INVX0 U27191 ( .INP(m3_stb_i), .ZN(n29292) );
  OA22X1 U27192 ( .IN1(n29349), .IN2(n23851), .IN3(n29292), .IN4(n23850), .Q(
        n23852) );
  NAND4X0 U27193 ( .IN1(n23855), .IN2(n23854), .IN3(n23853), .IN4(n23852), 
        .QN(s14_stb_o) );
  INVX0 U27194 ( .INP(n29218), .ZN(n24140) );
  INVX0 U27195 ( .INP(n29219), .ZN(n24127) );
  OA22X1 U27196 ( .IN1(n24140), .IN2(n28124), .IN3(n24127), .IN4(n28122), .Q(
        n23859) );
  INVX0 U27197 ( .INP(n29228), .ZN(n24128) );
  OA22X1 U27198 ( .IN1(n24139), .IN2(n28128), .IN3(n24128), .IN4(n28121), .Q(
        n23858) );
  INVX0 U27199 ( .INP(n29225), .ZN(n24138) );
  INVX0 U27200 ( .INP(n29226), .ZN(n24117) );
  OA22X1 U27201 ( .IN1(n24138), .IN2(n28126), .IN3(n24117), .IN4(n28125), .Q(
        n23857) );
  INVX0 U27202 ( .INP(n29217), .ZN(n24130) );
  OA22X1 U27203 ( .IN1(n24130), .IN2(n28123), .IN3(n24096), .IN4(n28127), .Q(
        n23856) );
  NAND4X0 U27204 ( .IN1(n23859), .IN2(n23858), .IN3(n23857), .IN4(n23856), 
        .QN(s14_we_o) );
  INVX0 U27205 ( .INP(n29225), .ZN(n24122) );
  OA22X1 U27206 ( .IN1(n24122), .IN2(n28139), .IN3(n24136), .IN4(n28135), .Q(
        n23863) );
  INVX0 U27207 ( .INP(n29227), .ZN(n24129) );
  OA22X1 U27208 ( .IN1(n24129), .IN2(n28140), .IN3(n24130), .IN4(n28133), .Q(
        n23862) );
  INVX0 U27209 ( .INP(n29219), .ZN(n24142) );
  OA22X1 U27210 ( .IN1(n24142), .IN2(n28138), .IN3(n24096), .IN4(n28137), .Q(
        n23861) );
  OA22X1 U27211 ( .IN1(n24131), .IN2(n28134), .IN3(n24117), .IN4(n28136), .Q(
        n23860) );
  NAND4X0 U27212 ( .IN1(n23863), .IN2(n23862), .IN3(n23861), .IN4(n23860), 
        .QN(s14_data_o[0]) );
  INVX0 U27213 ( .INP(n29226), .ZN(n24141) );
  OA22X1 U27214 ( .IN1(n24141), .IN2(n28152), .IN3(n24096), .IN4(n28151), .Q(
        n23867) );
  OA22X1 U27215 ( .IN1(n24127), .IN2(n28149), .IN3(n24136), .IN4(n28147), .Q(
        n23866) );
  OA22X1 U27216 ( .IN1(n24140), .IN2(n28150), .IN3(n24129), .IN4(n28146), .Q(
        n23865) );
  INVX0 U27217 ( .INP(n29217), .ZN(n24143) );
  OA22X1 U27218 ( .IN1(n24143), .IN2(n28148), .IN3(n24138), .IN4(n28145), .Q(
        n23864) );
  NAND4X0 U27219 ( .IN1(n23867), .IN2(n23866), .IN3(n23865), .IN4(n23864), 
        .QN(s14_data_o[1]) );
  OA22X1 U27220 ( .IN1(n24142), .IN2(n28158), .IN3(n24136), .IN4(n28161), .Q(
        n23871) );
  OA22X1 U27221 ( .IN1(n24141), .IN2(n28162), .IN3(n24096), .IN4(n28157), .Q(
        n23870) );
  OA22X1 U27222 ( .IN1(n24130), .IN2(n28163), .IN3(n24138), .IN4(n28159), .Q(
        n23869) );
  OA22X1 U27223 ( .IN1(n24140), .IN2(n28160), .IN3(n24129), .IN4(n28164), .Q(
        n23868) );
  NAND4X0 U27224 ( .IN1(n23871), .IN2(n23870), .IN3(n23869), .IN4(n23868), 
        .QN(s14_data_o[2]) );
  OA22X1 U27225 ( .IN1(n24140), .IN2(n28172), .IN3(n24127), .IN4(n28171), .Q(
        n23875) );
  OA22X1 U27226 ( .IN1(n24141), .IN2(n28175), .IN3(n24136), .IN4(n28173), .Q(
        n23874) );
  OA22X1 U27227 ( .IN1(n24130), .IN2(n28176), .IN3(n24096), .IN4(n28169), .Q(
        n23873) );
  OA22X1 U27228 ( .IN1(n24139), .IN2(n28174), .IN3(n24138), .IN4(n28170), .Q(
        n23872) );
  NAND4X0 U27229 ( .IN1(n23875), .IN2(n23874), .IN3(n23873), .IN4(n23872), 
        .QN(s14_data_o[3]) );
  OA22X1 U27230 ( .IN1(n24139), .IN2(n28184), .IN3(n24130), .IN4(n28186), .Q(
        n23879) );
  OA22X1 U27231 ( .IN1(n24117), .IN2(n28183), .IN3(n24128), .IN4(n28181), .Q(
        n23878) );
  OA22X1 U27232 ( .IN1(n24140), .IN2(n28182), .IN3(n24138), .IN4(n28188), .Q(
        n23877) );
  OA22X1 U27233 ( .IN1(n24127), .IN2(n28185), .IN3(n24096), .IN4(n28187), .Q(
        n23876) );
  NAND4X0 U27234 ( .IN1(n23879), .IN2(n23878), .IN3(n23877), .IN4(n23876), 
        .QN(s14_data_o[4]) );
  OA22X1 U27235 ( .IN1(n24143), .IN2(n28194), .IN3(n24117), .IN4(n28197), .Q(
        n23883) );
  OA22X1 U27236 ( .IN1(n24138), .IN2(n28193), .IN3(n24127), .IN4(n28198), .Q(
        n23882) );
  OA22X1 U27237 ( .IN1(n24140), .IN2(n28196), .IN3(n24096), .IN4(n28195), .Q(
        n23881) );
  OA22X1 U27238 ( .IN1(n24139), .IN2(n28200), .IN3(n24136), .IN4(n28199), .Q(
        n23880) );
  NAND4X0 U27239 ( .IN1(n23883), .IN2(n23882), .IN3(n23881), .IN4(n23880), 
        .QN(s14_data_o[5]) );
  OA22X1 U27240 ( .IN1(n24130), .IN2(n28206), .IN3(n24128), .IN4(n28209), .Q(
        n23887) );
  OA22X1 U27241 ( .IN1(n24131), .IN2(n28208), .IN3(n24138), .IN4(n28212), .Q(
        n23886) );
  OA22X1 U27242 ( .IN1(n24141), .IN2(n28205), .IN3(n24096), .IN4(n28210), .Q(
        n23885) );
  OA22X1 U27243 ( .IN1(n24139), .IN2(n28207), .IN3(n24127), .IN4(n28211), .Q(
        n23884) );
  NAND4X0 U27244 ( .IN1(n23887), .IN2(n23886), .IN3(n23885), .IN4(n23884), 
        .QN(s14_data_o[6]) );
  OA22X1 U27245 ( .IN1(n24142), .IN2(n28217), .IN3(n24117), .IN4(n28223), .Q(
        n23891) );
  OA22X1 U27246 ( .IN1(n24130), .IN2(n28224), .IN3(n24138), .IN4(n28218), .Q(
        n23890) );
  OA22X1 U27247 ( .IN1(n24139), .IN2(n28219), .IN3(n24136), .IN4(n28221), .Q(
        n23889) );
  OA22X1 U27248 ( .IN1(n24140), .IN2(n28220), .IN3(n24096), .IN4(n28222), .Q(
        n23888) );
  NAND4X0 U27249 ( .IN1(n23891), .IN2(n23890), .IN3(n23889), .IN4(n23888), 
        .QN(s14_data_o[7]) );
  INVX0 U27250 ( .INP(n24096), .ZN(n29220) );
  INVX0 U27251 ( .INP(n29220), .ZN(n24137) );
  OA22X1 U27252 ( .IN1(n24137), .IN2(n28233), .IN3(n24128), .IN4(n28235), .Q(
        n23895) );
  OA22X1 U27253 ( .IN1(n24139), .IN2(n28232), .IN3(n24117), .IN4(n28229), .Q(
        n23894) );
  OA22X1 U27254 ( .IN1(n24131), .IN2(n28230), .IN3(n24138), .IN4(n28234), .Q(
        n23893) );
  OA22X1 U27255 ( .IN1(n24143), .IN2(n28231), .IN3(n24127), .IN4(n28236), .Q(
        n23892) );
  NAND4X0 U27256 ( .IN1(n23895), .IN2(n23894), .IN3(n23893), .IN4(n23892), 
        .QN(s14_data_o[8]) );
  OA22X1 U27257 ( .IN1(n24140), .IN2(n28242), .IN3(n24129), .IN4(n28244), .Q(
        n23899) );
  OA22X1 U27258 ( .IN1(n24127), .IN2(n28241), .IN3(n24117), .IN4(n28245), .Q(
        n23898) );
  OA22X1 U27259 ( .IN1(n24138), .IN2(n28248), .IN3(n24136), .IN4(n28247), .Q(
        n23897) );
  OA22X1 U27260 ( .IN1(n24143), .IN2(n28246), .IN3(n24096), .IN4(n28243), .Q(
        n23896) );
  NAND4X0 U27261 ( .IN1(n23899), .IN2(n23898), .IN3(n23897), .IN4(n23896), 
        .QN(s14_data_o[9]) );
  OA22X1 U27262 ( .IN1(n24131), .IN2(n28258), .IN3(n24130), .IN4(n28260), .Q(
        n23903) );
  OA22X1 U27263 ( .IN1(n24139), .IN2(n28257), .IN3(n24138), .IN4(n28256), .Q(
        n23902) );
  OA22X1 U27264 ( .IN1(n24137), .IN2(n28253), .IN3(n24128), .IN4(n28259), .Q(
        n23901) );
  OA22X1 U27265 ( .IN1(n24142), .IN2(n28254), .IN3(n24117), .IN4(n28255), .Q(
        n23900) );
  NAND4X0 U27266 ( .IN1(n23903), .IN2(n23902), .IN3(n23901), .IN4(n23900), 
        .QN(s14_data_o[10]) );
  OA22X1 U27267 ( .IN1(n24140), .IN2(n28266), .IN3(n24117), .IN4(n28270), .Q(
        n23907) );
  OA22X1 U27268 ( .IN1(n24127), .IN2(n28268), .IN3(n24136), .IN4(n28269), .Q(
        n23906) );
  OA22X1 U27269 ( .IN1(n24139), .IN2(n28272), .IN3(n24138), .IN4(n28271), .Q(
        n23905) );
  OA22X1 U27270 ( .IN1(n24130), .IN2(n28265), .IN3(n24137), .IN4(n28267), .Q(
        n23904) );
  NAND4X0 U27271 ( .IN1(n23907), .IN2(n23906), .IN3(n23905), .IN4(n23904), 
        .QN(s14_data_o[11]) );
  OA22X1 U27272 ( .IN1(n24139), .IN2(n28278), .IN3(n24128), .IN4(n28277), .Q(
        n23911) );
  OA22X1 U27273 ( .IN1(n24131), .IN2(n28284), .IN3(n24138), .IN4(n28282), .Q(
        n23910) );
  OA22X1 U27274 ( .IN1(n24142), .IN2(n28283), .IN3(n24117), .IN4(n28281), .Q(
        n23909) );
  OA22X1 U27275 ( .IN1(n24143), .IN2(n28280), .IN3(n24137), .IN4(n28279), .Q(
        n23908) );
  NAND4X0 U27276 ( .IN1(n23911), .IN2(n23910), .IN3(n23909), .IN4(n23908), 
        .QN(s14_data_o[12]) );
  OA22X1 U27277 ( .IN1(n24139), .IN2(n28294), .IN3(n24130), .IN4(n28296), .Q(
        n23915) );
  OA22X1 U27278 ( .IN1(n24127), .IN2(n28289), .IN3(n24137), .IN4(n28291), .Q(
        n23914) );
  OA22X1 U27279 ( .IN1(n24140), .IN2(n28290), .IN3(n24136), .IN4(n28295), .Q(
        n23913) );
  OA22X1 U27280 ( .IN1(n24122), .IN2(n28292), .IN3(n24117), .IN4(n28293), .Q(
        n23912) );
  NAND4X0 U27281 ( .IN1(n23915), .IN2(n23914), .IN3(n23913), .IN4(n23912), 
        .QN(s14_data_o[13]) );
  OA22X1 U27282 ( .IN1(n24131), .IN2(n28306), .IN3(n24129), .IN4(n28304), .Q(
        n23919) );
  OA22X1 U27283 ( .IN1(n24130), .IN2(n28308), .IN3(n24141), .IN4(n28302), .Q(
        n23918) );
  OA22X1 U27284 ( .IN1(n24122), .IN2(n28305), .IN3(n24127), .IN4(n28307), .Q(
        n23917) );
  OA22X1 U27285 ( .IN1(n24096), .IN2(n28301), .IN3(n24128), .IN4(n28303), .Q(
        n23916) );
  NAND4X0 U27286 ( .IN1(n23919), .IN2(n23918), .IN3(n23917), .IN4(n23916), 
        .QN(s14_data_o[14]) );
  OA22X1 U27287 ( .IN1(n24130), .IN2(n28314), .IN3(n24127), .IN4(n28320), .Q(
        n23923) );
  OA22X1 U27288 ( .IN1(n24139), .IN2(n28315), .IN3(n24117), .IN4(n28318), .Q(
        n23922) );
  OA22X1 U27289 ( .IN1(n24140), .IN2(n28316), .IN3(n24137), .IN4(n28317), .Q(
        n23921) );
  OA22X1 U27290 ( .IN1(n24138), .IN2(n28313), .IN3(n24136), .IN4(n28319), .Q(
        n23920) );
  NAND4X0 U27291 ( .IN1(n23923), .IN2(n23922), .IN3(n23921), .IN4(n23920), 
        .QN(s14_data_o[15]) );
  OA22X1 U27292 ( .IN1(n24131), .IN2(n28330), .IN3(n24127), .IN4(n28329), .Q(
        n23927) );
  OA22X1 U27293 ( .IN1(n24129), .IN2(n28332), .IN3(n24130), .IN4(n28331), .Q(
        n23926) );
  OA22X1 U27294 ( .IN1(n24122), .IN2(n28326), .IN3(n24141), .IN4(n28325), .Q(
        n23925) );
  OA22X1 U27295 ( .IN1(n24096), .IN2(n28328), .IN3(n24128), .IN4(n28327), .Q(
        n23924) );
  NAND4X0 U27296 ( .IN1(n23927), .IN2(n23926), .IN3(n23925), .IN4(n23924), 
        .QN(s14_data_o[16]) );
  OA22X1 U27297 ( .IN1(n24140), .IN2(n28340), .IN3(n24141), .IN4(n28339), .Q(
        n23931) );
  OA22X1 U27298 ( .IN1(n24139), .IN2(n28344), .IN3(n24130), .IN4(n28342), .Q(
        n23930) );
  OA22X1 U27299 ( .IN1(n24122), .IN2(n28338), .IN3(n24142), .IN4(n28337), .Q(
        n23929) );
  OA22X1 U27300 ( .IN1(n24096), .IN2(n28343), .IN3(n24136), .IN4(n28341), .Q(
        n23928) );
  NAND4X0 U27301 ( .IN1(n23931), .IN2(n23930), .IN3(n23929), .IN4(n23928), 
        .QN(s14_data_o[17]) );
  OA22X1 U27302 ( .IN1(n24142), .IN2(n28354), .IN3(n24128), .IN4(n28353), .Q(
        n23935) );
  OA22X1 U27303 ( .IN1(n24143), .IN2(n28350), .IN3(n24117), .IN4(n28349), .Q(
        n23934) );
  OA22X1 U27304 ( .IN1(n24139), .IN2(n28356), .IN3(n24138), .IN4(n28355), .Q(
        n23933) );
  OA22X1 U27305 ( .IN1(n24131), .IN2(n28352), .IN3(n24137), .IN4(n28351), .Q(
        n23932) );
  NAND4X0 U27306 ( .IN1(n23935), .IN2(n23934), .IN3(n23933), .IN4(n23932), 
        .QN(s14_data_o[18]) );
  OA22X1 U27307 ( .IN1(n24131), .IN2(n28366), .IN3(n24136), .IN4(n28367), .Q(
        n23939) );
  OA22X1 U27308 ( .IN1(n24141), .IN2(n28361), .IN3(n24137), .IN4(n28368), .Q(
        n23938) );
  OA22X1 U27309 ( .IN1(n24129), .IN2(n28364), .IN3(n24130), .IN4(n28362), .Q(
        n23937) );
  OA22X1 U27310 ( .IN1(n24138), .IN2(n28363), .IN3(n24127), .IN4(n28365), .Q(
        n23936) );
  NAND4X0 U27311 ( .IN1(n23939), .IN2(n23938), .IN3(n23937), .IN4(n23936), 
        .QN(s14_data_o[19]) );
  OA22X1 U27312 ( .IN1(n24143), .IN2(n28374), .IN3(n24142), .IN4(n28376), .Q(
        n23943) );
  OA22X1 U27313 ( .IN1(n24138), .IN2(n28373), .IN3(n24137), .IN4(n28379), .Q(
        n23942) );
  OA22X1 U27314 ( .IN1(n24141), .IN2(n28380), .IN3(n24128), .IN4(n28375), .Q(
        n23941) );
  OA22X1 U27315 ( .IN1(n24131), .IN2(n28378), .IN3(n24129), .IN4(n28377), .Q(
        n23940) );
  NAND4X0 U27316 ( .IN1(n23943), .IN2(n23942), .IN3(n23941), .IN4(n23940), 
        .QN(s14_data_o[20]) );
  OA22X1 U27317 ( .IN1(n24131), .IN2(n28392), .IN3(n24137), .IN4(n28389), .Q(
        n23947) );
  OA22X1 U27318 ( .IN1(n24130), .IN2(n28390), .IN3(n24138), .IN4(n28388), .Q(
        n23946) );
  OA22X1 U27319 ( .IN1(n24127), .IN2(n28387), .IN3(n24128), .IN4(n28391), .Q(
        n23945) );
  OA22X1 U27320 ( .IN1(n24139), .IN2(n28386), .IN3(n24117), .IN4(n28385), .Q(
        n23944) );
  NAND4X0 U27321 ( .IN1(n23947), .IN2(n23946), .IN3(n23945), .IN4(n23944), 
        .QN(s14_data_o[21]) );
  OA22X1 U27322 ( .IN1(n24129), .IN2(n28402), .IN3(n24141), .IN4(n28399), .Q(
        n23951) );
  OA22X1 U27323 ( .IN1(n24137), .IN2(n28401), .IN3(n24128), .IN4(n28397), .Q(
        n23950) );
  OA22X1 U27324 ( .IN1(n24131), .IN2(n28400), .IN3(n24142), .IN4(n28398), .Q(
        n23949) );
  OA22X1 U27325 ( .IN1(n24143), .IN2(n28404), .IN3(n24138), .IN4(n28403), .Q(
        n23948) );
  NAND4X0 U27326 ( .IN1(n23951), .IN2(n23950), .IN3(n23949), .IN4(n23948), 
        .QN(s14_data_o[22]) );
  OA22X1 U27327 ( .IN1(n24122), .IN2(n28413), .IN3(n24117), .IN4(n28412), .Q(
        n23955) );
  OA22X1 U27328 ( .IN1(n24096), .IN2(n28409), .IN3(n24128), .IN4(n28411), .Q(
        n23954) );
  OA22X1 U27329 ( .IN1(n24139), .IN2(n28415), .IN3(n24127), .IN4(n28410), .Q(
        n23953) );
  OA22X1 U27330 ( .IN1(n24131), .IN2(n28416), .IN3(n24130), .IN4(n28414), .Q(
        n23952) );
  NAND4X0 U27331 ( .IN1(n23955), .IN2(n23954), .IN3(n23953), .IN4(n23952), 
        .QN(s14_data_o[23]) );
  OA22X1 U27332 ( .IN1(n24131), .IN2(n28426), .IN3(n24137), .IN4(n28427), .Q(
        n23959) );
  OA22X1 U27333 ( .IN1(n24141), .IN2(n28428), .IN3(n24128), .IN4(n28423), .Q(
        n23958) );
  OA22X1 U27334 ( .IN1(n24129), .IN2(n28424), .IN3(n24138), .IN4(n28421), .Q(
        n23957) );
  OA22X1 U27335 ( .IN1(n24130), .IN2(n28422), .IN3(n24127), .IN4(n28425), .Q(
        n23956) );
  NAND4X0 U27336 ( .IN1(n23959), .IN2(n23958), .IN3(n23957), .IN4(n23956), 
        .QN(s14_data_o[24]) );
  OA22X1 U27337 ( .IN1(n24138), .IN2(n28439), .IN3(n24128), .IN4(n28435), .Q(
        n23963) );
  OA22X1 U27338 ( .IN1(n24131), .IN2(n28438), .IN3(n24130), .IN4(n28434), .Q(
        n23962) );
  OA22X1 U27339 ( .IN1(n24139), .IN2(n28440), .IN3(n24141), .IN4(n28437), .Q(
        n23961) );
  OA22X1 U27340 ( .IN1(n24142), .IN2(n28433), .IN3(n24137), .IN4(n28436), .Q(
        n23960) );
  NAND4X0 U27341 ( .IN1(n23963), .IN2(n23962), .IN3(n23961), .IN4(n23960), 
        .QN(s14_data_o[25]) );
  OA22X1 U27342 ( .IN1(n24131), .IN2(n28452), .IN3(n24122), .IN4(n28446), .Q(
        n23967) );
  OA22X1 U27343 ( .IN1(n24129), .IN2(n28451), .IN3(n24130), .IN4(n28450), .Q(
        n23966) );
  OA22X1 U27344 ( .IN1(n24142), .IN2(n28449), .IN3(n24141), .IN4(n28448), .Q(
        n23965) );
  OA22X1 U27345 ( .IN1(n24096), .IN2(n28447), .IN3(n24128), .IN4(n28445), .Q(
        n23964) );
  NAND4X0 U27346 ( .IN1(n23967), .IN2(n23966), .IN3(n23965), .IN4(n23964), 
        .QN(s14_data_o[26]) );
  OA22X1 U27347 ( .IN1(n24131), .IN2(n28462), .IN3(n24127), .IN4(n28457), .Q(
        n23971) );
  OA22X1 U27348 ( .IN1(n24122), .IN2(n28458), .IN3(n24128), .IN4(n28459), .Q(
        n23970) );
  OA22X1 U27349 ( .IN1(n24139), .IN2(n28461), .IN3(n24117), .IN4(n28463), .Q(
        n23969) );
  OA22X1 U27350 ( .IN1(n24130), .IN2(n28464), .IN3(n24137), .IN4(n28460), .Q(
        n23968) );
  NAND4X0 U27351 ( .IN1(n23971), .IN2(n23970), .IN3(n23969), .IN4(n23968), 
        .QN(s14_data_o[27]) );
  OA22X1 U27352 ( .IN1(n24131), .IN2(n28474), .IN3(n24129), .IN4(n28476), .Q(
        n23975) );
  OA22X1 U27353 ( .IN1(n24138), .IN2(n28470), .IN3(n24117), .IN4(n28475), .Q(
        n23974) );
  OA22X1 U27354 ( .IN1(n24143), .IN2(n28472), .IN3(n24128), .IN4(n28473), .Q(
        n23973) );
  OA22X1 U27355 ( .IN1(n24142), .IN2(n28471), .IN3(n24137), .IN4(n28469), .Q(
        n23972) );
  NAND4X0 U27356 ( .IN1(n23975), .IN2(n23974), .IN3(n23973), .IN4(n23972), 
        .QN(s14_data_o[28]) );
  OA22X1 U27357 ( .IN1(n24122), .IN2(n28486), .IN3(n24127), .IN4(n28487), .Q(
        n23979) );
  OA22X1 U27358 ( .IN1(n24131), .IN2(n28484), .IN3(n24129), .IN4(n28482), .Q(
        n23978) );
  OA22X1 U27359 ( .IN1(n24117), .IN2(n28483), .IN3(n24137), .IN4(n28485), .Q(
        n23977) );
  OA22X1 U27360 ( .IN1(n24143), .IN2(n28488), .IN3(n24128), .IN4(n28481), .Q(
        n23976) );
  NAND4X0 U27361 ( .IN1(n23979), .IN2(n23978), .IN3(n23977), .IN4(n23976), 
        .QN(s14_data_o[29]) );
  OA22X1 U27362 ( .IN1(n24142), .IN2(n28493), .IN3(n24141), .IN4(n28495), .Q(
        n23983) );
  OA22X1 U27363 ( .IN1(n24129), .IN2(n28498), .IN3(n24128), .IN4(n28499), .Q(
        n23982) );
  OA22X1 U27364 ( .IN1(n24130), .IN2(n28497), .IN3(n24138), .IN4(n28496), .Q(
        n23981) );
  OA22X1 U27365 ( .IN1(n24131), .IN2(n28494), .IN3(n24137), .IN4(n28500), .Q(
        n23980) );
  NAND4X0 U27366 ( .IN1(n23983), .IN2(n23982), .IN3(n23981), .IN4(n23980), 
        .QN(s14_data_o[30]) );
  OA22X1 U27367 ( .IN1(n24131), .IN2(n28510), .IN3(n24129), .IN4(n28509), .Q(
        n23987) );
  OA22X1 U27368 ( .IN1(n24142), .IN2(n28512), .IN3(n24117), .IN4(n28508), .Q(
        n23986) );
  OA22X1 U27369 ( .IN1(n24138), .IN2(n28505), .IN3(n24128), .IN4(n28507), .Q(
        n23985) );
  OA22X1 U27370 ( .IN1(n24130), .IN2(n28506), .IN3(n24137), .IN4(n28511), .Q(
        n23984) );
  NAND4X0 U27371 ( .IN1(n23987), .IN2(n23986), .IN3(n23985), .IN4(n23984), 
        .QN(s14_data_o[31]) );
  OA22X1 U27372 ( .IN1(n24122), .IN2(n28524), .IN3(n24137), .IN4(n28521), .Q(
        n23991) );
  OA22X1 U27373 ( .IN1(n24131), .IN2(n28518), .IN3(n24127), .IN4(n28523), .Q(
        n23990) );
  OA22X1 U27374 ( .IN1(n24130), .IN2(n28522), .IN3(n24141), .IN4(n28520), .Q(
        n23989) );
  OA22X1 U27375 ( .IN1(n24139), .IN2(n28517), .IN3(n24128), .IN4(n28519), .Q(
        n23988) );
  NAND4X0 U27376 ( .IN1(n23991), .IN2(n23990), .IN3(n23989), .IN4(n23988), 
        .QN(s14_sel_o[0]) );
  OA22X1 U27377 ( .IN1(n24143), .IN2(n28530), .IN3(n24142), .IN4(n28535), .Q(
        n23995) );
  OA22X1 U27378 ( .IN1(n24129), .IN2(n28532), .IN3(n24122), .IN4(n28536), .Q(
        n23994) );
  OA22X1 U27379 ( .IN1(n24140), .IN2(n28534), .IN3(n24128), .IN4(n28529), .Q(
        n23993) );
  OA22X1 U27380 ( .IN1(n24141), .IN2(n28533), .IN3(n24096), .IN4(n28531), .Q(
        n23992) );
  NAND4X0 U27381 ( .IN1(n23995), .IN2(n23994), .IN3(n23993), .IN4(n23992), 
        .QN(s14_sel_o[1]) );
  OA22X1 U27382 ( .IN1(n24129), .IN2(n28546), .IN3(n24096), .IN4(n28545), .Q(
        n23999) );
  OA22X1 U27383 ( .IN1(n24138), .IN2(n28548), .IN3(n24142), .IN4(n28547), .Q(
        n23998) );
  OA22X1 U27384 ( .IN1(n24140), .IN2(n28544), .IN3(n24130), .IN4(n28543), .Q(
        n23997) );
  OA22X1 U27385 ( .IN1(n24117), .IN2(n28542), .IN3(n24128), .IN4(n28541), .Q(
        n23996) );
  NAND4X0 U27386 ( .IN1(n23999), .IN2(n23998), .IN3(n23997), .IN4(n23996), 
        .QN(s14_sel_o[2]) );
  OA22X1 U27387 ( .IN1(n24143), .IN2(n28553), .IN3(n24128), .IN4(n28555), .Q(
        n24003) );
  OA22X1 U27388 ( .IN1(n24122), .IN2(n28557), .IN3(n24141), .IN4(n28560), .Q(
        n24002) );
  OA22X1 U27389 ( .IN1(n24140), .IN2(n28558), .IN3(n24096), .IN4(n28559), .Q(
        n24001) );
  OA22X1 U27390 ( .IN1(n24129), .IN2(n28554), .IN3(n24127), .IN4(n28556), .Q(
        n24000) );
  NAND4X0 U27391 ( .IN1(n24003), .IN2(n24002), .IN3(n24001), .IN4(n24000), 
        .QN(s14_sel_o[3]) );
  OA22X1 U27392 ( .IN1(n24129), .IN2(n28570), .IN3(n24128), .IN4(n28569), .Q(
        n24007) );
  OA22X1 U27393 ( .IN1(n24142), .IN2(n28568), .IN3(n24117), .IN4(n28567), .Q(
        n24006) );
  OA22X1 U27394 ( .IN1(n24143), .IN2(n28571), .IN3(n24096), .IN4(n28565), .Q(
        n24005) );
  OA22X1 U27395 ( .IN1(n24140), .IN2(n28572), .IN3(n24122), .IN4(n28566), .Q(
        n24004) );
  NAND4X0 U27396 ( .IN1(n24007), .IN2(n24006), .IN3(n24005), .IN4(n24004), 
        .QN(s14_addr_o[0]) );
  OA22X1 U27397 ( .IN1(n24129), .IN2(n28578), .IN3(n24127), .IN4(n28579), .Q(
        n24011) );
  OA22X1 U27398 ( .IN1(n24143), .IN2(n28582), .IN3(n24122), .IN4(n28581), .Q(
        n24010) );
  OA22X1 U27399 ( .IN1(n24140), .IN2(n28580), .IN3(n24136), .IN4(n28583), .Q(
        n24009) );
  OA22X1 U27400 ( .IN1(n24141), .IN2(n28584), .IN3(n24096), .IN4(n28577), .Q(
        n24008) );
  NAND4X0 U27401 ( .IN1(n24011), .IN2(n24010), .IN3(n24009), .IN4(n24008), 
        .QN(s14_addr_o[1]) );
  OA22X1 U27402 ( .IN1(n28592), .IN2(n24122), .IN3(n28593), .IN4(n24141), .Q(
        n24015) );
  OA22X1 U27403 ( .IN1(n28591), .IN2(n24140), .IN3(n28590), .IN4(n24127), .Q(
        n24014) );
  OA22X1 U27404 ( .IN1(n28589), .IN2(n24139), .IN3(n28595), .IN4(n24096), .Q(
        n24013) );
  OA22X1 U27405 ( .IN1(n28596), .IN2(n24128), .IN3(n28594), .IN4(n24143), .Q(
        n24012) );
  NAND4X0 U27406 ( .IN1(n24015), .IN2(n24014), .IN3(n24013), .IN4(n24012), 
        .QN(s14_addr_o[2]) );
  OA22X1 U27407 ( .IN1(n28601), .IN2(n24131), .IN3(n28603), .IN4(n24096), .Q(
        n24019) );
  OA22X1 U27408 ( .IN1(n28602), .IN2(n24141), .IN3(n28608), .IN4(n24136), .Q(
        n24018) );
  OA22X1 U27409 ( .IN1(n28604), .IN2(n24130), .IN3(n28605), .IN4(n24139), .Q(
        n24017) );
  OA22X1 U27410 ( .IN1(n28606), .IN2(n24127), .IN3(n28607), .IN4(n24138), .Q(
        n24016) );
  NAND4X0 U27411 ( .IN1(n24019), .IN2(n24018), .IN3(n24017), .IN4(n24016), 
        .QN(s14_addr_o[3]) );
  OA22X1 U27412 ( .IN1(n28616), .IN2(n24129), .IN3(n28614), .IN4(n24117), .Q(
        n24023) );
  OA22X1 U27413 ( .IN1(n28617), .IN2(n24140), .IN3(n28613), .IN4(n24143), .Q(
        n24022) );
  OA22X1 U27414 ( .IN1(n28620), .IN2(n24137), .IN3(n28619), .IN4(n24136), .Q(
        n24021) );
  OA22X1 U27415 ( .IN1(n28618), .IN2(n24122), .IN3(n28615), .IN4(n24127), .Q(
        n24020) );
  NAND4X0 U27416 ( .IN1(n24023), .IN2(n24022), .IN3(n24021), .IN4(n24020), 
        .QN(s14_addr_o[4]) );
  OA22X1 U27417 ( .IN1(n28625), .IN2(n24136), .IN3(n28629), .IN4(n24140), .Q(
        n24027) );
  OA22X1 U27418 ( .IN1(n28626), .IN2(n24122), .IN3(n28631), .IN4(n24127), .Q(
        n24026) );
  OA22X1 U27419 ( .IN1(n28632), .IN2(n24143), .IN3(n28630), .IN4(n24139), .Q(
        n24025) );
  OA22X1 U27420 ( .IN1(n28628), .IN2(n24137), .IN3(n28627), .IN4(n24141), .Q(
        n24024) );
  NAND4X0 U27421 ( .IN1(n24027), .IN2(n24026), .IN3(n24025), .IN4(n24024), 
        .QN(s14_addr_o[5]) );
  OA22X1 U27422 ( .IN1(n24143), .IN2(n28644), .IN3(n24117), .IN4(n28637), .Q(
        n24031) );
  OA22X1 U27423 ( .IN1(n24131), .IN2(n28642), .IN3(n24142), .IN4(n28638), .Q(
        n24030) );
  OA22X1 U27424 ( .IN1(n24139), .IN2(n28640), .IN3(n24138), .IN4(n28643), .Q(
        n24029) );
  OA22X1 U27425 ( .IN1(n24096), .IN2(n28641), .IN3(n24136), .IN4(n28639), .Q(
        n24028) );
  NAND4X0 U27426 ( .IN1(n24031), .IN2(n24030), .IN3(n24029), .IN4(n24028), 
        .QN(s14_addr_o[6]) );
  OA22X1 U27427 ( .IN1(n24138), .IN2(n28653), .IN3(n24117), .IN4(n28649), .Q(
        n24035) );
  OA22X1 U27428 ( .IN1(n24142), .IN2(n28650), .IN3(n24136), .IN4(n28655), .Q(
        n24034) );
  OA22X1 U27429 ( .IN1(n24131), .IN2(n28654), .IN3(n24096), .IN4(n28651), .Q(
        n24033) );
  OA22X1 U27430 ( .IN1(n24129), .IN2(n28652), .IN3(n24130), .IN4(n28656), .Q(
        n24032) );
  NAND4X0 U27431 ( .IN1(n24035), .IN2(n24034), .IN3(n24033), .IN4(n24032), 
        .QN(s14_addr_o[7]) );
  OA22X1 U27432 ( .IN1(n24140), .IN2(n28664), .IN3(n24142), .IN4(n28668), .Q(
        n24039) );
  OA22X1 U27433 ( .IN1(n24139), .IN2(n28663), .IN3(n24117), .IN4(n28662), .Q(
        n24038) );
  OA22X1 U27434 ( .IN1(n24143), .IN2(n28666), .IN3(n24138), .IN4(n28665), .Q(
        n24037) );
  OA22X1 U27435 ( .IN1(n24096), .IN2(n28661), .IN3(n24136), .IN4(n28667), .Q(
        n24036) );
  NAND4X0 U27436 ( .IN1(n24039), .IN2(n24038), .IN3(n24037), .IN4(n24036), 
        .QN(s14_addr_o[8]) );
  OA22X1 U27437 ( .IN1(n24143), .IN2(n28674), .IN3(n24136), .IN4(n28677), .Q(
        n24043) );
  OA22X1 U27438 ( .IN1(n24142), .IN2(n28673), .IN3(n24117), .IN4(n28678), .Q(
        n24042) );
  OA22X1 U27439 ( .IN1(n24140), .IN2(n28680), .IN3(n24122), .IN4(n28676), .Q(
        n24041) );
  OA22X1 U27440 ( .IN1(n24129), .IN2(n28679), .IN3(n24096), .IN4(n28675), .Q(
        n24040) );
  NAND4X0 U27441 ( .IN1(n24043), .IN2(n24042), .IN3(n24041), .IN4(n24040), 
        .QN(s14_addr_o[9]) );
  OA22X1 U27442 ( .IN1(n24140), .IN2(n28692), .IN3(n24136), .IN4(n28689), .Q(
        n24047) );
  OA22X1 U27443 ( .IN1(n24139), .IN2(n28686), .IN3(n24096), .IN4(n28690), .Q(
        n24046) );
  OA22X1 U27444 ( .IN1(n24143), .IN2(n28688), .IN3(n24122), .IN4(n28687), .Q(
        n24045) );
  OA22X1 U27445 ( .IN1(n24142), .IN2(n28685), .IN3(n24117), .IN4(n28691), .Q(
        n24044) );
  NAND4X0 U27446 ( .IN1(n24047), .IN2(n24046), .IN3(n24045), .IN4(n24044), 
        .QN(s14_addr_o[10]) );
  OA22X1 U27447 ( .IN1(n24129), .IN2(n28698), .IN3(n24096), .IN4(n28700), .Q(
        n24051) );
  OA22X1 U27448 ( .IN1(n24143), .IN2(n28697), .IN3(n24117), .IN4(n28703), .Q(
        n24050) );
  OA22X1 U27449 ( .IN1(n24131), .IN2(n28702), .IN3(n24136), .IN4(n28699), .Q(
        n24049) );
  OA22X1 U27450 ( .IN1(n24122), .IN2(n28704), .IN3(n24127), .IN4(n28701), .Q(
        n24048) );
  NAND4X0 U27451 ( .IN1(n24051), .IN2(n24050), .IN3(n24049), .IN4(n24048), 
        .QN(s14_addr_o[11]) );
  OA22X1 U27452 ( .IN1(n24129), .IN2(n28710), .IN3(n24136), .IN4(n28713), .Q(
        n24055) );
  OA22X1 U27453 ( .IN1(n24131), .IN2(n28714), .IN3(n24141), .IN4(n28715), .Q(
        n24054) );
  OA22X1 U27454 ( .IN1(n24143), .IN2(n28712), .IN3(n24096), .IN4(n28711), .Q(
        n24053) );
  OA22X1 U27455 ( .IN1(n24122), .IN2(n28716), .IN3(n24142), .IN4(n28709), .Q(
        n24052) );
  NAND4X0 U27456 ( .IN1(n24055), .IN2(n24054), .IN3(n24053), .IN4(n24052), 
        .QN(s14_addr_o[12]) );
  OA22X1 U27457 ( .IN1(n24140), .IN2(n28722), .IN3(n24117), .IN4(n28721), .Q(
        n24059) );
  OA22X1 U27458 ( .IN1(n24143), .IN2(n28726), .IN3(n24142), .IN4(n28723), .Q(
        n24058) );
  OA22X1 U27459 ( .IN1(n24129), .IN2(n28728), .IN3(n24138), .IN4(n28724), .Q(
        n24057) );
  OA22X1 U27460 ( .IN1(n24096), .IN2(n28725), .IN3(n24136), .IN4(n28727), .Q(
        n24056) );
  NAND4X0 U27461 ( .IN1(n24059), .IN2(n24058), .IN3(n24057), .IN4(n24056), 
        .QN(s14_addr_o[13]) );
  OA22X1 U27462 ( .IN1(n24140), .IN2(n28734), .IN3(n24127), .IN4(n28740), .Q(
        n24063) );
  OA22X1 U27463 ( .IN1(n24117), .IN2(n28737), .IN3(n24136), .IN4(n28739), .Q(
        n24062) );
  OA22X1 U27464 ( .IN1(n24139), .IN2(n28738), .IN3(n24096), .IN4(n28733), .Q(
        n24061) );
  OA22X1 U27465 ( .IN1(n24143), .IN2(n28736), .IN3(n24138), .IN4(n28735), .Q(
        n24060) );
  NAND4X0 U27466 ( .IN1(n24063), .IN2(n24062), .IN3(n24061), .IN4(n24060), 
        .QN(s14_addr_o[14]) );
  OA22X1 U27467 ( .IN1(n24129), .IN2(n28748), .IN3(n24117), .IN4(n28751), .Q(
        n24067) );
  OA22X1 U27468 ( .IN1(n24130), .IN2(n28750), .IN3(n24128), .IN4(n28745), .Q(
        n24066) );
  OA22X1 U27469 ( .IN1(n24142), .IN2(n28747), .IN3(n24096), .IN4(n28749), .Q(
        n24065) );
  OA22X1 U27470 ( .IN1(n24131), .IN2(n28746), .IN3(n24138), .IN4(n28752), .Q(
        n24064) );
  NAND4X0 U27471 ( .IN1(n24067), .IN2(n24066), .IN3(n24065), .IN4(n24064), 
        .QN(s14_addr_o[15]) );
  OA22X1 U27472 ( .IN1(n24143), .IN2(n28760), .IN3(n24136), .IN4(n28763), .Q(
        n24071) );
  OA22X1 U27473 ( .IN1(n24139), .IN2(n28762), .IN3(n24117), .IN4(n28757), .Q(
        n24070) );
  OA22X1 U27474 ( .IN1(n24122), .IN2(n28761), .IN3(n24096), .IN4(n28764), .Q(
        n24069) );
  OA22X1 U27475 ( .IN1(n24131), .IN2(n28758), .IN3(n24127), .IN4(n28759), .Q(
        n24068) );
  NAND4X0 U27476 ( .IN1(n24071), .IN2(n24070), .IN3(n24069), .IN4(n24068), 
        .QN(s14_addr_o[16]) );
  OA22X1 U27477 ( .IN1(n24122), .IN2(n28773), .IN3(n24136), .IN4(n28769), .Q(
        n24075) );
  OA22X1 U27478 ( .IN1(n24131), .IN2(n28772), .IN3(n24130), .IN4(n28774), .Q(
        n24074) );
  OA22X1 U27479 ( .IN1(n24129), .IN2(n28776), .IN3(n24141), .IN4(n28771), .Q(
        n24073) );
  OA22X1 U27480 ( .IN1(n24142), .IN2(n28775), .IN3(n24096), .IN4(n28770), .Q(
        n24072) );
  NAND4X0 U27481 ( .IN1(n24075), .IN2(n24074), .IN3(n24073), .IN4(n24072), 
        .QN(s14_addr_o[17]) );
  OA22X1 U27482 ( .IN1(n24143), .IN2(n28787), .IN3(n24138), .IN4(n28782), .Q(
        n24079) );
  OA22X1 U27483 ( .IN1(n24129), .IN2(n28788), .IN3(n24117), .IN4(n28783), .Q(
        n24078) );
  OA22X1 U27484 ( .IN1(n24142), .IN2(n28784), .IN3(n24136), .IN4(n28781), .Q(
        n24077) );
  OA22X1 U27485 ( .IN1(n24131), .IN2(n28786), .IN3(n24096), .IN4(n28785), .Q(
        n24076) );
  NAND4X0 U27486 ( .IN1(n24079), .IN2(n24078), .IN3(n24077), .IN4(n24076), 
        .QN(s14_addr_o[18]) );
  OA22X1 U27487 ( .IN1(n24131), .IN2(n28796), .IN3(n24136), .IN4(n28799), .Q(
        n24083) );
  OA22X1 U27488 ( .IN1(n24122), .IN2(n28794), .IN3(n24142), .IN4(n28797), .Q(
        n24082) );
  OA22X1 U27489 ( .IN1(n24129), .IN2(n28800), .IN3(n24130), .IN4(n28798), .Q(
        n24081) );
  OA22X1 U27490 ( .IN1(n24141), .IN2(n28795), .IN3(n24096), .IN4(n28793), .Q(
        n24080) );
  NAND4X0 U27491 ( .IN1(n24083), .IN2(n24082), .IN3(n24081), .IN4(n24080), 
        .QN(s14_addr_o[19]) );
  OA22X1 U27492 ( .IN1(n24122), .IN2(n28810), .IN3(n24127), .IN4(n28806), .Q(
        n24087) );
  OA22X1 U27493 ( .IN1(n24143), .IN2(n28807), .IN3(n24096), .IN4(n28809), .Q(
        n24086) );
  OA22X1 U27494 ( .IN1(n24141), .IN2(n28811), .IN3(n24128), .IN4(n28805), .Q(
        n24085) );
  OA22X1 U27495 ( .IN1(n24140), .IN2(n28812), .IN3(n24129), .IN4(n28808), .Q(
        n24084) );
  NAND4X0 U27496 ( .IN1(n24087), .IN2(n24086), .IN3(n24085), .IN4(n24084), 
        .QN(s14_addr_o[20]) );
  OA22X1 U27497 ( .IN1(n24131), .IN2(n28822), .IN3(n24096), .IN4(n28818), .Q(
        n24091) );
  OA22X1 U27498 ( .IN1(n24122), .IN2(n28819), .IN3(n24141), .IN4(n28823), .Q(
        n24090) );
  OA22X1 U27499 ( .IN1(n24139), .IN2(n28824), .IN3(n24142), .IN4(n28821), .Q(
        n24089) );
  OA22X1 U27500 ( .IN1(n24143), .IN2(n28820), .IN3(n24128), .IN4(n28817), .Q(
        n24088) );
  NAND4X0 U27501 ( .IN1(n24091), .IN2(n24090), .IN3(n24089), .IN4(n24088), 
        .QN(s14_addr_o[21]) );
  OA22X1 U27502 ( .IN1(n24140), .IN2(n28833), .IN3(n24096), .IN4(n28837), .Q(
        n24095) );
  OA22X1 U27503 ( .IN1(n24129), .IN2(n28832), .IN3(n24117), .IN4(n28834), .Q(
        n24094) );
  OA22X1 U27504 ( .IN1(n24130), .IN2(n28831), .IN3(n24136), .IN4(n28829), .Q(
        n24093) );
  OA22X1 U27505 ( .IN1(n24122), .IN2(n28838), .IN3(n24142), .IN4(n28836), .Q(
        n24092) );
  NAND4X0 U27506 ( .IN1(n24095), .IN2(n24094), .IN3(n24093), .IN4(n24092), 
        .QN(s14_addr_o[22]) );
  OA22X1 U27507 ( .IN1(n24122), .IN2(n28850), .IN3(n24136), .IN4(n28851), .Q(
        n24100) );
  OA22X1 U27508 ( .IN1(n24139), .IN2(n28845), .IN3(n24141), .IN4(n28849), .Q(
        n24099) );
  OA22X1 U27509 ( .IN1(n24143), .IN2(n28843), .IN3(n24127), .IN4(n28852), .Q(
        n24098) );
  OA22X1 U27510 ( .IN1(n24140), .IN2(n28848), .IN3(n24096), .IN4(n28846), .Q(
        n24097) );
  NAND4X0 U27511 ( .IN1(n24100), .IN2(n24099), .IN3(n24098), .IN4(n24097), 
        .QN(s14_addr_o[23]) );
  OA22X1 U27512 ( .IN1(n28864), .IN2(n24129), .IN3(n28863), .IN4(n24140), .Q(
        n24104) );
  OA22X1 U27513 ( .IN1(n28865), .IN2(n24137), .IN3(n28857), .IN4(n24122), .Q(
        n24103) );
  OA22X1 U27514 ( .IN1(n28860), .IN2(n24128), .IN3(n28859), .IN4(n24117), .Q(
        n24102) );
  OA22X1 U27515 ( .IN1(n28858), .IN2(n24130), .IN3(n28861), .IN4(n24127), .Q(
        n24101) );
  NAND4X0 U27516 ( .IN1(n24104), .IN2(n24103), .IN3(n24102), .IN4(n24101), 
        .QN(s14_addr_o[24]) );
  OA22X1 U27517 ( .IN1(n28877), .IN2(n24139), .IN3(n28870), .IN4(n24140), .Q(
        n24108) );
  OA22X1 U27518 ( .IN1(n28871), .IN2(n24137), .IN3(n28872), .IN4(n24142), .Q(
        n24107) );
  OA22X1 U27519 ( .IN1(n28873), .IN2(n24143), .IN3(n28875), .IN4(n24128), .Q(
        n24106) );
  OA22X1 U27520 ( .IN1(n28876), .IN2(n24141), .IN3(n28874), .IN4(n24122), .Q(
        n24105) );
  NAND4X0 U27521 ( .IN1(n24108), .IN2(n24107), .IN3(n24106), .IN4(n24105), 
        .QN(s14_addr_o[25]) );
  OA22X1 U27522 ( .IN1(n28885), .IN2(n24130), .IN3(n28889), .IN4(n24136), .Q(
        n24112) );
  OA22X1 U27523 ( .IN1(n28887), .IN2(n24129), .IN3(n28882), .IN4(n24138), .Q(
        n24111) );
  OA22X1 U27524 ( .IN1(n28884), .IN2(n24140), .IN3(n28886), .IN4(n24142), .Q(
        n24110) );
  OA22X1 U27525 ( .IN1(n28883), .IN2(n24137), .IN3(n28888), .IN4(n24141), .Q(
        n24109) );
  NAND4X0 U27526 ( .IN1(n24112), .IN2(n24111), .IN3(n24110), .IN4(n24109), 
        .QN(s14_addr_o[26]) );
  OA22X1 U27527 ( .IN1(n28896), .IN2(n24141), .IN3(n28894), .IN4(n24140), .Q(
        n24116) );
  OA22X1 U27528 ( .IN1(n28897), .IN2(n24137), .IN3(n28901), .IN4(n24122), .Q(
        n24115) );
  OA22X1 U27529 ( .IN1(n28898), .IN2(n24128), .IN3(n28900), .IN4(n24142), .Q(
        n24114) );
  OA22X1 U27530 ( .IN1(n28899), .IN2(n24143), .IN3(n28895), .IN4(n24139), .Q(
        n24113) );
  NAND4X0 U27531 ( .IN1(n24116), .IN2(n24115), .IN3(n24114), .IN4(n24113), 
        .QN(s14_addr_o[27]) );
  OA22X1 U27532 ( .IN1(n28908), .IN2(n24122), .IN3(n28906), .IN4(n24127), .Q(
        n24121) );
  OA22X1 U27533 ( .IN1(n28913), .IN2(n24136), .IN3(n28910), .IN4(n24117), .Q(
        n24120) );
  OA22X1 U27534 ( .IN1(n28907), .IN2(n24137), .IN3(n28911), .IN4(n24139), .Q(
        n24119) );
  OA22X1 U27535 ( .IN1(n28909), .IN2(n24130), .IN3(n28912), .IN4(n24140), .Q(
        n24118) );
  NAND4X0 U27536 ( .IN1(n24121), .IN2(n24120), .IN3(n24119), .IN4(n24118), 
        .QN(s14_addr_o[28]) );
  OA22X1 U27537 ( .IN1(n28926), .IN2(n24143), .IN3(n28924), .IN4(n24129), .Q(
        n24126) );
  OA22X1 U27538 ( .IN1(n28919), .IN2(n24122), .IN3(n28923), .IN4(n24127), .Q(
        n24125) );
  OA22X1 U27539 ( .IN1(n28920), .IN2(n24141), .IN3(n28925), .IN4(n24140), .Q(
        n24124) );
  OA22X1 U27540 ( .IN1(n28922), .IN2(n24137), .IN3(n28921), .IN4(n24128), .Q(
        n24123) );
  NAND4X0 U27541 ( .IN1(n24126), .IN2(n24125), .IN3(n24124), .IN4(n24123), 
        .QN(s14_addr_o[29]) );
  OA22X1 U27542 ( .IN1(n28937), .IN2(n24137), .IN3(n28936), .IN4(n24141), .Q(
        n24135) );
  OA22X1 U27543 ( .IN1(n28933), .IN2(n24128), .IN3(n28939), .IN4(n24127), .Q(
        n24134) );
  OA22X1 U27544 ( .IN1(n28932), .IN2(n24130), .IN3(n28935), .IN4(n24129), .Q(
        n24133) );
  OA22X1 U27545 ( .IN1(n28931), .IN2(n24131), .IN3(n28940), .IN4(n24138), .Q(
        n24132) );
  NAND4X0 U27546 ( .IN1(n24135), .IN2(n24134), .IN3(n24133), .IN4(n24132), 
        .QN(s14_addr_o[30]) );
  OA22X1 U27547 ( .IN1(n28956), .IN2(n24137), .IN3(n28960), .IN4(n24136), .Q(
        n24147) );
  OA22X1 U27548 ( .IN1(n28952), .IN2(n24139), .IN3(n28958), .IN4(n24138), .Q(
        n24146) );
  OA22X1 U27549 ( .IN1(n28954), .IN2(n24141), .IN3(n28950), .IN4(n24140), .Q(
        n24145) );
  OA22X1 U27550 ( .IN1(n28948), .IN2(n24143), .IN3(n28946), .IN4(n24142), .Q(
        n24144) );
  NAND4X0 U27551 ( .IN1(n24147), .IN2(n24146), .IN3(n24145), .IN4(n24144), 
        .QN(s14_addr_o[31]) );
  INVX0 U27552 ( .INP(m7_stb_i), .ZN(n29368) );
  OA22X1 U27553 ( .IN1(n29368), .IN2(n24149), .IN3(n29330), .IN4(n24148), .Q(
        n24159) );
  OA22X1 U27554 ( .IN1(n29273), .IN2(n24151), .IN3(n29349), .IN4(n24150), .Q(
        n24158) );
  INVX0 U27555 ( .INP(m1_stb_i), .ZN(n29254) );
  OA22X1 U27556 ( .IN1(n29254), .IN2(n24153), .IN3(n29292), .IN4(n24152), .Q(
        n24157) );
  OA22X1 U27557 ( .IN1(n29235), .IN2(n24155), .IN3(n29311), .IN4(n24154), .Q(
        n24156) );
  NAND4X0 U27558 ( .IN1(n24159), .IN2(n24158), .IN3(n24157), .IN4(n24156), 
        .QN(s13_stb_o) );
  INVX0 U27559 ( .INP(n29207), .ZN(n24445) );
  INVX0 U27560 ( .INP(n29209), .ZN(n24427) );
  OA22X1 U27561 ( .IN1(n24445), .IN2(n28123), .IN3(n24427), .IN4(n28122), .Q(
        n24163) );
  INVX0 U27562 ( .INP(n29200), .ZN(n24442) );
  OA22X1 U27563 ( .IN1(n24392), .IN2(n28124), .IN3(n24442), .IN4(n28128), .Q(
        n24162) );
  INVX0 U27564 ( .INP(n29208), .ZN(n24432) );
  INVX0 U27565 ( .INP(n24397), .ZN(n29201) );
  INVX0 U27566 ( .INP(n29201), .ZN(n24444) );
  OA22X1 U27567 ( .IN1(n24432), .IN2(n28127), .IN3(n24444), .IN4(n28121), .Q(
        n24161) );
  INVX0 U27568 ( .INP(n29210), .ZN(n24435) );
  OA22X1 U27569 ( .IN1(n24435), .IN2(n28126), .IN3(n24418), .IN4(n28125), .Q(
        n24160) );
  NAND4X0 U27570 ( .IN1(n24163), .IN2(n24162), .IN3(n24161), .IN4(n24160), 
        .QN(s13_we_o) );
  INVX0 U27571 ( .INP(n24418), .ZN(n29199) );
  INVX0 U27572 ( .INP(n29199), .ZN(n24441) );
  OA22X1 U27573 ( .IN1(n24441), .IN2(n28136), .IN3(n24397), .IN4(n28135), .Q(
        n24167) );
  INVX0 U27574 ( .INP(n29207), .ZN(n24434) );
  INVX0 U27575 ( .INP(n29210), .ZN(n24440) );
  OA22X1 U27576 ( .IN1(n24434), .IN2(n28133), .IN3(n24440), .IN4(n28139), .Q(
        n24166) );
  INVX0 U27577 ( .INP(n29202), .ZN(n24447) );
  OA22X1 U27578 ( .IN1(n24447), .IN2(n28134), .IN3(n24442), .IN4(n28140), .Q(
        n24165) );
  INVX0 U27579 ( .INP(n29208), .ZN(n24443) );
  OA22X1 U27580 ( .IN1(n24427), .IN2(n28138), .IN3(n24443), .IN4(n28137), .Q(
        n24164) );
  NAND4X0 U27581 ( .IN1(n24167), .IN2(n24166), .IN3(n24165), .IN4(n24164), 
        .QN(s13_data_o[0]) );
  OA22X1 U27582 ( .IN1(n24440), .IN2(n28145), .IN3(n24432), .IN4(n28151), .Q(
        n24171) );
  INVX0 U27583 ( .INP(n29200), .ZN(n24433) );
  INVX0 U27584 ( .INP(n29209), .ZN(n24446) );
  OA22X1 U27585 ( .IN1(n24433), .IN2(n28146), .IN3(n24446), .IN4(n28149), .Q(
        n24170) );
  OA22X1 U27586 ( .IN1(n24441), .IN2(n28152), .IN3(n24397), .IN4(n28147), .Q(
        n24169) );
  OA22X1 U27587 ( .IN1(n24447), .IN2(n28150), .IN3(n24434), .IN4(n28148), .Q(
        n24168) );
  NAND4X0 U27588 ( .IN1(n24171), .IN2(n24170), .IN3(n24169), .IN4(n24168), 
        .QN(s13_data_o[1]) );
  OA22X1 U27589 ( .IN1(n24442), .IN2(n28164), .IN3(n24397), .IN4(n28161), .Q(
        n24175) );
  OA22X1 U27590 ( .IN1(n24434), .IN2(n28163), .IN3(n24446), .IN4(n28158), .Q(
        n24174) );
  OA22X1 U27591 ( .IN1(n24447), .IN2(n28160), .IN3(n24418), .IN4(n28162), .Q(
        n24173) );
  OA22X1 U27592 ( .IN1(n24435), .IN2(n28159), .IN3(n24432), .IN4(n28157), .Q(
        n24172) );
  NAND4X0 U27593 ( .IN1(n24175), .IN2(n24174), .IN3(n24173), .IN4(n24172), 
        .QN(s13_data_o[2]) );
  OA22X1 U27594 ( .IN1(n24441), .IN2(n28175), .IN3(n24397), .IN4(n28173), .Q(
        n24179) );
  OA22X1 U27595 ( .IN1(n24446), .IN2(n28171), .IN3(n24432), .IN4(n28169), .Q(
        n24178) );
  OA22X1 U27596 ( .IN1(n24392), .IN2(n28172), .IN3(n24434), .IN4(n28176), .Q(
        n24177) );
  OA22X1 U27597 ( .IN1(n24433), .IN2(n28174), .IN3(n24440), .IN4(n28170), .Q(
        n24176) );
  NAND4X0 U27598 ( .IN1(n24179), .IN2(n24178), .IN3(n24177), .IN4(n24176), 
        .QN(s13_data_o[3]) );
  OA22X1 U27599 ( .IN1(n24447), .IN2(n28182), .IN3(n24432), .IN4(n28187), .Q(
        n24183) );
  OA22X1 U27600 ( .IN1(n24427), .IN2(n28185), .IN3(n24418), .IN4(n28183), .Q(
        n24182) );
  OA22X1 U27601 ( .IN1(n24440), .IN2(n28188), .IN3(n24397), .IN4(n28181), .Q(
        n24181) );
  OA22X1 U27602 ( .IN1(n24442), .IN2(n28184), .IN3(n24434), .IN4(n28186), .Q(
        n24180) );
  NAND4X0 U27603 ( .IN1(n24183), .IN2(n24182), .IN3(n24181), .IN4(n24180), 
        .QN(s13_data_o[4]) );
  OA22X1 U27604 ( .IN1(n24435), .IN2(n28193), .IN3(n24432), .IN4(n28195), .Q(
        n24187) );
  OA22X1 U27605 ( .IN1(n24434), .IN2(n28194), .IN3(n24397), .IN4(n28199), .Q(
        n24186) );
  OA22X1 U27606 ( .IN1(n24442), .IN2(n28200), .IN3(n24446), .IN4(n28198), .Q(
        n24185) );
  OA22X1 U27607 ( .IN1(n24392), .IN2(n28196), .IN3(n24418), .IN4(n28197), .Q(
        n24184) );
  NAND4X0 U27608 ( .IN1(n24187), .IN2(n24186), .IN3(n24185), .IN4(n24184), 
        .QN(s13_data_o[5]) );
  OA22X1 U27609 ( .IN1(n24442), .IN2(n28207), .IN3(n24434), .IN4(n28206), .Q(
        n24191) );
  OA22X1 U27610 ( .IN1(n24447), .IN2(n28208), .IN3(n24418), .IN4(n28205), .Q(
        n24190) );
  OA22X1 U27611 ( .IN1(n24443), .IN2(n28210), .IN3(n24397), .IN4(n28209), .Q(
        n24189) );
  OA22X1 U27612 ( .IN1(n24435), .IN2(n28212), .IN3(n24446), .IN4(n28211), .Q(
        n24188) );
  NAND4X0 U27613 ( .IN1(n24191), .IN2(n24190), .IN3(n24189), .IN4(n24188), 
        .QN(s13_data_o[6]) );
  OA22X1 U27614 ( .IN1(n24434), .IN2(n28224), .IN3(n24418), .IN4(n28223), .Q(
        n24195) );
  OA22X1 U27615 ( .IN1(n24392), .IN2(n28220), .IN3(n24432), .IN4(n28222), .Q(
        n24194) );
  OA22X1 U27616 ( .IN1(n24435), .IN2(n28218), .IN3(n24446), .IN4(n28217), .Q(
        n24193) );
  OA22X1 U27617 ( .IN1(n24433), .IN2(n28219), .IN3(n24444), .IN4(n28221), .Q(
        n24192) );
  NAND4X0 U27618 ( .IN1(n24195), .IN2(n24194), .IN3(n24193), .IN4(n24192), 
        .QN(s13_data_o[7]) );
  OA22X1 U27619 ( .IN1(n24434), .IN2(n28231), .IN3(n24446), .IN4(n28236), .Q(
        n24199) );
  OA22X1 U27620 ( .IN1(n24447), .IN2(n28230), .IN3(n24444), .IN4(n28235), .Q(
        n24198) );
  OA22X1 U27621 ( .IN1(n24441), .IN2(n28229), .IN3(n24432), .IN4(n28233), .Q(
        n24197) );
  OA22X1 U27622 ( .IN1(n24442), .IN2(n28232), .IN3(n24435), .IN4(n28234), .Q(
        n24196) );
  NAND4X0 U27623 ( .IN1(n24199), .IN2(n24198), .IN3(n24197), .IN4(n24196), 
        .QN(s13_data_o[8]) );
  OA22X1 U27624 ( .IN1(n24446), .IN2(n28241), .IN3(n24418), .IN4(n28245), .Q(
        n24203) );
  OA22X1 U27625 ( .IN1(n24392), .IN2(n28242), .IN3(n24444), .IN4(n28247), .Q(
        n24202) );
  OA22X1 U27626 ( .IN1(n24445), .IN2(n28246), .IN3(n24435), .IN4(n28248), .Q(
        n24201) );
  OA22X1 U27627 ( .IN1(n24433), .IN2(n28244), .IN3(n24432), .IN4(n28243), .Q(
        n24200) );
  NAND4X0 U27628 ( .IN1(n24203), .IN2(n24202), .IN3(n24201), .IN4(n24200), 
        .QN(s13_data_o[9]) );
  OA22X1 U27629 ( .IN1(n24440), .IN2(n28256), .IN3(n24418), .IN4(n28255), .Q(
        n24207) );
  OA22X1 U27630 ( .IN1(n24442), .IN2(n28257), .IN3(n24446), .IN4(n28254), .Q(
        n24206) );
  OA22X1 U27631 ( .IN1(n24445), .IN2(n28260), .IN3(n24444), .IN4(n28259), .Q(
        n24205) );
  OA22X1 U27632 ( .IN1(n24447), .IN2(n28258), .IN3(n24432), .IN4(n28253), .Q(
        n24204) );
  NAND4X0 U27633 ( .IN1(n24207), .IN2(n24206), .IN3(n24205), .IN4(n24204), 
        .QN(s13_data_o[10]) );
  OA22X1 U27634 ( .IN1(n24392), .IN2(n28266), .IN3(n24434), .IN4(n28265), .Q(
        n24211) );
  OA22X1 U27635 ( .IN1(n24441), .IN2(n28270), .IN3(n24444), .IN4(n28269), .Q(
        n24210) );
  OA22X1 U27636 ( .IN1(n24433), .IN2(n28272), .IN3(n24446), .IN4(n28268), .Q(
        n24209) );
  OA22X1 U27637 ( .IN1(n24440), .IN2(n28271), .IN3(n24443), .IN4(n28267), .Q(
        n24208) );
  NAND4X0 U27638 ( .IN1(n24211), .IN2(n24210), .IN3(n24209), .IN4(n24208), 
        .QN(s13_data_o[11]) );
  OA22X1 U27639 ( .IN1(n24433), .IN2(n28278), .IN3(n24443), .IN4(n28279), .Q(
        n24215) );
  OA22X1 U27640 ( .IN1(n24447), .IN2(n28284), .IN3(n24446), .IN4(n28283), .Q(
        n24214) );
  OA22X1 U27641 ( .IN1(n24445), .IN2(n28280), .IN3(n24444), .IN4(n28277), .Q(
        n24213) );
  OA22X1 U27642 ( .IN1(n24435), .IN2(n28282), .IN3(n24418), .IN4(n28281), .Q(
        n24212) );
  NAND4X0 U27643 ( .IN1(n24215), .IN2(n24214), .IN3(n24213), .IN4(n24212), 
        .QN(s13_data_o[12]) );
  OA22X1 U27644 ( .IN1(n24442), .IN2(n28294), .IN3(n24434), .IN4(n28296), .Q(
        n24219) );
  OA22X1 U27645 ( .IN1(n24418), .IN2(n28293), .IN3(n24443), .IN4(n28291), .Q(
        n24218) );
  OA22X1 U27646 ( .IN1(n24440), .IN2(n28292), .IN3(n24444), .IN4(n28295), .Q(
        n24217) );
  OA22X1 U27647 ( .IN1(n24392), .IN2(n28290), .IN3(n24446), .IN4(n28289), .Q(
        n24216) );
  NAND4X0 U27648 ( .IN1(n24219), .IN2(n24218), .IN3(n24217), .IN4(n24216), 
        .QN(s13_data_o[13]) );
  OA22X1 U27649 ( .IN1(n24418), .IN2(n28302), .IN3(n24443), .IN4(n28301), .Q(
        n24223) );
  OA22X1 U27650 ( .IN1(n24427), .IN2(n28307), .IN3(n24444), .IN4(n28303), .Q(
        n24222) );
  OA22X1 U27651 ( .IN1(n24447), .IN2(n28306), .IN3(n24434), .IN4(n28308), .Q(
        n24221) );
  OA22X1 U27652 ( .IN1(n24433), .IN2(n28304), .IN3(n24440), .IN4(n28305), .Q(
        n24220) );
  NAND4X0 U27653 ( .IN1(n24223), .IN2(n24222), .IN3(n24221), .IN4(n24220), 
        .QN(s13_data_o[14]) );
  OA22X1 U27654 ( .IN1(n24442), .IN2(n28315), .IN3(n24444), .IN4(n28319), .Q(
        n24227) );
  OA22X1 U27655 ( .IN1(n24392), .IN2(n28316), .IN3(n24435), .IN4(n28313), .Q(
        n24226) );
  OA22X1 U27656 ( .IN1(n24446), .IN2(n28320), .IN3(n24418), .IN4(n28318), .Q(
        n24225) );
  OA22X1 U27657 ( .IN1(n24445), .IN2(n28314), .IN3(n24443), .IN4(n28317), .Q(
        n24224) );
  NAND4X0 U27658 ( .IN1(n24227), .IN2(n24226), .IN3(n24225), .IN4(n24224), 
        .QN(s13_data_o[15]) );
  OA22X1 U27659 ( .IN1(n24442), .IN2(n28332), .IN3(n24434), .IN4(n28331), .Q(
        n24231) );
  OA22X1 U27660 ( .IN1(n24427), .IN2(n28329), .IN3(n24418), .IN4(n28325), .Q(
        n24230) );
  OA22X1 U27661 ( .IN1(n24432), .IN2(n28328), .IN3(n24444), .IN4(n28327), .Q(
        n24229) );
  OA22X1 U27662 ( .IN1(n24447), .IN2(n28330), .IN3(n24440), .IN4(n28326), .Q(
        n24228) );
  NAND4X0 U27663 ( .IN1(n24231), .IN2(n24230), .IN3(n24229), .IN4(n24228), 
        .QN(s13_data_o[16]) );
  OA22X1 U27664 ( .IN1(n24434), .IN2(n28342), .IN3(n24441), .IN4(n28339), .Q(
        n24235) );
  OA22X1 U27665 ( .IN1(n24392), .IN2(n28340), .IN3(n24444), .IN4(n28341), .Q(
        n24234) );
  OA22X1 U27666 ( .IN1(n24435), .IN2(n28338), .IN3(n24446), .IN4(n28337), .Q(
        n24233) );
  OA22X1 U27667 ( .IN1(n24433), .IN2(n28344), .IN3(n24443), .IN4(n28343), .Q(
        n24232) );
  NAND4X0 U27668 ( .IN1(n24235), .IN2(n24234), .IN3(n24233), .IN4(n24232), 
        .QN(s13_data_o[17]) );
  OA22X1 U27669 ( .IN1(n24435), .IN2(n28355), .IN3(n24441), .IN4(n28349), .Q(
        n24239) );
  OA22X1 U27670 ( .IN1(n24392), .IN2(n28352), .IN3(n24444), .IN4(n28353), .Q(
        n24238) );
  OA22X1 U27671 ( .IN1(n24442), .IN2(n28356), .IN3(n24443), .IN4(n28351), .Q(
        n24237) );
  OA22X1 U27672 ( .IN1(n24445), .IN2(n28350), .IN3(n24427), .IN4(n28354), .Q(
        n24236) );
  NAND4X0 U27673 ( .IN1(n24239), .IN2(n24238), .IN3(n24237), .IN4(n24236), 
        .QN(s13_data_o[18]) );
  OA22X1 U27674 ( .IN1(n24392), .IN2(n28366), .IN3(n24443), .IN4(n28368), .Q(
        n24243) );
  OA22X1 U27675 ( .IN1(n24446), .IN2(n28365), .IN3(n24444), .IN4(n28367), .Q(
        n24242) );
  OA22X1 U27676 ( .IN1(n24434), .IN2(n28362), .IN3(n24441), .IN4(n28361), .Q(
        n24241) );
  OA22X1 U27677 ( .IN1(n24442), .IN2(n28364), .IN3(n24435), .IN4(n28363), .Q(
        n24240) );
  NAND4X0 U27678 ( .IN1(n24243), .IN2(n24242), .IN3(n24241), .IN4(n24240), 
        .QN(s13_data_o[19]) );
  OA22X1 U27679 ( .IN1(n24440), .IN2(n28373), .IN3(n24443), .IN4(n28379), .Q(
        n24247) );
  OA22X1 U27680 ( .IN1(n24392), .IN2(n28378), .IN3(n24442), .IN4(n28377), .Q(
        n24246) );
  OA22X1 U27681 ( .IN1(n24427), .IN2(n28376), .IN3(n24441), .IN4(n28380), .Q(
        n24245) );
  OA22X1 U27682 ( .IN1(n24434), .IN2(n28374), .IN3(n24444), .IN4(n28375), .Q(
        n24244) );
  NAND4X0 U27683 ( .IN1(n24247), .IN2(n24246), .IN3(n24245), .IN4(n24244), 
        .QN(s13_data_o[20]) );
  OA22X1 U27684 ( .IN1(n24440), .IN2(n28388), .IN3(n24441), .IN4(n28385), .Q(
        n24251) );
  OA22X1 U27685 ( .IN1(n24433), .IN2(n28386), .IN3(n24445), .IN4(n28390), .Q(
        n24250) );
  OA22X1 U27686 ( .IN1(n24392), .IN2(n28392), .IN3(n24444), .IN4(n28391), .Q(
        n24249) );
  OA22X1 U27687 ( .IN1(n24427), .IN2(n28387), .IN3(n24443), .IN4(n28389), .Q(
        n24248) );
  NAND4X0 U27688 ( .IN1(n24251), .IN2(n24250), .IN3(n24249), .IN4(n24248), 
        .QN(s13_data_o[21]) );
  OA22X1 U27689 ( .IN1(n24392), .IN2(n28400), .IN3(n24427), .IN4(n28398), .Q(
        n24255) );
  OA22X1 U27690 ( .IN1(n24435), .IN2(n28403), .IN3(n24443), .IN4(n28401), .Q(
        n24254) );
  OA22X1 U27691 ( .IN1(n24433), .IN2(n28402), .IN3(n24441), .IN4(n28399), .Q(
        n24253) );
  OA22X1 U27692 ( .IN1(n24445), .IN2(n28404), .IN3(n24444), .IN4(n28397), .Q(
        n24252) );
  NAND4X0 U27693 ( .IN1(n24255), .IN2(n24254), .IN3(n24253), .IN4(n24252), 
        .QN(s13_data_o[22]) );
  OA22X1 U27694 ( .IN1(n24392), .IN2(n28416), .IN3(n24434), .IN4(n28414), .Q(
        n24259) );
  OA22X1 U27695 ( .IN1(n24418), .IN2(n28412), .IN3(n24443), .IN4(n28409), .Q(
        n24258) );
  OA22X1 U27696 ( .IN1(n24435), .IN2(n28413), .IN3(n24397), .IN4(n28411), .Q(
        n24257) );
  OA22X1 U27697 ( .IN1(n24442), .IN2(n28415), .IN3(n24446), .IN4(n28410), .Q(
        n24256) );
  NAND4X0 U27698 ( .IN1(n24259), .IN2(n24258), .IN3(n24257), .IN4(n24256), 
        .QN(s13_data_o[23]) );
  OA22X1 U27699 ( .IN1(n24392), .IN2(n28426), .IN3(n24443), .IN4(n28427), .Q(
        n24263) );
  OA22X1 U27700 ( .IN1(n24435), .IN2(n28421), .IN3(n24441), .IN4(n28428), .Q(
        n24262) );
  OA22X1 U27701 ( .IN1(n24445), .IN2(n28422), .IN3(n24397), .IN4(n28423), .Q(
        n24261) );
  OA22X1 U27702 ( .IN1(n24433), .IN2(n28424), .IN3(n24446), .IN4(n28425), .Q(
        n24260) );
  NAND4X0 U27703 ( .IN1(n24263), .IN2(n24262), .IN3(n24261), .IN4(n24260), 
        .QN(s13_data_o[24]) );
  OA22X1 U27704 ( .IN1(n24435), .IN2(n28439), .IN3(n24427), .IN4(n28433), .Q(
        n24267) );
  OA22X1 U27705 ( .IN1(n24392), .IN2(n28438), .IN3(n24397), .IN4(n28435), .Q(
        n24266) );
  OA22X1 U27706 ( .IN1(n24434), .IN2(n28434), .IN3(n24443), .IN4(n28436), .Q(
        n24265) );
  OA22X1 U27707 ( .IN1(n24442), .IN2(n28440), .IN3(n24441), .IN4(n28437), .Q(
        n24264) );
  NAND4X0 U27708 ( .IN1(n24267), .IN2(n24266), .IN3(n24265), .IN4(n24264), 
        .QN(s13_data_o[25]) );
  OA22X1 U27709 ( .IN1(n24392), .IN2(n28452), .IN3(n24442), .IN4(n28451), .Q(
        n24271) );
  OA22X1 U27710 ( .IN1(n24435), .IN2(n28446), .IN3(n24441), .IN4(n28448), .Q(
        n24270) );
  OA22X1 U27711 ( .IN1(n24446), .IN2(n28449), .IN3(n24397), .IN4(n28445), .Q(
        n24269) );
  OA22X1 U27712 ( .IN1(n24445), .IN2(n28450), .IN3(n24443), .IN4(n28447), .Q(
        n24268) );
  NAND4X0 U27713 ( .IN1(n24271), .IN2(n24270), .IN3(n24269), .IN4(n24268), 
        .QN(s13_data_o[26]) );
  OA22X1 U27714 ( .IN1(n24442), .IN2(n28461), .IN3(n24440), .IN4(n28458), .Q(
        n24275) );
  OA22X1 U27715 ( .IN1(n24392), .IN2(n28462), .IN3(n24397), .IN4(n28459), .Q(
        n24274) );
  OA22X1 U27716 ( .IN1(n24434), .IN2(n28464), .IN3(n24443), .IN4(n28460), .Q(
        n24273) );
  OA22X1 U27717 ( .IN1(n24427), .IN2(n28457), .IN3(n24441), .IN4(n28463), .Q(
        n24272) );
  NAND4X0 U27718 ( .IN1(n24275), .IN2(n24274), .IN3(n24273), .IN4(n24272), 
        .QN(s13_data_o[27]) );
  OA22X1 U27719 ( .IN1(n24445), .IN2(n28472), .IN3(n24441), .IN4(n28475), .Q(
        n24279) );
  OA22X1 U27720 ( .IN1(n24392), .IN2(n28474), .IN3(n24442), .IN4(n28476), .Q(
        n24278) );
  OA22X1 U27721 ( .IN1(n24435), .IN2(n28470), .IN3(n24446), .IN4(n28471), .Q(
        n24277) );
  OA22X1 U27722 ( .IN1(n24443), .IN2(n28469), .IN3(n24397), .IN4(n28473), .Q(
        n24276) );
  NAND4X0 U27723 ( .IN1(n24279), .IN2(n24278), .IN3(n24277), .IN4(n24276), 
        .QN(s13_data_o[28]) );
  OA22X1 U27724 ( .IN1(n24432), .IN2(n28485), .IN3(n24397), .IN4(n28481), .Q(
        n24283) );
  OA22X1 U27725 ( .IN1(n24392), .IN2(n28484), .IN3(n24441), .IN4(n28483), .Q(
        n24282) );
  OA22X1 U27726 ( .IN1(n24445), .IN2(n28488), .IN3(n24435), .IN4(n28486), .Q(
        n24281) );
  OA22X1 U27727 ( .IN1(n24433), .IN2(n28482), .IN3(n24427), .IN4(n28487), .Q(
        n24280) );
  NAND4X0 U27728 ( .IN1(n24283), .IN2(n24282), .IN3(n24281), .IN4(n24280), 
        .QN(s13_data_o[29]) );
  OA22X1 U27729 ( .IN1(n24445), .IN2(n28497), .IN3(n24432), .IN4(n28500), .Q(
        n24287) );
  OA22X1 U27730 ( .IN1(n24392), .IN2(n28494), .IN3(n24427), .IN4(n28493), .Q(
        n24286) );
  OA22X1 U27731 ( .IN1(n24435), .IN2(n28496), .IN3(n24441), .IN4(n28495), .Q(
        n24285) );
  OA22X1 U27732 ( .IN1(n24433), .IN2(n28498), .IN3(n24397), .IN4(n28499), .Q(
        n24284) );
  NAND4X0 U27733 ( .IN1(n24287), .IN2(n24286), .IN3(n24285), .IN4(n24284), 
        .QN(s13_data_o[30]) );
  OA22X1 U27734 ( .IN1(n24442), .IN2(n28509), .IN3(n24432), .IN4(n28511), .Q(
        n24291) );
  OA22X1 U27735 ( .IN1(n24435), .IN2(n28505), .IN3(n24441), .IN4(n28508), .Q(
        n24290) );
  OA22X1 U27736 ( .IN1(n24392), .IN2(n28510), .IN3(n24397), .IN4(n28507), .Q(
        n24289) );
  OA22X1 U27737 ( .IN1(n24445), .IN2(n28506), .IN3(n24446), .IN4(n28512), .Q(
        n24288) );
  NAND4X0 U27738 ( .IN1(n24291), .IN2(n24290), .IN3(n24289), .IN4(n24288), 
        .QN(s13_data_o[31]) );
  OA22X1 U27739 ( .IN1(n24435), .IN2(n28524), .IN3(n24441), .IN4(n28520), .Q(
        n24295) );
  OA22X1 U27740 ( .IN1(n24433), .IN2(n28517), .IN3(n24397), .IN4(n28519), .Q(
        n24294) );
  OA22X1 U27741 ( .IN1(n24447), .IN2(n28518), .IN3(n24445), .IN4(n28522), .Q(
        n24293) );
  OA22X1 U27742 ( .IN1(n24427), .IN2(n28523), .IN3(n24432), .IN4(n28521), .Q(
        n24292) );
  NAND4X0 U27743 ( .IN1(n24295), .IN2(n24294), .IN3(n24293), .IN4(n24292), 
        .QN(s13_sel_o[0]) );
  OA22X1 U27744 ( .IN1(n24442), .IN2(n28532), .IN3(n24435), .IN4(n28536), .Q(
        n24299) );
  OA22X1 U27745 ( .IN1(n24432), .IN2(n28531), .IN3(n24397), .IN4(n28529), .Q(
        n24298) );
  OA22X1 U27746 ( .IN1(n24445), .IN2(n28530), .IN3(n24441), .IN4(n28533), .Q(
        n24297) );
  OA22X1 U27747 ( .IN1(n24447), .IN2(n28534), .IN3(n24446), .IN4(n28535), .Q(
        n24296) );
  NAND4X0 U27748 ( .IN1(n24299), .IN2(n24298), .IN3(n24297), .IN4(n24296), 
        .QN(s13_sel_o[1]) );
  OA22X1 U27749 ( .IN1(n24435), .IN2(n28548), .IN3(n24432), .IN4(n28545), .Q(
        n24303) );
  OA22X1 U27750 ( .IN1(n24442), .IN2(n28546), .IN3(n24418), .IN4(n28542), .Q(
        n24302) );
  OA22X1 U27751 ( .IN1(n24447), .IN2(n28544), .IN3(n24445), .IN4(n28543), .Q(
        n24301) );
  OA22X1 U27752 ( .IN1(n24427), .IN2(n28547), .IN3(n24397), .IN4(n28541), .Q(
        n24300) );
  NAND4X0 U27753 ( .IN1(n24303), .IN2(n24302), .IN3(n24301), .IN4(n24300), 
        .QN(s13_sel_o[2]) );
  OA22X1 U27754 ( .IN1(n24447), .IN2(n28558), .IN3(n24440), .IN4(n28557), .Q(
        n24307) );
  OA22X1 U27755 ( .IN1(n24427), .IN2(n28556), .IN3(n24397), .IN4(n28555), .Q(
        n24306) );
  OA22X1 U27756 ( .IN1(n24445), .IN2(n28553), .IN3(n24418), .IN4(n28560), .Q(
        n24305) );
  OA22X1 U27757 ( .IN1(n24433), .IN2(n28554), .IN3(n24432), .IN4(n28559), .Q(
        n24304) );
  NAND4X0 U27758 ( .IN1(n24307), .IN2(n24306), .IN3(n24305), .IN4(n24304), 
        .QN(s13_sel_o[3]) );
  OA22X1 U27759 ( .IN1(n24447), .IN2(n28572), .IN3(n24427), .IN4(n28568), .Q(
        n24311) );
  OA22X1 U27760 ( .IN1(n24435), .IN2(n28566), .IN3(n24397), .IN4(n28569), .Q(
        n24310) );
  OA22X1 U27761 ( .IN1(n24442), .IN2(n28570), .IN3(n24434), .IN4(n28571), .Q(
        n24309) );
  OA22X1 U27762 ( .IN1(n24418), .IN2(n28567), .IN3(n24432), .IN4(n28565), .Q(
        n24308) );
  NAND4X0 U27763 ( .IN1(n24311), .IN2(n24310), .IN3(n24309), .IN4(n24308), 
        .QN(s13_addr_o[0]) );
  OA22X1 U27764 ( .IN1(n24435), .IN2(n28581), .IN3(n24397), .IN4(n28583), .Q(
        n24315) );
  OA22X1 U27765 ( .IN1(n24392), .IN2(n28580), .IN3(n24445), .IN4(n28582), .Q(
        n24314) );
  OA22X1 U27766 ( .IN1(n24427), .IN2(n28579), .IN3(n24418), .IN4(n28584), .Q(
        n24313) );
  OA22X1 U27767 ( .IN1(n24433), .IN2(n28578), .IN3(n24432), .IN4(n28577), .Q(
        n24312) );
  NAND4X0 U27768 ( .IN1(n24315), .IN2(n24314), .IN3(n24313), .IN4(n24312), 
        .QN(s13_addr_o[1]) );
  OA22X1 U27769 ( .IN1(n28594), .IN2(n24434), .IN3(n28590), .IN4(n24446), .Q(
        n24319) );
  OA22X1 U27770 ( .IN1(n28591), .IN2(n24447), .IN3(n28593), .IN4(n24418), .Q(
        n24318) );
  OA22X1 U27771 ( .IN1(n28589), .IN2(n24433), .IN3(n28595), .IN4(n24432), .Q(
        n24317) );
  OA22X1 U27772 ( .IN1(n28592), .IN2(n24440), .IN3(n28596), .IN4(n24444), .Q(
        n24316) );
  NAND4X0 U27773 ( .IN1(n24319), .IN2(n24318), .IN3(n24317), .IN4(n24316), 
        .QN(s13_addr_o[2]) );
  OA22X1 U27774 ( .IN1(n28602), .IN2(n24441), .IN3(n28604), .IN4(n24434), .Q(
        n24323) );
  OA22X1 U27775 ( .IN1(n28601), .IN2(n24392), .IN3(n28608), .IN4(n24444), .Q(
        n24322) );
  OA22X1 U27776 ( .IN1(n28606), .IN2(n24446), .IN3(n28605), .IN4(n24442), .Q(
        n24321) );
  OA22X1 U27777 ( .IN1(n28603), .IN2(n24432), .IN3(n28607), .IN4(n24440), .Q(
        n24320) );
  NAND4X0 U27778 ( .IN1(n24323), .IN2(n24322), .IN3(n24321), .IN4(n24320), 
        .QN(s13_addr_o[3]) );
  OA22X1 U27779 ( .IN1(n28618), .IN2(n24435), .IN3(n28615), .IN4(n24446), .Q(
        n24327) );
  OA22X1 U27780 ( .IN1(n28620), .IN2(n24443), .IN3(n28614), .IN4(n24418), .Q(
        n24326) );
  OA22X1 U27781 ( .IN1(n28619), .IN2(n24444), .IN3(n28617), .IN4(n24447), .Q(
        n24325) );
  OA22X1 U27782 ( .IN1(n28616), .IN2(n24433), .IN3(n28613), .IN4(n24434), .Q(
        n24324) );
  NAND4X0 U27783 ( .IN1(n24327), .IN2(n24326), .IN3(n24325), .IN4(n24324), 
        .QN(s13_addr_o[4]) );
  OA22X1 U27784 ( .IN1(n28632), .IN2(n24445), .IN3(n28628), .IN4(n24443), .Q(
        n24331) );
  OA22X1 U27785 ( .IN1(n28630), .IN2(n24433), .IN3(n28629), .IN4(n24447), .Q(
        n24330) );
  OA22X1 U27786 ( .IN1(n28627), .IN2(n24441), .IN3(n28631), .IN4(n24446), .Q(
        n24329) );
  OA22X1 U27787 ( .IN1(n28626), .IN2(n24440), .IN3(n28625), .IN4(n24444), .Q(
        n24328) );
  NAND4X0 U27788 ( .IN1(n24331), .IN2(n24330), .IN3(n24329), .IN4(n24328), 
        .QN(s13_addr_o[5]) );
  OA22X1 U27789 ( .IN1(n24440), .IN2(n28643), .IN3(n24397), .IN4(n28639), .Q(
        n24335) );
  OA22X1 U27790 ( .IN1(n24427), .IN2(n28638), .IN3(n24443), .IN4(n28641), .Q(
        n24334) );
  OA22X1 U27791 ( .IN1(n24392), .IN2(n28642), .IN3(n24442), .IN4(n28640), .Q(
        n24333) );
  OA22X1 U27792 ( .IN1(n24445), .IN2(n28644), .IN3(n24418), .IN4(n28637), .Q(
        n24332) );
  NAND4X0 U27793 ( .IN1(n24335), .IN2(n24334), .IN3(n24333), .IN4(n24332), 
        .QN(s13_addr_o[6]) );
  OA22X1 U27794 ( .IN1(n24442), .IN2(n28652), .IN3(n24434), .IN4(n28656), .Q(
        n24339) );
  OA22X1 U27795 ( .IN1(n24392), .IN2(n28654), .IN3(n24440), .IN4(n28653), .Q(
        n24338) );
  OA22X1 U27796 ( .IN1(n24427), .IN2(n28650), .IN3(n24432), .IN4(n28651), .Q(
        n24337) );
  OA22X1 U27797 ( .IN1(n24418), .IN2(n28649), .IN3(n24397), .IN4(n28655), .Q(
        n24336) );
  NAND4X0 U27798 ( .IN1(n24339), .IN2(n24338), .IN3(n24337), .IN4(n24336), 
        .QN(s13_addr_o[7]) );
  OA22X1 U27799 ( .IN1(n24435), .IN2(n28665), .IN3(n24397), .IN4(n28667), .Q(
        n24343) );
  OA22X1 U27800 ( .IN1(n24441), .IN2(n28662), .IN3(n24443), .IN4(n28661), .Q(
        n24342) );
  OA22X1 U27801 ( .IN1(n24447), .IN2(n28664), .IN3(n24445), .IN4(n28666), .Q(
        n24341) );
  OA22X1 U27802 ( .IN1(n24433), .IN2(n28663), .IN3(n24446), .IN4(n28668), .Q(
        n24340) );
  NAND4X0 U27803 ( .IN1(n24343), .IN2(n24342), .IN3(n24341), .IN4(n24340), 
        .QN(s13_addr_o[8]) );
  OA22X1 U27804 ( .IN1(n24447), .IN2(n28680), .IN3(n24427), .IN4(n28673), .Q(
        n24347) );
  OA22X1 U27805 ( .IN1(n24443), .IN2(n28675), .IN3(n24397), .IN4(n28677), .Q(
        n24346) );
  OA22X1 U27806 ( .IN1(n24445), .IN2(n28674), .IN3(n24418), .IN4(n28678), .Q(
        n24345) );
  OA22X1 U27807 ( .IN1(n24433), .IN2(n28679), .IN3(n24440), .IN4(n28676), .Q(
        n24344) );
  NAND4X0 U27808 ( .IN1(n24347), .IN2(n24346), .IN3(n24345), .IN4(n24344), 
        .QN(s13_addr_o[9]) );
  OA22X1 U27809 ( .IN1(n24445), .IN2(n28688), .IN3(n24443), .IN4(n28690), .Q(
        n24351) );
  OA22X1 U27810 ( .IN1(n24442), .IN2(n28686), .IN3(n24427), .IN4(n28685), .Q(
        n24350) );
  OA22X1 U27811 ( .IN1(n24392), .IN2(n28692), .IN3(n24397), .IN4(n28689), .Q(
        n24349) );
  OA22X1 U27812 ( .IN1(n24440), .IN2(n28687), .IN3(n24418), .IN4(n28691), .Q(
        n24348) );
  NAND4X0 U27813 ( .IN1(n24351), .IN2(n24350), .IN3(n24349), .IN4(n24348), 
        .QN(s13_addr_o[10]) );
  OA22X1 U27814 ( .IN1(n24447), .IN2(n28702), .IN3(n24440), .IN4(n28704), .Q(
        n24355) );
  OA22X1 U27815 ( .IN1(n24427), .IN2(n28701), .IN3(n24397), .IN4(n28699), .Q(
        n24354) );
  OA22X1 U27816 ( .IN1(n24442), .IN2(n28698), .IN3(n24434), .IN4(n28697), .Q(
        n24353) );
  OA22X1 U27817 ( .IN1(n24418), .IN2(n28703), .IN3(n24432), .IN4(n28700), .Q(
        n24352) );
  NAND4X0 U27818 ( .IN1(n24355), .IN2(n24354), .IN3(n24353), .IN4(n24352), 
        .QN(s13_addr_o[11]) );
  OA22X1 U27819 ( .IN1(n24433), .IN2(n28710), .IN3(n24432), .IN4(n28711), .Q(
        n24359) );
  OA22X1 U27820 ( .IN1(n24435), .IN2(n28716), .IN3(n24427), .IN4(n28709), .Q(
        n24358) );
  OA22X1 U27821 ( .IN1(n24445), .IN2(n28712), .IN3(n24397), .IN4(n28713), .Q(
        n24357) );
  OA22X1 U27822 ( .IN1(n24447), .IN2(n28714), .IN3(n24418), .IN4(n28715), .Q(
        n24356) );
  NAND4X0 U27823 ( .IN1(n24359), .IN2(n24358), .IN3(n24357), .IN4(n24356), 
        .QN(s13_addr_o[12]) );
  OA22X1 U27824 ( .IN1(n24433), .IN2(n28728), .IN3(n24446), .IN4(n28723), .Q(
        n24363) );
  OA22X1 U27825 ( .IN1(n24443), .IN2(n28725), .IN3(n24397), .IN4(n28727), .Q(
        n24362) );
  OA22X1 U27826 ( .IN1(n24392), .IN2(n28722), .IN3(n24434), .IN4(n28726), .Q(
        n24361) );
  OA22X1 U27827 ( .IN1(n24440), .IN2(n28724), .IN3(n24418), .IN4(n28721), .Q(
        n24360) );
  NAND4X0 U27828 ( .IN1(n24363), .IN2(n24362), .IN3(n24361), .IN4(n24360), 
        .QN(s13_addr_o[13]) );
  OA22X1 U27829 ( .IN1(n24442), .IN2(n28738), .IN3(n24432), .IN4(n28733), .Q(
        n24367) );
  OA22X1 U27830 ( .IN1(n24427), .IN2(n28740), .IN3(n24397), .IN4(n28739), .Q(
        n24366) );
  OA22X1 U27831 ( .IN1(n24392), .IN2(n28734), .IN3(n24440), .IN4(n28735), .Q(
        n24365) );
  OA22X1 U27832 ( .IN1(n24445), .IN2(n28736), .IN3(n24418), .IN4(n28737), .Q(
        n24364) );
  NAND4X0 U27833 ( .IN1(n24367), .IN2(n24366), .IN3(n24365), .IN4(n24364), 
        .QN(s13_addr_o[14]) );
  OA22X1 U27834 ( .IN1(n24434), .IN2(n28750), .IN3(n24440), .IN4(n28752), .Q(
        n24371) );
  OA22X1 U27835 ( .IN1(n24442), .IN2(n28748), .IN3(n24397), .IN4(n28745), .Q(
        n24370) );
  OA22X1 U27836 ( .IN1(n24427), .IN2(n28747), .IN3(n24418), .IN4(n28751), .Q(
        n24369) );
  OA22X1 U27837 ( .IN1(n24392), .IN2(n28746), .IN3(n24443), .IN4(n28749), .Q(
        n24368) );
  NAND4X0 U27838 ( .IN1(n24371), .IN2(n24370), .IN3(n24369), .IN4(n24368), 
        .QN(s13_addr_o[15]) );
  OA22X1 U27839 ( .IN1(n24447), .IN2(n28758), .IN3(n24397), .IN4(n28763), .Q(
        n24375) );
  OA22X1 U27840 ( .IN1(n24433), .IN2(n28762), .IN3(n24434), .IN4(n28760), .Q(
        n24374) );
  OA22X1 U27841 ( .IN1(n24427), .IN2(n28759), .IN3(n24418), .IN4(n28757), .Q(
        n24373) );
  OA22X1 U27842 ( .IN1(n24435), .IN2(n28761), .IN3(n24432), .IN4(n28764), .Q(
        n24372) );
  NAND4X0 U27843 ( .IN1(n24375), .IN2(n24374), .IN3(n24373), .IN4(n24372), 
        .QN(s13_addr_o[16]) );
  OA22X1 U27844 ( .IN1(n24442), .IN2(n28776), .IN3(n24443), .IN4(n28770), .Q(
        n24379) );
  OA22X1 U27845 ( .IN1(n24447), .IN2(n28772), .IN3(n24418), .IN4(n28771), .Q(
        n24378) );
  OA22X1 U27846 ( .IN1(n24427), .IN2(n28775), .IN3(n24397), .IN4(n28769), .Q(
        n24377) );
  OA22X1 U27847 ( .IN1(n24445), .IN2(n28774), .IN3(n24440), .IN4(n28773), .Q(
        n24376) );
  NAND4X0 U27848 ( .IN1(n24379), .IN2(n24378), .IN3(n24377), .IN4(n24376), 
        .QN(s13_addr_o[17]) );
  OA22X1 U27849 ( .IN1(n24433), .IN2(n28788), .IN3(n24434), .IN4(n28787), .Q(
        n24383) );
  OA22X1 U27850 ( .IN1(n24392), .IN2(n28786), .IN3(n24440), .IN4(n28782), .Q(
        n24382) );
  OA22X1 U27851 ( .IN1(n24427), .IN2(n28784), .IN3(n24418), .IN4(n28783), .Q(
        n24381) );
  OA22X1 U27852 ( .IN1(n24432), .IN2(n28785), .IN3(n24397), .IN4(n28781), .Q(
        n24380) );
  NAND4X0 U27853 ( .IN1(n24383), .IN2(n24382), .IN3(n24381), .IN4(n24380), 
        .QN(s13_addr_o[18]) );
  OA22X1 U27854 ( .IN1(n24440), .IN2(n28794), .IN3(n24397), .IN4(n28799), .Q(
        n24387) );
  OA22X1 U27855 ( .IN1(n24447), .IN2(n28796), .IN3(n24442), .IN4(n28800), .Q(
        n24386) );
  OA22X1 U27856 ( .IN1(n24445), .IN2(n28798), .IN3(n24432), .IN4(n28793), .Q(
        n24385) );
  OA22X1 U27857 ( .IN1(n24427), .IN2(n28797), .IN3(n24418), .IN4(n28795), .Q(
        n24384) );
  NAND4X0 U27858 ( .IN1(n24387), .IN2(n24386), .IN3(n24385), .IN4(n24384), 
        .QN(s13_addr_o[19]) );
  OA22X1 U27859 ( .IN1(n24392), .IN2(n28812), .IN3(n24427), .IN4(n28806), .Q(
        n24391) );
  OA22X1 U27860 ( .IN1(n24434), .IN2(n28807), .IN3(n24397), .IN4(n28805), .Q(
        n24390) );
  OA22X1 U27861 ( .IN1(n24435), .IN2(n28810), .IN3(n24418), .IN4(n28811), .Q(
        n24389) );
  OA22X1 U27862 ( .IN1(n24433), .IN2(n28808), .IN3(n24432), .IN4(n28809), .Q(
        n24388) );
  NAND4X0 U27863 ( .IN1(n24391), .IN2(n24390), .IN3(n24389), .IN4(n24388), 
        .QN(s13_addr_o[20]) );
  OA22X1 U27864 ( .IN1(n24392), .IN2(n28822), .IN3(n24418), .IN4(n28823), .Q(
        n24396) );
  OA22X1 U27865 ( .IN1(n24446), .IN2(n28821), .IN3(n24397), .IN4(n28817), .Q(
        n24395) );
  OA22X1 U27866 ( .IN1(n24445), .IN2(n28820), .IN3(n24443), .IN4(n28818), .Q(
        n24394) );
  OA22X1 U27867 ( .IN1(n24433), .IN2(n28824), .IN3(n24440), .IN4(n28819), .Q(
        n24393) );
  NAND4X0 U27868 ( .IN1(n24396), .IN2(n24395), .IN3(n24394), .IN4(n24393), 
        .QN(s13_addr_o[21]) );
  OA22X1 U27869 ( .IN1(n24427), .IN2(n28836), .IN3(n24397), .IN4(n28829), .Q(
        n24401) );
  OA22X1 U27870 ( .IN1(n24445), .IN2(n28831), .IN3(n24443), .IN4(n28837), .Q(
        n24400) );
  OA22X1 U27871 ( .IN1(n24433), .IN2(n28832), .IN3(n24418), .IN4(n28834), .Q(
        n24399) );
  OA22X1 U27872 ( .IN1(n24447), .IN2(n28833), .IN3(n24440), .IN4(n28838), .Q(
        n24398) );
  NAND4X0 U27873 ( .IN1(n24401), .IN2(n24400), .IN3(n24399), .IN4(n24398), 
        .QN(s13_addr_o[22]) );
  OA22X1 U27874 ( .IN1(n24433), .IN2(n28845), .IN3(n24434), .IN4(n28843), .Q(
        n24405) );
  OA22X1 U27875 ( .IN1(n24418), .IN2(n28849), .IN3(n24444), .IN4(n28851), .Q(
        n24404) );
  OA22X1 U27876 ( .IN1(n24447), .IN2(n28848), .IN3(n24443), .IN4(n28846), .Q(
        n24403) );
  OA22X1 U27877 ( .IN1(n24435), .IN2(n28850), .IN3(n24446), .IN4(n28852), .Q(
        n24402) );
  NAND4X0 U27878 ( .IN1(n24405), .IN2(n24404), .IN3(n24403), .IN4(n24402), 
        .QN(s13_addr_o[23]) );
  OA22X1 U27879 ( .IN1(n28858), .IN2(n24434), .IN3(n28857), .IN4(n24440), .Q(
        n24409) );
  OA22X1 U27880 ( .IN1(n28864), .IN2(n24433), .IN3(n28863), .IN4(n24447), .Q(
        n24408) );
  OA22X1 U27881 ( .IN1(n28865), .IN2(n24432), .IN3(n28861), .IN4(n24446), .Q(
        n24407) );
  OA22X1 U27882 ( .IN1(n28860), .IN2(n24444), .IN3(n28859), .IN4(n24418), .Q(
        n24406) );
  NAND4X0 U27883 ( .IN1(n24409), .IN2(n24408), .IN3(n24407), .IN4(n24406), 
        .QN(s13_addr_o[24]) );
  OA22X1 U27884 ( .IN1(n28871), .IN2(n24443), .IN3(n28872), .IN4(n24446), .Q(
        n24413) );
  OA22X1 U27885 ( .IN1(n28877), .IN2(n24433), .IN3(n28876), .IN4(n24418), .Q(
        n24412) );
  OA22X1 U27886 ( .IN1(n28873), .IN2(n24445), .IN3(n28875), .IN4(n24444), .Q(
        n24411) );
  OA22X1 U27887 ( .IN1(n28870), .IN2(n24447), .IN3(n28874), .IN4(n24440), .Q(
        n24410) );
  NAND4X0 U27888 ( .IN1(n24413), .IN2(n24412), .IN3(n24411), .IN4(n24410), 
        .QN(s13_addr_o[25]) );
  OA22X1 U27889 ( .IN1(n28885), .IN2(n24434), .IN3(n28887), .IN4(n24442), .Q(
        n24417) );
  OA22X1 U27890 ( .IN1(n28889), .IN2(n24444), .IN3(n28884), .IN4(n24447), .Q(
        n24416) );
  OA22X1 U27891 ( .IN1(n28888), .IN2(n24441), .IN3(n28886), .IN4(n24446), .Q(
        n24415) );
  OA22X1 U27892 ( .IN1(n28883), .IN2(n24432), .IN3(n28882), .IN4(n24440), .Q(
        n24414) );
  NAND4X0 U27893 ( .IN1(n24417), .IN2(n24416), .IN3(n24415), .IN4(n24414), 
        .QN(s13_addr_o[26]) );
  OA22X1 U27894 ( .IN1(n28901), .IN2(n24435), .IN3(n28900), .IN4(n24446), .Q(
        n24422) );
  OA22X1 U27895 ( .IN1(n28898), .IN2(n24444), .IN3(n28896), .IN4(n24418), .Q(
        n24421) );
  OA22X1 U27896 ( .IN1(n28897), .IN2(n24443), .IN3(n28895), .IN4(n24442), .Q(
        n24420) );
  OA22X1 U27897 ( .IN1(n28899), .IN2(n24445), .IN3(n28894), .IN4(n24447), .Q(
        n24419) );
  NAND4X0 U27898 ( .IN1(n24422), .IN2(n24421), .IN3(n24420), .IN4(n24419), 
        .QN(s13_addr_o[27]) );
  OA22X1 U27899 ( .IN1(n28910), .IN2(n24441), .IN3(n28906), .IN4(n24427), .Q(
        n24426) );
  OA22X1 U27900 ( .IN1(n28907), .IN2(n24432), .IN3(n28913), .IN4(n24444), .Q(
        n24425) );
  OA22X1 U27901 ( .IN1(n28909), .IN2(n24434), .IN3(n28908), .IN4(n24440), .Q(
        n24424) );
  OA22X1 U27902 ( .IN1(n28911), .IN2(n24433), .IN3(n28912), .IN4(n24447), .Q(
        n24423) );
  NAND4X0 U27903 ( .IN1(n24426), .IN2(n24425), .IN3(n24424), .IN4(n24423), 
        .QN(s13_addr_o[28]) );
  OA22X1 U27904 ( .IN1(n28921), .IN2(n24444), .IN3(n28919), .IN4(n24440), .Q(
        n24431) );
  OA22X1 U27905 ( .IN1(n28920), .IN2(n24441), .IN3(n28923), .IN4(n24427), .Q(
        n24430) );
  OA22X1 U27906 ( .IN1(n28922), .IN2(n24443), .IN3(n28925), .IN4(n24447), .Q(
        n24429) );
  OA22X1 U27907 ( .IN1(n28926), .IN2(n24445), .IN3(n28924), .IN4(n24442), .Q(
        n24428) );
  NAND4X0 U27908 ( .IN1(n24431), .IN2(n24430), .IN3(n24429), .IN4(n24428), 
        .QN(s13_addr_o[29]) );
  OA22X1 U27909 ( .IN1(n28937), .IN2(n24432), .IN3(n28939), .IN4(n24446), .Q(
        n24439) );
  OA22X1 U27910 ( .IN1(n28935), .IN2(n24433), .IN3(n28931), .IN4(n24447), .Q(
        n24438) );
  OA22X1 U27911 ( .IN1(n28932), .IN2(n24434), .IN3(n28933), .IN4(n24444), .Q(
        n24437) );
  OA22X1 U27912 ( .IN1(n28936), .IN2(n24441), .IN3(n28940), .IN4(n24435), .Q(
        n24436) );
  NAND4X0 U27913 ( .IN1(n24439), .IN2(n24438), .IN3(n24437), .IN4(n24436), 
        .QN(s13_addr_o[30]) );
  OA22X1 U27914 ( .IN1(n28954), .IN2(n24441), .IN3(n28958), .IN4(n24440), .Q(
        n24451) );
  OA22X1 U27915 ( .IN1(n28956), .IN2(n24443), .IN3(n28952), .IN4(n24442), .Q(
        n24450) );
  OA22X1 U27916 ( .IN1(n28948), .IN2(n24445), .IN3(n28960), .IN4(n24444), .Q(
        n24449) );
  OA22X1 U27917 ( .IN1(n28950), .IN2(n24447), .IN3(n28946), .IN4(n24446), .Q(
        n24448) );
  NAND4X0 U27918 ( .IN1(n24451), .IN2(n24450), .IN3(n24449), .IN4(n24448), 
        .QN(s13_addr_o[31]) );
  OA22X1 U27919 ( .IN1(n29349), .IN2(n24453), .IN3(n29311), .IN4(n24452), .Q(
        n24464) );
  INVX0 U27920 ( .INP(n24454), .ZN(n24456) );
  OA22X1 U27921 ( .IN1(n29254), .IN2(n24456), .IN3(n29292), .IN4(n24455), .Q(
        n24463) );
  OA22X1 U27922 ( .IN1(n29273), .IN2(n24458), .IN3(n29330), .IN4(n24457), .Q(
        n24462) );
  OA22X1 U27923 ( .IN1(n29368), .IN2(n24460), .IN3(n29235), .IN4(n24459), .Q(
        n24461) );
  NAND4X0 U27924 ( .IN1(n24464), .IN2(n24463), .IN3(n24462), .IN4(n24461), 
        .QN(s12_stb_o) );
  INVX0 U27925 ( .INP(n29192), .ZN(n24748) );
  INVX0 U27926 ( .INP(n29184), .ZN(n24740) );
  OA22X1 U27927 ( .IN1(n24748), .IN2(n28123), .IN3(n24740), .IN4(n28126), .Q(
        n24468) );
  INVX0 U27928 ( .INP(n29191), .ZN(n24752) );
  INVX0 U27929 ( .INP(n29181), .ZN(n24731) );
  OA22X1 U27930 ( .IN1(n24752), .IN2(n28124), .IN3(n24731), .IN4(n28128), .Q(
        n24467) );
  INVX0 U27931 ( .INP(n29182), .ZN(n24736) );
  INVX0 U27932 ( .INP(n29189), .ZN(n24722) );
  OA22X1 U27933 ( .IN1(n24736), .IN2(n28122), .IN3(n24722), .IN4(n28125), .Q(
        n24466) );
  INVX0 U27934 ( .INP(n24738), .ZN(n29183) );
  INVX0 U27935 ( .INP(n29183), .ZN(n24746) );
  INVX0 U27936 ( .INP(n24701), .ZN(n29190) );
  INVX0 U27937 ( .INP(n29190), .ZN(n24745) );
  OA22X1 U27938 ( .IN1(n24746), .IN2(n28127), .IN3(n24745), .IN4(n28121), .Q(
        n24465) );
  NAND4X0 U27939 ( .IN1(n24468), .IN2(n24467), .IN3(n24466), .IN4(n24465), 
        .QN(s12_we_o) );
  OA22X1 U27940 ( .IN1(n24722), .IN2(n28136), .IN3(n24738), .IN4(n28137), .Q(
        n24472) );
  OA22X1 U27941 ( .IN1(n24752), .IN2(n28134), .IN3(n24740), .IN4(n28139), .Q(
        n24471) );
  OA22X1 U27942 ( .IN1(n24736), .IN2(n28138), .IN3(n24701), .IN4(n28135), .Q(
        n24470) );
  INVX0 U27943 ( .INP(n29192), .ZN(n24739) );
  OA22X1 U27944 ( .IN1(n24747), .IN2(n28140), .IN3(n24739), .IN4(n28133), .Q(
        n24469) );
  NAND4X0 U27945 ( .IN1(n24472), .IN2(n24471), .IN3(n24470), .IN4(n24469), 
        .QN(s12_data_o[0]) );
  INVX0 U27946 ( .INP(n29182), .ZN(n24751) );
  OA22X1 U27947 ( .IN1(n24751), .IN2(n28149), .IN3(n24701), .IN4(n28147), .Q(
        n24476) );
  OA22X1 U27948 ( .IN1(n24731), .IN2(n28146), .IN3(n24739), .IN4(n28148), .Q(
        n24475) );
  OA22X1 U27949 ( .IN1(n24737), .IN2(n28150), .IN3(n24722), .IN4(n28152), .Q(
        n24474) );
  OA22X1 U27950 ( .IN1(n24740), .IN2(n28145), .IN3(n24738), .IN4(n28151), .Q(
        n24473) );
  NAND4X0 U27951 ( .IN1(n24476), .IN2(n24475), .IN3(n24474), .IN4(n24473), 
        .QN(s12_data_o[1]) );
  OA22X1 U27952 ( .IN1(n24747), .IN2(n28164), .IN3(n24738), .IN4(n28157), .Q(
        n24480) );
  OA22X1 U27953 ( .IN1(n24737), .IN2(n28160), .IN3(n24722), .IN4(n28162), .Q(
        n24479) );
  OA22X1 U27954 ( .IN1(n24739), .IN2(n28163), .IN3(n24740), .IN4(n28159), .Q(
        n24478) );
  OA22X1 U27955 ( .IN1(n24751), .IN2(n28158), .IN3(n24701), .IN4(n28161), .Q(
        n24477) );
  NAND4X0 U27956 ( .IN1(n24480), .IN2(n24479), .IN3(n24478), .IN4(n24477), 
        .QN(s12_data_o[2]) );
  OA22X1 U27957 ( .IN1(n24737), .IN2(n28172), .IN3(n24736), .IN4(n28171), .Q(
        n24484) );
  OA22X1 U27958 ( .IN1(n24748), .IN2(n28176), .IN3(n24738), .IN4(n28169), .Q(
        n24483) );
  INVX0 U27959 ( .INP(n29184), .ZN(n24749) );
  OA22X1 U27960 ( .IN1(n24749), .IN2(n28170), .IN3(n24722), .IN4(n28175), .Q(
        n24482) );
  OA22X1 U27961 ( .IN1(n24731), .IN2(n28174), .IN3(n24701), .IN4(n28173), .Q(
        n24481) );
  NAND4X0 U27962 ( .IN1(n24484), .IN2(n24483), .IN3(n24482), .IN4(n24481), 
        .QN(s12_data_o[3]) );
  OA22X1 U27963 ( .IN1(n24747), .IN2(n28184), .IN3(n24701), .IN4(n28181), .Q(
        n24488) );
  OA22X1 U27964 ( .IN1(n24736), .IN2(n28185), .IN3(n24738), .IN4(n28187), .Q(
        n24487) );
  OA22X1 U27965 ( .IN1(n24740), .IN2(n28188), .IN3(n24722), .IN4(n28183), .Q(
        n24486) );
  OA22X1 U27966 ( .IN1(n24737), .IN2(n28182), .IN3(n24739), .IN4(n28186), .Q(
        n24485) );
  NAND4X0 U27967 ( .IN1(n24488), .IN2(n24487), .IN3(n24486), .IN4(n24485), 
        .QN(s12_data_o[4]) );
  OA22X1 U27968 ( .IN1(n24739), .IN2(n28194), .IN3(n24740), .IN4(n28193), .Q(
        n24492) );
  OA22X1 U27969 ( .IN1(n24747), .IN2(n28200), .IN3(n24701), .IN4(n28199), .Q(
        n24491) );
  OA22X1 U27970 ( .IN1(n24737), .IN2(n28196), .IN3(n24736), .IN4(n28198), .Q(
        n24490) );
  INVX0 U27971 ( .INP(n29189), .ZN(n24750) );
  OA22X1 U27972 ( .IN1(n24750), .IN2(n28197), .IN3(n24738), .IN4(n28195), .Q(
        n24489) );
  NAND4X0 U27973 ( .IN1(n24492), .IN2(n24491), .IN3(n24490), .IN4(n24489), 
        .QN(s12_data_o[5]) );
  OA22X1 U27974 ( .IN1(n24737), .IN2(n28208), .IN3(n24739), .IN4(n28206), .Q(
        n24496) );
  OA22X1 U27975 ( .IN1(n24751), .IN2(n28211), .IN3(n24701), .IN4(n28209), .Q(
        n24495) );
  OA22X1 U27976 ( .IN1(n24731), .IN2(n28207), .IN3(n24750), .IN4(n28205), .Q(
        n24494) );
  OA22X1 U27977 ( .IN1(n24749), .IN2(n28212), .IN3(n24738), .IN4(n28210), .Q(
        n24493) );
  NAND4X0 U27978 ( .IN1(n24496), .IN2(n24495), .IN3(n24494), .IN4(n24493), 
        .QN(s12_data_o[6]) );
  OA22X1 U27979 ( .IN1(n24737), .IN2(n28220), .IN3(n24731), .IN4(n28219), .Q(
        n24500) );
  OA22X1 U27980 ( .IN1(n24739), .IN2(n28224), .IN3(n24740), .IN4(n28218), .Q(
        n24499) );
  OA22X1 U27981 ( .IN1(n24736), .IN2(n28217), .IN3(n24745), .IN4(n28221), .Q(
        n24498) );
  OA22X1 U27982 ( .IN1(n24722), .IN2(n28223), .IN3(n24738), .IN4(n28222), .Q(
        n24497) );
  NAND4X0 U27983 ( .IN1(n24500), .IN2(n24499), .IN3(n24498), .IN4(n24497), 
        .QN(s12_data_o[7]) );
  OA22X1 U27984 ( .IN1(n24747), .IN2(n28232), .IN3(n24745), .IN4(n28235), .Q(
        n24504) );
  OA22X1 U27985 ( .IN1(n24736), .IN2(n28236), .IN3(n24722), .IN4(n28229), .Q(
        n24503) );
  OA22X1 U27986 ( .IN1(n24752), .IN2(n28230), .IN3(n24738), .IN4(n28233), .Q(
        n24502) );
  OA22X1 U27987 ( .IN1(n24739), .IN2(n28231), .IN3(n24740), .IN4(n28234), .Q(
        n24501) );
  NAND4X0 U27988 ( .IN1(n24504), .IN2(n24503), .IN3(n24502), .IN4(n24501), 
        .QN(s12_data_o[8]) );
  OA22X1 U27989 ( .IN1(n24740), .IN2(n28248), .IN3(n24745), .IN4(n28247), .Q(
        n24508) );
  OA22X1 U27990 ( .IN1(n24748), .IN2(n28246), .IN3(n24750), .IN4(n28245), .Q(
        n24507) );
  OA22X1 U27991 ( .IN1(n24731), .IN2(n28244), .IN3(n24736), .IN4(n28241), .Q(
        n24506) );
  OA22X1 U27992 ( .IN1(n24737), .IN2(n28242), .IN3(n24738), .IN4(n28243), .Q(
        n24505) );
  NAND4X0 U27993 ( .IN1(n24508), .IN2(n24507), .IN3(n24506), .IN4(n24505), 
        .QN(s12_data_o[9]) );
  OA22X1 U27994 ( .IN1(n24751), .IN2(n28254), .IN3(n24745), .IN4(n28259), .Q(
        n24512) );
  OA22X1 U27995 ( .IN1(n24749), .IN2(n28256), .IN3(n24746), .IN4(n28253), .Q(
        n24511) );
  OA22X1 U27996 ( .IN1(n24752), .IN2(n28258), .IN3(n24739), .IN4(n28260), .Q(
        n24510) );
  OA22X1 U27997 ( .IN1(n24747), .IN2(n28257), .IN3(n24750), .IN4(n28255), .Q(
        n24509) );
  NAND4X0 U27998 ( .IN1(n24512), .IN2(n24511), .IN3(n24510), .IN4(n24509), 
        .QN(s12_data_o[10]) );
  OA22X1 U27999 ( .IN1(n24748), .IN2(n28265), .IN3(n24745), .IN4(n28269), .Q(
        n24516) );
  OA22X1 U28000 ( .IN1(n24740), .IN2(n28271), .IN3(n24746), .IN4(n28267), .Q(
        n24515) );
  OA22X1 U28001 ( .IN1(n24737), .IN2(n28266), .IN3(n24731), .IN4(n28272), .Q(
        n24514) );
  OA22X1 U28002 ( .IN1(n24751), .IN2(n28268), .IN3(n24722), .IN4(n28270), .Q(
        n24513) );
  NAND4X0 U28003 ( .IN1(n24516), .IN2(n24515), .IN3(n24514), .IN4(n24513), 
        .QN(s12_data_o[11]) );
  OA22X1 U28004 ( .IN1(n24752), .IN2(n28284), .IN3(n24736), .IN4(n28283), .Q(
        n24520) );
  OA22X1 U28005 ( .IN1(n24750), .IN2(n28281), .IN3(n24745), .IN4(n28277), .Q(
        n24519) );
  OA22X1 U28006 ( .IN1(n24739), .IN2(n28280), .IN3(n24740), .IN4(n28282), .Q(
        n24518) );
  OA22X1 U28007 ( .IN1(n24747), .IN2(n28278), .IN3(n24746), .IN4(n28279), .Q(
        n24517) );
  NAND4X0 U28008 ( .IN1(n24520), .IN2(n24519), .IN3(n24518), .IN4(n24517), 
        .QN(s12_data_o[12]) );
  OA22X1 U28009 ( .IN1(n24747), .IN2(n28294), .IN3(n24739), .IN4(n28296), .Q(
        n24524) );
  OA22X1 U28010 ( .IN1(n24737), .IN2(n28290), .IN3(n24722), .IN4(n28293), .Q(
        n24523) );
  OA22X1 U28011 ( .IN1(n24751), .IN2(n28289), .IN3(n24746), .IN4(n28291), .Q(
        n24522) );
  OA22X1 U28012 ( .IN1(n24749), .IN2(n28292), .IN3(n24745), .IN4(n28295), .Q(
        n24521) );
  NAND4X0 U28013 ( .IN1(n24524), .IN2(n24523), .IN3(n24522), .IN4(n24521), 
        .QN(s12_data_o[13]) );
  OA22X1 U28014 ( .IN1(n24752), .IN2(n28306), .IN3(n24731), .IN4(n28304), .Q(
        n24528) );
  OA22X1 U28015 ( .IN1(n24739), .IN2(n28308), .IN3(n24745), .IN4(n28303), .Q(
        n24527) );
  OA22X1 U28016 ( .IN1(n24736), .IN2(n28307), .IN3(n24722), .IN4(n28302), .Q(
        n24526) );
  OA22X1 U28017 ( .IN1(n24749), .IN2(n28305), .IN3(n24746), .IN4(n28301), .Q(
        n24525) );
  NAND4X0 U28018 ( .IN1(n24528), .IN2(n24527), .IN3(n24526), .IN4(n24525), 
        .QN(s12_data_o[14]) );
  OA22X1 U28019 ( .IN1(n24747), .IN2(n28315), .IN3(n24739), .IN4(n28314), .Q(
        n24532) );
  OA22X1 U28020 ( .IN1(n24737), .IN2(n28316), .IN3(n24722), .IN4(n28318), .Q(
        n24531) );
  OA22X1 U28021 ( .IN1(n24738), .IN2(n28317), .IN3(n24745), .IN4(n28319), .Q(
        n24530) );
  OA22X1 U28022 ( .IN1(n24749), .IN2(n28313), .IN3(n24736), .IN4(n28320), .Q(
        n24529) );
  NAND4X0 U28023 ( .IN1(n24532), .IN2(n24531), .IN3(n24530), .IN4(n24529), 
        .QN(s12_data_o[15]) );
  OA22X1 U28024 ( .IN1(n24739), .IN2(n28331), .IN3(n24740), .IN4(n28326), .Q(
        n24536) );
  OA22X1 U28025 ( .IN1(n24738), .IN2(n28328), .IN3(n24745), .IN4(n28327), .Q(
        n24535) );
  OA22X1 U28026 ( .IN1(n24747), .IN2(n28332), .IN3(n24722), .IN4(n28325), .Q(
        n24534) );
  OA22X1 U28027 ( .IN1(n24752), .IN2(n28330), .IN3(n24751), .IN4(n28329), .Q(
        n24533) );
  NAND4X0 U28028 ( .IN1(n24536), .IN2(n24535), .IN3(n24534), .IN4(n24533), 
        .QN(s12_data_o[16]) );
  OA22X1 U28029 ( .IN1(n24737), .IN2(n28340), .IN3(n24731), .IN4(n28344), .Q(
        n24540) );
  OA22X1 U28030 ( .IN1(n24746), .IN2(n28343), .IN3(n24745), .IN4(n28341), .Q(
        n24539) );
  OA22X1 U28031 ( .IN1(n24748), .IN2(n28342), .IN3(n24740), .IN4(n28338), .Q(
        n24538) );
  OA22X1 U28032 ( .IN1(n24751), .IN2(n28337), .IN3(n24722), .IN4(n28339), .Q(
        n24537) );
  NAND4X0 U28033 ( .IN1(n24540), .IN2(n24539), .IN3(n24538), .IN4(n24537), 
        .QN(s12_data_o[17]) );
  OA22X1 U28034 ( .IN1(n24749), .IN2(n28355), .IN3(n24722), .IN4(n28349), .Q(
        n24544) );
  OA22X1 U28035 ( .IN1(n24747), .IN2(n28356), .IN3(n24746), .IN4(n28351), .Q(
        n24543) );
  OA22X1 U28036 ( .IN1(n24736), .IN2(n28354), .IN3(n24745), .IN4(n28353), .Q(
        n24542) );
  OA22X1 U28037 ( .IN1(n24752), .IN2(n28352), .IN3(n24739), .IN4(n28350), .Q(
        n24541) );
  NAND4X0 U28038 ( .IN1(n24544), .IN2(n24543), .IN3(n24542), .IN4(n24541), 
        .QN(s12_data_o[18]) );
  OA22X1 U28039 ( .IN1(n24747), .IN2(n28364), .IN3(n24746), .IN4(n28368), .Q(
        n24548) );
  OA22X1 U28040 ( .IN1(n24752), .IN2(n28366), .IN3(n24722), .IN4(n28361), .Q(
        n24547) );
  OA22X1 U28041 ( .IN1(n24748), .IN2(n28362), .IN3(n24749), .IN4(n28363), .Q(
        n24546) );
  OA22X1 U28042 ( .IN1(n24751), .IN2(n28365), .IN3(n24745), .IN4(n28367), .Q(
        n24545) );
  NAND4X0 U28043 ( .IN1(n24548), .IN2(n24547), .IN3(n24546), .IN4(n24545), 
        .QN(s12_data_o[19]) );
  OA22X1 U28044 ( .IN1(n24739), .IN2(n28374), .IN3(n24746), .IN4(n28379), .Q(
        n24552) );
  OA22X1 U28045 ( .IN1(n24737), .IN2(n28378), .IN3(n24731), .IN4(n28377), .Q(
        n24551) );
  OA22X1 U28046 ( .IN1(n24749), .IN2(n28373), .IN3(n24736), .IN4(n28376), .Q(
        n24550) );
  OA22X1 U28047 ( .IN1(n24722), .IN2(n28380), .IN3(n24745), .IN4(n28375), .Q(
        n24549) );
  NAND4X0 U28048 ( .IN1(n24552), .IN2(n24551), .IN3(n24550), .IN4(n24549), 
        .QN(s12_data_o[20]) );
  OA22X1 U28049 ( .IN1(n24752), .IN2(n28392), .IN3(n24739), .IN4(n28390), .Q(
        n24556) );
  OA22X1 U28050 ( .IN1(n24747), .IN2(n28386), .IN3(n24740), .IN4(n28388), .Q(
        n24555) );
  OA22X1 U28051 ( .IN1(n24736), .IN2(n28387), .IN3(n24722), .IN4(n28385), .Q(
        n24554) );
  OA22X1 U28052 ( .IN1(n24738), .IN2(n28389), .IN3(n24745), .IN4(n28391), .Q(
        n24553) );
  NAND4X0 U28053 ( .IN1(n24556), .IN2(n24555), .IN3(n24554), .IN4(n24553), 
        .QN(s12_data_o[21]) );
  OA22X1 U28054 ( .IN1(n24739), .IN2(n28404), .IN3(n24745), .IN4(n28397), .Q(
        n24560) );
  OA22X1 U28055 ( .IN1(n24747), .IN2(n28402), .IN3(n24722), .IN4(n28399), .Q(
        n24559) );
  OA22X1 U28056 ( .IN1(n24749), .IN2(n28403), .IN3(n24751), .IN4(n28398), .Q(
        n24558) );
  OA22X1 U28057 ( .IN1(n24752), .IN2(n28400), .IN3(n24746), .IN4(n28401), .Q(
        n24557) );
  NAND4X0 U28058 ( .IN1(n24560), .IN2(n24559), .IN3(n24558), .IN4(n24557), 
        .QN(s12_data_o[22]) );
  OA22X1 U28059 ( .IN1(n24752), .IN2(n28416), .IN3(n24750), .IN4(n28412), .Q(
        n24564) );
  OA22X1 U28060 ( .IN1(n24749), .IN2(n28413), .IN3(n24701), .IN4(n28411), .Q(
        n24563) );
  OA22X1 U28061 ( .IN1(n24751), .IN2(n28410), .IN3(n24746), .IN4(n28409), .Q(
        n24562) );
  OA22X1 U28062 ( .IN1(n24747), .IN2(n28415), .IN3(n24748), .IN4(n28414), .Q(
        n24561) );
  NAND4X0 U28063 ( .IN1(n24564), .IN2(n24563), .IN3(n24562), .IN4(n24561), 
        .QN(s12_data_o[23]) );
  OA22X1 U28064 ( .IN1(n24746), .IN2(n28427), .IN3(n24701), .IN4(n28423), .Q(
        n24568) );
  OA22X1 U28065 ( .IN1(n24747), .IN2(n28424), .IN3(n24736), .IN4(n28425), .Q(
        n24567) );
  OA22X1 U28066 ( .IN1(n24752), .IN2(n28426), .IN3(n24749), .IN4(n28421), .Q(
        n24566) );
  OA22X1 U28067 ( .IN1(n24739), .IN2(n28422), .IN3(n24722), .IN4(n28428), .Q(
        n24565) );
  NAND4X0 U28068 ( .IN1(n24568), .IN2(n24567), .IN3(n24566), .IN4(n24565), 
        .QN(s12_data_o[24]) );
  OA22X1 U28069 ( .IN1(n24747), .IN2(n28440), .IN3(n24749), .IN4(n28439), .Q(
        n24572) );
  OA22X1 U28070 ( .IN1(n24752), .IN2(n28438), .IN3(n24722), .IN4(n28437), .Q(
        n24571) );
  OA22X1 U28071 ( .IN1(n24739), .IN2(n28434), .IN3(n24746), .IN4(n28436), .Q(
        n24570) );
  OA22X1 U28072 ( .IN1(n24736), .IN2(n28433), .IN3(n24701), .IN4(n28435), .Q(
        n24569) );
  NAND4X0 U28073 ( .IN1(n24572), .IN2(n24571), .IN3(n24570), .IN4(n24569), 
        .QN(s12_data_o[25]) );
  OA22X1 U28074 ( .IN1(n24752), .IN2(n28452), .IN3(n24731), .IN4(n28451), .Q(
        n24576) );
  OA22X1 U28075 ( .IN1(n24736), .IN2(n28449), .IN3(n24701), .IN4(n28445), .Q(
        n24575) );
  OA22X1 U28076 ( .IN1(n24750), .IN2(n28448), .IN3(n24746), .IN4(n28447), .Q(
        n24574) );
  OA22X1 U28077 ( .IN1(n24748), .IN2(n28450), .IN3(n24740), .IN4(n28446), .Q(
        n24573) );
  NAND4X0 U28078 ( .IN1(n24576), .IN2(n24575), .IN3(n24574), .IN4(n24573), 
        .QN(s12_data_o[26]) );
  OA22X1 U28079 ( .IN1(n24749), .IN2(n28458), .IN3(n24701), .IN4(n28459), .Q(
        n24580) );
  OA22X1 U28080 ( .IN1(n24752), .IN2(n28462), .IN3(n24748), .IN4(n28464), .Q(
        n24579) );
  OA22X1 U28081 ( .IN1(n24736), .IN2(n28457), .IN3(n24746), .IN4(n28460), .Q(
        n24578) );
  OA22X1 U28082 ( .IN1(n24747), .IN2(n28461), .IN3(n24722), .IN4(n28463), .Q(
        n24577) );
  NAND4X0 U28083 ( .IN1(n24580), .IN2(n24579), .IN3(n24578), .IN4(n24577), 
        .QN(s12_data_o[27]) );
  OA22X1 U28084 ( .IN1(n24748), .IN2(n28472), .IN3(n24740), .IN4(n28470), .Q(
        n24584) );
  OA22X1 U28085 ( .IN1(n24752), .IN2(n28474), .IN3(n24701), .IN4(n28473), .Q(
        n24583) );
  OA22X1 U28086 ( .IN1(n24722), .IN2(n28475), .IN3(n24746), .IN4(n28469), .Q(
        n24582) );
  OA22X1 U28087 ( .IN1(n24747), .IN2(n28476), .IN3(n24751), .IN4(n28471), .Q(
        n24581) );
  NAND4X0 U28088 ( .IN1(n24584), .IN2(n24583), .IN3(n24582), .IN4(n24581), 
        .QN(s12_data_o[28]) );
  OA22X1 U28089 ( .IN1(n24736), .IN2(n28487), .IN3(n24750), .IN4(n28483), .Q(
        n24588) );
  OA22X1 U28090 ( .IN1(n24731), .IN2(n28482), .IN3(n24746), .IN4(n28485), .Q(
        n24587) );
  OA22X1 U28091 ( .IN1(n24752), .IN2(n28484), .IN3(n24749), .IN4(n28486), .Q(
        n24586) );
  OA22X1 U28092 ( .IN1(n24748), .IN2(n28488), .IN3(n24701), .IN4(n28481), .Q(
        n24585) );
  NAND4X0 U28093 ( .IN1(n24588), .IN2(n24587), .IN3(n24586), .IN4(n24585), 
        .QN(s12_data_o[29]) );
  OA22X1 U28094 ( .IN1(n24740), .IN2(n28496), .IN3(n24751), .IN4(n28493), .Q(
        n24592) );
  OA22X1 U28095 ( .IN1(n24738), .IN2(n28500), .IN3(n24701), .IN4(n28499), .Q(
        n24591) );
  OA22X1 U28096 ( .IN1(n24739), .IN2(n28497), .IN3(n24722), .IN4(n28495), .Q(
        n24590) );
  OA22X1 U28097 ( .IN1(n24752), .IN2(n28494), .IN3(n24731), .IN4(n28498), .Q(
        n24589) );
  NAND4X0 U28098 ( .IN1(n24592), .IN2(n24591), .IN3(n24590), .IN4(n24589), 
        .QN(s12_data_o[30]) );
  OA22X1 U28099 ( .IN1(n24752), .IN2(n28510), .IN3(n24739), .IN4(n28506), .Q(
        n24596) );
  OA22X1 U28100 ( .IN1(n24738), .IN2(n28511), .IN3(n24701), .IN4(n28507), .Q(
        n24595) );
  OA22X1 U28101 ( .IN1(n24731), .IN2(n28509), .IN3(n24751), .IN4(n28512), .Q(
        n24594) );
  OA22X1 U28102 ( .IN1(n24740), .IN2(n28505), .IN3(n24750), .IN4(n28508), .Q(
        n24593) );
  NAND4X0 U28103 ( .IN1(n24596), .IN2(n24595), .IN3(n24594), .IN4(n24593), 
        .QN(s12_data_o[31]) );
  OA22X1 U28104 ( .IN1(n24752), .IN2(n28518), .IN3(n24739), .IN4(n28522), .Q(
        n24600) );
  OA22X1 U28105 ( .IN1(n24738), .IN2(n28521), .IN3(n24701), .IN4(n28519), .Q(
        n24599) );
  OA22X1 U28106 ( .IN1(n24751), .IN2(n28523), .IN3(n24722), .IN4(n28520), .Q(
        n24598) );
  OA22X1 U28107 ( .IN1(n24731), .IN2(n28517), .IN3(n24740), .IN4(n28524), .Q(
        n24597) );
  NAND4X0 U28108 ( .IN1(n24600), .IN2(n24599), .IN3(n24598), .IN4(n24597), 
        .QN(s12_sel_o[0]) );
  OA22X1 U28109 ( .IN1(n24740), .IN2(n28536), .IN3(n24746), .IN4(n28531), .Q(
        n24604) );
  OA22X1 U28110 ( .IN1(n24750), .IN2(n28533), .IN3(n24701), .IN4(n28529), .Q(
        n24603) );
  OA22X1 U28111 ( .IN1(n24731), .IN2(n28532), .IN3(n24751), .IN4(n28535), .Q(
        n24602) );
  OA22X1 U28112 ( .IN1(n24752), .IN2(n28534), .IN3(n24739), .IN4(n28530), .Q(
        n24601) );
  NAND4X0 U28113 ( .IN1(n24604), .IN2(n24603), .IN3(n24602), .IN4(n24601), 
        .QN(s12_sel_o[1]) );
  OA22X1 U28114 ( .IN1(n24752), .IN2(n28544), .IN3(n24701), .IN4(n28541), .Q(
        n24608) );
  OA22X1 U28115 ( .IN1(n24731), .IN2(n28546), .IN3(n24750), .IN4(n28542), .Q(
        n24607) );
  OA22X1 U28116 ( .IN1(n24736), .IN2(n28547), .IN3(n24738), .IN4(n28545), .Q(
        n24606) );
  OA22X1 U28117 ( .IN1(n24748), .IN2(n28543), .IN3(n24740), .IN4(n28548), .Q(
        n24605) );
  NAND4X0 U28118 ( .IN1(n24608), .IN2(n24607), .IN3(n24606), .IN4(n24605), 
        .QN(s12_sel_o[2]) );
  OA22X1 U28119 ( .IN1(n24731), .IN2(n28554), .IN3(n24738), .IN4(n28559), .Q(
        n24612) );
  OA22X1 U28120 ( .IN1(n24739), .IN2(n28553), .IN3(n24751), .IN4(n28556), .Q(
        n24611) );
  OA22X1 U28121 ( .IN1(n24737), .IN2(n28558), .IN3(n24749), .IN4(n28557), .Q(
        n24610) );
  OA22X1 U28122 ( .IN1(n24750), .IN2(n28560), .IN3(n24701), .IN4(n28555), .Q(
        n24609) );
  NAND4X0 U28123 ( .IN1(n24612), .IN2(n24611), .IN3(n24610), .IN4(n24609), 
        .QN(s12_sel_o[3]) );
  OA22X1 U28124 ( .IN1(n24738), .IN2(n28565), .IN3(n24701), .IN4(n28569), .Q(
        n24616) );
  OA22X1 U28125 ( .IN1(n24731), .IN2(n28570), .IN3(n24751), .IN4(n28568), .Q(
        n24615) );
  OA22X1 U28126 ( .IN1(n24737), .IN2(n28572), .IN3(n24750), .IN4(n28567), .Q(
        n24614) );
  OA22X1 U28127 ( .IN1(n24748), .IN2(n28571), .IN3(n24740), .IN4(n28566), .Q(
        n24613) );
  NAND4X0 U28128 ( .IN1(n24616), .IN2(n24615), .IN3(n24614), .IN4(n24613), 
        .QN(s12_addr_o[0]) );
  OA22X1 U28129 ( .IN1(n24747), .IN2(n28578), .IN3(n24739), .IN4(n28582), .Q(
        n24620) );
  OA22X1 U28130 ( .IN1(n24750), .IN2(n28584), .IN3(n24701), .IN4(n28583), .Q(
        n24619) );
  OA22X1 U28131 ( .IN1(n24737), .IN2(n28580), .IN3(n24738), .IN4(n28577), .Q(
        n24618) );
  OA22X1 U28132 ( .IN1(n24740), .IN2(n28581), .IN3(n24751), .IN4(n28579), .Q(
        n24617) );
  NAND4X0 U28133 ( .IN1(n24620), .IN2(n24619), .IN3(n24618), .IN4(n24617), 
        .QN(s12_addr_o[1]) );
  OA22X1 U28134 ( .IN1(n28596), .IN2(n24745), .IN3(n28594), .IN4(n24739), .Q(
        n24624) );
  OA22X1 U28135 ( .IN1(n28589), .IN2(n24747), .IN3(n28595), .IN4(n24738), .Q(
        n24623) );
  OA22X1 U28136 ( .IN1(n28592), .IN2(n24740), .IN3(n28593), .IN4(n24722), .Q(
        n24622) );
  OA22X1 U28137 ( .IN1(n28591), .IN2(n24752), .IN3(n28590), .IN4(n24751), .Q(
        n24621) );
  NAND4X0 U28138 ( .IN1(n24624), .IN2(n24623), .IN3(n24622), .IN4(n24621), 
        .QN(s12_addr_o[2]) );
  OA22X1 U28139 ( .IN1(n28605), .IN2(n24731), .IN3(n28607), .IN4(n24740), .Q(
        n24628) );
  OA22X1 U28140 ( .IN1(n28603), .IN2(n24746), .IN3(n28608), .IN4(n24745), .Q(
        n24627) );
  OA22X1 U28141 ( .IN1(n28602), .IN2(n24750), .IN3(n28606), .IN4(n24751), .Q(
        n24626) );
  OA22X1 U28142 ( .IN1(n28604), .IN2(n24739), .IN3(n28601), .IN4(n24737), .Q(
        n24625) );
  NAND4X0 U28143 ( .IN1(n24628), .IN2(n24627), .IN3(n24626), .IN4(n24625), 
        .QN(s12_addr_o[3]) );
  OA22X1 U28144 ( .IN1(n28617), .IN2(n24752), .IN3(n28615), .IN4(n24751), .Q(
        n24632) );
  OA22X1 U28145 ( .IN1(n28616), .IN2(n24747), .IN3(n28613), .IN4(n24748), .Q(
        n24631) );
  OA22X1 U28146 ( .IN1(n28620), .IN2(n24746), .IN3(n28619), .IN4(n24745), .Q(
        n24630) );
  OA22X1 U28147 ( .IN1(n28618), .IN2(n24749), .IN3(n28614), .IN4(n24750), .Q(
        n24629) );
  NAND4X0 U28148 ( .IN1(n24632), .IN2(n24631), .IN3(n24630), .IN4(n24629), 
        .QN(s12_addr_o[4]) );
  OA22X1 U28149 ( .IN1(n28627), .IN2(n24750), .IN3(n28625), .IN4(n24745), .Q(
        n24636) );
  OA22X1 U28150 ( .IN1(n28628), .IN2(n24746), .IN3(n28631), .IN4(n24751), .Q(
        n24635) );
  OA22X1 U28151 ( .IN1(n28626), .IN2(n24740), .IN3(n28630), .IN4(n24731), .Q(
        n24634) );
  OA22X1 U28152 ( .IN1(n28632), .IN2(n24748), .IN3(n28629), .IN4(n24737), .Q(
        n24633) );
  NAND4X0 U28153 ( .IN1(n24636), .IN2(n24635), .IN3(n24634), .IN4(n24633), 
        .QN(s12_addr_o[5]) );
  OA22X1 U28154 ( .IN1(n24747), .IN2(n28640), .IN3(n24722), .IN4(n28637), .Q(
        n24640) );
  OA22X1 U28155 ( .IN1(n24748), .IN2(n28644), .IN3(n24701), .IN4(n28639), .Q(
        n24639) );
  OA22X1 U28156 ( .IN1(n24737), .IN2(n28642), .IN3(n24738), .IN4(n28641), .Q(
        n24638) );
  OA22X1 U28157 ( .IN1(n24749), .IN2(n28643), .IN3(n24751), .IN4(n28638), .Q(
        n24637) );
  NAND4X0 U28158 ( .IN1(n24640), .IN2(n24639), .IN3(n24638), .IN4(n24637), 
        .QN(s12_addr_o[6]) );
  OA22X1 U28159 ( .IN1(n24736), .IN2(n28650), .IN3(n24701), .IN4(n28655), .Q(
        n24644) );
  OA22X1 U28160 ( .IN1(n24748), .IN2(n28656), .IN3(n24738), .IN4(n28651), .Q(
        n24643) );
  OA22X1 U28161 ( .IN1(n24737), .IN2(n28654), .IN3(n24731), .IN4(n28652), .Q(
        n24642) );
  OA22X1 U28162 ( .IN1(n24749), .IN2(n28653), .IN3(n24750), .IN4(n28649), .Q(
        n24641) );
  NAND4X0 U28163 ( .IN1(n24644), .IN2(n24643), .IN3(n24642), .IN4(n24641), 
        .QN(s12_addr_o[7]) );
  OA22X1 U28164 ( .IN1(n24731), .IN2(n28663), .IN3(n24751), .IN4(n28668), .Q(
        n24648) );
  OA22X1 U28165 ( .IN1(n24750), .IN2(n28662), .IN3(n24701), .IN4(n28667), .Q(
        n24647) );
  OA22X1 U28166 ( .IN1(n24748), .IN2(n28666), .IN3(n24749), .IN4(n28665), .Q(
        n24646) );
  OA22X1 U28167 ( .IN1(n24752), .IN2(n28664), .IN3(n24738), .IN4(n28661), .Q(
        n24645) );
  NAND4X0 U28168 ( .IN1(n24648), .IN2(n24647), .IN3(n24646), .IN4(n24645), 
        .QN(s12_addr_o[8]) );
  OA22X1 U28169 ( .IN1(n24731), .IN2(n28679), .IN3(n24749), .IN4(n28676), .Q(
        n24652) );
  OA22X1 U28170 ( .IN1(n24748), .IN2(n28674), .IN3(n24701), .IN4(n28677), .Q(
        n24651) );
  OA22X1 U28171 ( .IN1(n24736), .IN2(n28673), .IN3(n24738), .IN4(n28675), .Q(
        n24650) );
  OA22X1 U28172 ( .IN1(n24752), .IN2(n28680), .IN3(n24750), .IN4(n28678), .Q(
        n24649) );
  NAND4X0 U28173 ( .IN1(n24652), .IN2(n24651), .IN3(n24650), .IN4(n24649), 
        .QN(s12_addr_o[9]) );
  OA22X1 U28174 ( .IN1(n24737), .IN2(n28692), .IN3(n24739), .IN4(n28688), .Q(
        n24656) );
  OA22X1 U28175 ( .IN1(n24749), .IN2(n28687), .IN3(n24722), .IN4(n28691), .Q(
        n24655) );
  OA22X1 U28176 ( .IN1(n24731), .IN2(n28686), .IN3(n24738), .IN4(n28690), .Q(
        n24654) );
  OA22X1 U28177 ( .IN1(n24736), .IN2(n28685), .IN3(n24701), .IN4(n28689), .Q(
        n24653) );
  NAND4X0 U28178 ( .IN1(n24656), .IN2(n24655), .IN3(n24654), .IN4(n24653), 
        .QN(s12_addr_o[10]) );
  OA22X1 U28179 ( .IN1(n24748), .IN2(n28697), .IN3(n24738), .IN4(n28700), .Q(
        n24660) );
  OA22X1 U28180 ( .IN1(n24751), .IN2(n28701), .IN3(n24701), .IN4(n28699), .Q(
        n24659) );
  OA22X1 U28181 ( .IN1(n24749), .IN2(n28704), .IN3(n24722), .IN4(n28703), .Q(
        n24658) );
  OA22X1 U28182 ( .IN1(n24737), .IN2(n28702), .IN3(n24731), .IN4(n28698), .Q(
        n24657) );
  NAND4X0 U28183 ( .IN1(n24660), .IN2(n24659), .IN3(n24658), .IN4(n24657), 
        .QN(s12_addr_o[11]) );
  OA22X1 U28184 ( .IN1(n24752), .IN2(n28714), .IN3(n24731), .IN4(n28710), .Q(
        n24664) );
  OA22X1 U28185 ( .IN1(n24748), .IN2(n28712), .IN3(n24740), .IN4(n28716), .Q(
        n24663) );
  OA22X1 U28186 ( .IN1(n24736), .IN2(n28709), .IN3(n24750), .IN4(n28715), .Q(
        n24662) );
  OA22X1 U28187 ( .IN1(n24746), .IN2(n28711), .IN3(n24701), .IN4(n28713), .Q(
        n24661) );
  NAND4X0 U28188 ( .IN1(n24664), .IN2(n24663), .IN3(n24662), .IN4(n24661), 
        .QN(s12_addr_o[12]) );
  OA22X1 U28189 ( .IN1(n24747), .IN2(n28728), .IN3(n24740), .IN4(n28724), .Q(
        n24668) );
  OA22X1 U28190 ( .IN1(n24748), .IN2(n28726), .IN3(n24738), .IN4(n28725), .Q(
        n24667) );
  OA22X1 U28191 ( .IN1(n24736), .IN2(n28723), .IN3(n24701), .IN4(n28727), .Q(
        n24666) );
  OA22X1 U28192 ( .IN1(n24752), .IN2(n28722), .IN3(n24722), .IN4(n28721), .Q(
        n24665) );
  NAND4X0 U28193 ( .IN1(n24668), .IN2(n24667), .IN3(n24666), .IN4(n24665), 
        .QN(s12_addr_o[13]) );
  OA22X1 U28194 ( .IN1(n24737), .IN2(n28734), .IN3(n24701), .IN4(n28739), .Q(
        n24672) );
  OA22X1 U28195 ( .IN1(n24748), .IN2(n28736), .IN3(n24749), .IN4(n28735), .Q(
        n24671) );
  OA22X1 U28196 ( .IN1(n24750), .IN2(n28737), .IN3(n24738), .IN4(n28733), .Q(
        n24670) );
  OA22X1 U28197 ( .IN1(n24747), .IN2(n28738), .IN3(n24736), .IN4(n28740), .Q(
        n24669) );
  NAND4X0 U28198 ( .IN1(n24672), .IN2(n24671), .IN3(n24670), .IN4(n24669), 
        .QN(s12_addr_o[14]) );
  OA22X1 U28199 ( .IN1(n24752), .IN2(n28746), .IN3(n24751), .IN4(n28747), .Q(
        n24676) );
  OA22X1 U28200 ( .IN1(n24747), .IN2(n28748), .IN3(n24701), .IN4(n28745), .Q(
        n24675) );
  OA22X1 U28201 ( .IN1(n24749), .IN2(n28752), .IN3(n24738), .IN4(n28749), .Q(
        n24674) );
  OA22X1 U28202 ( .IN1(n24748), .IN2(n28750), .IN3(n24722), .IN4(n28751), .Q(
        n24673) );
  NAND4X0 U28203 ( .IN1(n24676), .IN2(n24675), .IN3(n24674), .IN4(n24673), 
        .QN(s12_addr_o[15]) );
  OA22X1 U28204 ( .IN1(n24731), .IN2(n28762), .IN3(n24736), .IN4(n28759), .Q(
        n24680) );
  OA22X1 U28205 ( .IN1(n24738), .IN2(n28764), .IN3(n24701), .IN4(n28763), .Q(
        n24679) );
  OA22X1 U28206 ( .IN1(n24737), .IN2(n28758), .IN3(n24740), .IN4(n28761), .Q(
        n24678) );
  OA22X1 U28207 ( .IN1(n24748), .IN2(n28760), .IN3(n24750), .IN4(n28757), .Q(
        n24677) );
  NAND4X0 U28208 ( .IN1(n24680), .IN2(n24679), .IN3(n24678), .IN4(n24677), 
        .QN(s12_addr_o[16]) );
  OA22X1 U28209 ( .IN1(n24748), .IN2(n28774), .IN3(n24701), .IN4(n28769), .Q(
        n24684) );
  OA22X1 U28210 ( .IN1(n24749), .IN2(n28773), .IN3(n24751), .IN4(n28775), .Q(
        n24683) );
  OA22X1 U28211 ( .IN1(n24752), .IN2(n28772), .IN3(n24738), .IN4(n28770), .Q(
        n24682) );
  OA22X1 U28212 ( .IN1(n24747), .IN2(n28776), .IN3(n24750), .IN4(n28771), .Q(
        n24681) );
  NAND4X0 U28213 ( .IN1(n24684), .IN2(n24683), .IN3(n24682), .IN4(n24681), 
        .QN(s12_addr_o[17]) );
  OA22X1 U28214 ( .IN1(n24752), .IN2(n28786), .IN3(n24739), .IN4(n28787), .Q(
        n24688) );
  OA22X1 U28215 ( .IN1(n24749), .IN2(n28782), .IN3(n24736), .IN4(n28784), .Q(
        n24687) );
  OA22X1 U28216 ( .IN1(n24731), .IN2(n28788), .IN3(n24701), .IN4(n28781), .Q(
        n24686) );
  OA22X1 U28217 ( .IN1(n24750), .IN2(n28783), .IN3(n24738), .IN4(n28785), .Q(
        n24685) );
  NAND4X0 U28218 ( .IN1(n24688), .IN2(n24687), .IN3(n24686), .IN4(n24685), 
        .QN(s12_addr_o[18]) );
  OA22X1 U28219 ( .IN1(n24748), .IN2(n28798), .IN3(n24701), .IN4(n28799), .Q(
        n24692) );
  OA22X1 U28220 ( .IN1(n24750), .IN2(n28795), .IN3(n24738), .IN4(n28793), .Q(
        n24691) );
  OA22X1 U28221 ( .IN1(n24731), .IN2(n28800), .IN3(n24749), .IN4(n28794), .Q(
        n24690) );
  OA22X1 U28222 ( .IN1(n24737), .IN2(n28796), .IN3(n24751), .IN4(n28797), .Q(
        n24689) );
  NAND4X0 U28223 ( .IN1(n24692), .IN2(n24691), .IN3(n24690), .IN4(n24689), 
        .QN(s12_addr_o[19]) );
  OA22X1 U28224 ( .IN1(n24748), .IN2(n28807), .IN3(n24701), .IN4(n28805), .Q(
        n24696) );
  OA22X1 U28225 ( .IN1(n24751), .IN2(n28806), .IN3(n24722), .IN4(n28811), .Q(
        n24695) );
  OA22X1 U28226 ( .IN1(n24737), .IN2(n28812), .IN3(n24749), .IN4(n28810), .Q(
        n24694) );
  OA22X1 U28227 ( .IN1(n24747), .IN2(n28808), .IN3(n24738), .IN4(n28809), .Q(
        n24693) );
  NAND4X0 U28228 ( .IN1(n24696), .IN2(n24695), .IN3(n24694), .IN4(n24693), 
        .QN(s12_addr_o[20]) );
  OA22X1 U28229 ( .IN1(n24747), .IN2(n28824), .IN3(n24740), .IN4(n28819), .Q(
        n24700) );
  OA22X1 U28230 ( .IN1(n24737), .IN2(n28822), .IN3(n24738), .IN4(n28818), .Q(
        n24699) );
  OA22X1 U28231 ( .IN1(n24739), .IN2(n28820), .IN3(n24722), .IN4(n28823), .Q(
        n24698) );
  OA22X1 U28232 ( .IN1(n24736), .IN2(n28821), .IN3(n24701), .IN4(n28817), .Q(
        n24697) );
  NAND4X0 U28233 ( .IN1(n24700), .IN2(n24699), .IN3(n24698), .IN4(n24697), 
        .QN(s12_addr_o[21]) );
  OA22X1 U28234 ( .IN1(n24731), .IN2(n28832), .IN3(n24722), .IN4(n28834), .Q(
        n24705) );
  OA22X1 U28235 ( .IN1(n24752), .IN2(n28833), .IN3(n24736), .IN4(n28836), .Q(
        n24704) );
  OA22X1 U28236 ( .IN1(n24748), .IN2(n28831), .IN3(n24738), .IN4(n28837), .Q(
        n24703) );
  OA22X1 U28237 ( .IN1(n24749), .IN2(n28838), .IN3(n24701), .IN4(n28829), .Q(
        n24702) );
  NAND4X0 U28238 ( .IN1(n24705), .IN2(n24704), .IN3(n24703), .IN4(n24702), 
        .QN(s12_addr_o[22]) );
  OA22X1 U28239 ( .IN1(n24731), .IN2(n28845), .IN3(n24751), .IN4(n28852), .Q(
        n24709) );
  OA22X1 U28240 ( .IN1(n24748), .IN2(n28843), .IN3(n24740), .IN4(n28850), .Q(
        n24708) );
  OA22X1 U28241 ( .IN1(n24737), .IN2(n28848), .IN3(n24745), .IN4(n28851), .Q(
        n24707) );
  OA22X1 U28242 ( .IN1(n24750), .IN2(n28849), .IN3(n24738), .IN4(n28846), .Q(
        n24706) );
  NAND4X0 U28243 ( .IN1(n24709), .IN2(n24708), .IN3(n24707), .IN4(n24706), 
        .QN(s12_addr_o[23]) );
  OA22X1 U28244 ( .IN1(n28865), .IN2(n24746), .IN3(n28864), .IN4(n24747), .Q(
        n24713) );
  OA22X1 U28245 ( .IN1(n28858), .IN2(n24739), .IN3(n28860), .IN4(n24745), .Q(
        n24712) );
  OA22X1 U28246 ( .IN1(n28857), .IN2(n24749), .IN3(n28861), .IN4(n24751), .Q(
        n24711) );
  OA22X1 U28247 ( .IN1(n28859), .IN2(n24750), .IN3(n28863), .IN4(n24737), .Q(
        n24710) );
  NAND4X0 U28248 ( .IN1(n24713), .IN2(n24712), .IN3(n24711), .IN4(n24710), 
        .QN(s12_addr_o[24]) );
  OA22X1 U28249 ( .IN1(n28877), .IN2(n24731), .IN3(n28872), .IN4(n24736), .Q(
        n24717) );
  OA22X1 U28250 ( .IN1(n28870), .IN2(n24737), .IN3(n28874), .IN4(n24749), .Q(
        n24716) );
  OA22X1 U28251 ( .IN1(n28875), .IN2(n24745), .IN3(n28876), .IN4(n24722), .Q(
        n24715) );
  OA22X1 U28252 ( .IN1(n28873), .IN2(n24748), .IN3(n28871), .IN4(n24738), .Q(
        n24714) );
  NAND4X0 U28253 ( .IN1(n24717), .IN2(n24716), .IN3(n24715), .IN4(n24714), 
        .QN(s12_addr_o[25]) );
  OA22X1 U28254 ( .IN1(n28885), .IN2(n24739), .IN3(n28882), .IN4(n24749), .Q(
        n24721) );
  OA22X1 U28255 ( .IN1(n28889), .IN2(n24745), .IN3(n28888), .IN4(n24750), .Q(
        n24720) );
  OA22X1 U28256 ( .IN1(n28884), .IN2(n24752), .IN3(n28886), .IN4(n24736), .Q(
        n24719) );
  OA22X1 U28257 ( .IN1(n28883), .IN2(n24746), .IN3(n28887), .IN4(n24731), .Q(
        n24718) );
  NAND4X0 U28258 ( .IN1(n24721), .IN2(n24720), .IN3(n24719), .IN4(n24718), 
        .QN(s12_addr_o[26]) );
  OA22X1 U28259 ( .IN1(n28897), .IN2(n24746), .IN3(n28895), .IN4(n24747), .Q(
        n24726) );
  OA22X1 U28260 ( .IN1(n28898), .IN2(n24745), .IN3(n28901), .IN4(n24740), .Q(
        n24725) );
  OA22X1 U28261 ( .IN1(n28894), .IN2(n24737), .IN3(n28900), .IN4(n24736), .Q(
        n24724) );
  OA22X1 U28262 ( .IN1(n28899), .IN2(n24748), .IN3(n28896), .IN4(n24722), .Q(
        n24723) );
  NAND4X0 U28263 ( .IN1(n24726), .IN2(n24725), .IN3(n24724), .IN4(n24723), 
        .QN(s12_addr_o[27]) );
  OA22X1 U28264 ( .IN1(n28907), .IN2(n24746), .IN3(n28912), .IN4(n24737), .Q(
        n24730) );
  OA22X1 U28265 ( .IN1(n28913), .IN2(n24745), .IN3(n28910), .IN4(n24750), .Q(
        n24729) );
  OA22X1 U28266 ( .IN1(n28909), .IN2(n24739), .IN3(n28911), .IN4(n24731), .Q(
        n24728) );
  OA22X1 U28267 ( .IN1(n28908), .IN2(n24740), .IN3(n28906), .IN4(n24751), .Q(
        n24727) );
  NAND4X0 U28268 ( .IN1(n24730), .IN2(n24729), .IN3(n24728), .IN4(n24727), 
        .QN(s12_addr_o[28]) );
  OA22X1 U28269 ( .IN1(n28922), .IN2(n24746), .IN3(n28925), .IN4(n24737), .Q(
        n24735) );
  OA22X1 U28270 ( .IN1(n28924), .IN2(n24731), .IN3(n28919), .IN4(n24740), .Q(
        n24734) );
  OA22X1 U28271 ( .IN1(n28920), .IN2(n24750), .IN3(n28923), .IN4(n24751), .Q(
        n24733) );
  OA22X1 U28272 ( .IN1(n28926), .IN2(n24748), .IN3(n28921), .IN4(n24745), .Q(
        n24732) );
  NAND4X0 U28273 ( .IN1(n24735), .IN2(n24734), .IN3(n24733), .IN4(n24732), 
        .QN(s12_addr_o[29]) );
  OA22X1 U28274 ( .IN1(n28931), .IN2(n24737), .IN3(n28939), .IN4(n24736), .Q(
        n24744) );
  OA22X1 U28275 ( .IN1(n28932), .IN2(n24739), .IN3(n28937), .IN4(n24738), .Q(
        n24743) );
  OA22X1 U28276 ( .IN1(n28936), .IN2(n24750), .IN3(n28940), .IN4(n24740), .Q(
        n24742) );
  OA22X1 U28277 ( .IN1(n28935), .IN2(n24747), .IN3(n28933), .IN4(n24745), .Q(
        n24741) );
  NAND4X0 U28278 ( .IN1(n24744), .IN2(n24743), .IN3(n24742), .IN4(n24741), 
        .QN(s12_addr_o[30]) );
  OA22X1 U28279 ( .IN1(n28956), .IN2(n24746), .IN3(n28960), .IN4(n24745), .Q(
        n24756) );
  OA22X1 U28280 ( .IN1(n28948), .IN2(n24748), .IN3(n28952), .IN4(n24747), .Q(
        n24755) );
  OA22X1 U28281 ( .IN1(n28954), .IN2(n24750), .IN3(n28958), .IN4(n24749), .Q(
        n24754) );
  OA22X1 U28282 ( .IN1(n28950), .IN2(n24752), .IN3(n28946), .IN4(n24751), .Q(
        n24753) );
  NAND4X0 U28283 ( .IN1(n24756), .IN2(n24755), .IN3(n24754), .IN4(n24753), 
        .QN(s12_addr_o[31]) );
  OA22X1 U28284 ( .IN1(n29349), .IN2(n24758), .IN3(n29254), .IN4(n24757), .Q(
        n24769) );
  INVX0 U28285 ( .INP(n24759), .ZN(n24761) );
  OA22X1 U28286 ( .IN1(n29235), .IN2(n24761), .IN3(n29311), .IN4(n24760), .Q(
        n24768) );
  OA22X1 U28287 ( .IN1(n29368), .IN2(n24763), .IN3(n29292), .IN4(n24762), .Q(
        n24767) );
  OA22X1 U28288 ( .IN1(n29273), .IN2(n24765), .IN3(n29330), .IN4(n24764), .Q(
        n24766) );
  NAND4X0 U28289 ( .IN1(n24769), .IN2(n24768), .IN3(n24767), .IN4(n24766), 
        .QN(s11_stb_o) );
  INVX0 U28290 ( .INP(n29166), .ZN(n25028) );
  INVX0 U28291 ( .INP(n29172), .ZN(n25050) );
  OA22X1 U28292 ( .IN1(n25028), .IN2(n28126), .IN3(n25050), .IN4(n28122), .Q(
        n24773) );
  INVX0 U28293 ( .INP(n29163), .ZN(n25055) );
  INVX0 U28294 ( .INP(n29164), .ZN(n25011) );
  OA22X1 U28295 ( .IN1(n25055), .IN2(n28128), .IN3(n25011), .IN4(n28123), .Q(
        n24772) );
  INVX0 U28296 ( .INP(n29171), .ZN(n25056) );
  INVX0 U28297 ( .INP(n25006), .ZN(n29174) );
  INVX0 U28298 ( .INP(n29174), .ZN(n25051) );
  OA22X1 U28299 ( .IN1(n25056), .IN2(n28127), .IN3(n25051), .IN4(n28121), .Q(
        n24771) );
  INVX0 U28300 ( .INP(n29165), .ZN(n25038) );
  INVX0 U28301 ( .INP(n29173), .ZN(n25054) );
  OA22X1 U28302 ( .IN1(n25038), .IN2(n28124), .IN3(n25054), .IN4(n28125), .Q(
        n24770) );
  NAND4X0 U28303 ( .IN1(n24773), .IN2(n24772), .IN3(n24771), .IN4(n24770), 
        .QN(s11_we_o) );
  OA22X1 U28304 ( .IN1(n25055), .IN2(n28140), .IN3(n25050), .IN4(n28138), .Q(
        n24777) );
  OA22X1 U28305 ( .IN1(n25054), .IN2(n28136), .IN3(n25056), .IN4(n28137), .Q(
        n24776) );
  OA22X1 U28306 ( .IN1(n25038), .IN2(n28134), .IN3(n25011), .IN4(n28133), .Q(
        n24775) );
  OA22X1 U28307 ( .IN1(n25028), .IN2(n28139), .IN3(n25006), .IN4(n28135), .Q(
        n24774) );
  NAND4X0 U28308 ( .IN1(n24777), .IN2(n24776), .IN3(n24775), .IN4(n24774), 
        .QN(s11_data_o[0]) );
  INVX0 U28309 ( .INP(n29173), .ZN(n25039) );
  OA22X1 U28310 ( .IN1(n25039), .IN2(n28152), .IN3(n25006), .IN4(n28147), .Q(
        n24781) );
  OA22X1 U28311 ( .IN1(n25055), .IN2(n28146), .IN3(n25050), .IN4(n28149), .Q(
        n24780) );
  INVX0 U28312 ( .INP(n29166), .ZN(n25052) );
  INVX0 U28313 ( .INP(n29171), .ZN(n25045) );
  OA22X1 U28314 ( .IN1(n25052), .IN2(n28145), .IN3(n25045), .IN4(n28151), .Q(
        n24779) );
  OA22X1 U28315 ( .IN1(n25038), .IN2(n28150), .IN3(n25011), .IN4(n28148), .Q(
        n24778) );
  NAND4X0 U28316 ( .IN1(n24781), .IN2(n24780), .IN3(n24779), .IN4(n24778), 
        .QN(s11_data_o[1]) );
  INVX0 U28317 ( .INP(n29164), .ZN(n25057) );
  OA22X1 U28318 ( .IN1(n25057), .IN2(n28163), .IN3(n25052), .IN4(n28159), .Q(
        n24785) );
  OA22X1 U28319 ( .IN1(n25055), .IN2(n28164), .IN3(n25050), .IN4(n28158), .Q(
        n24784) );
  OA22X1 U28320 ( .IN1(n25054), .IN2(n28162), .IN3(n25045), .IN4(n28157), .Q(
        n24783) );
  OA22X1 U28321 ( .IN1(n25038), .IN2(n28160), .IN3(n25006), .IN4(n28161), .Q(
        n24782) );
  NAND4X0 U28322 ( .IN1(n24785), .IN2(n24784), .IN3(n24783), .IN4(n24782), 
        .QN(s11_data_o[2]) );
  OA22X1 U28323 ( .IN1(n25050), .IN2(n28171), .IN3(n25045), .IN4(n28169), .Q(
        n24789) );
  OA22X1 U28324 ( .IN1(n25038), .IN2(n28172), .IN3(n25011), .IN4(n28176), .Q(
        n24788) );
  OA22X1 U28325 ( .IN1(n25039), .IN2(n28175), .IN3(n25006), .IN4(n28173), .Q(
        n24787) );
  OA22X1 U28326 ( .IN1(n25055), .IN2(n28174), .IN3(n25052), .IN4(n28170), .Q(
        n24786) );
  NAND4X0 U28327 ( .IN1(n24789), .IN2(n24788), .IN3(n24787), .IN4(n24786), 
        .QN(s11_data_o[3]) );
  OA22X1 U28328 ( .IN1(n25011), .IN2(n28186), .IN3(n25052), .IN4(n28188), .Q(
        n24793) );
  INVX0 U28329 ( .INP(n29172), .ZN(n25029) );
  OA22X1 U28330 ( .IN1(n25029), .IN2(n28185), .IN3(n25006), .IN4(n28181), .Q(
        n24792) );
  OA22X1 U28331 ( .IN1(n25054), .IN2(n28183), .IN3(n25045), .IN4(n28187), .Q(
        n24791) );
  OA22X1 U28332 ( .IN1(n25038), .IN2(n28182), .IN3(n25044), .IN4(n28184), .Q(
        n24790) );
  NAND4X0 U28333 ( .IN1(n24793), .IN2(n24792), .IN3(n24791), .IN4(n24790), 
        .QN(s11_data_o[4]) );
  OA22X1 U28334 ( .IN1(n25039), .IN2(n28197), .IN3(n25006), .IN4(n28199), .Q(
        n24797) );
  OA22X1 U28335 ( .IN1(n25052), .IN2(n28193), .IN3(n25029), .IN4(n28198), .Q(
        n24796) );
  OA22X1 U28336 ( .IN1(n25055), .IN2(n28200), .IN3(n25045), .IN4(n28195), .Q(
        n24795) );
  OA22X1 U28337 ( .IN1(n25053), .IN2(n28196), .IN3(n25011), .IN4(n28194), .Q(
        n24794) );
  NAND4X0 U28338 ( .IN1(n24797), .IN2(n24796), .IN3(n24795), .IN4(n24794), 
        .QN(s11_data_o[5]) );
  OA22X1 U28339 ( .IN1(n25011), .IN2(n28206), .IN3(n25045), .IN4(n28210), .Q(
        n24801) );
  OA22X1 U28340 ( .IN1(n25028), .IN2(n28212), .IN3(n25050), .IN4(n28211), .Q(
        n24800) );
  OA22X1 U28341 ( .IN1(n25044), .IN2(n28207), .IN3(n25006), .IN4(n28209), .Q(
        n24799) );
  OA22X1 U28342 ( .IN1(n25038), .IN2(n28208), .IN3(n25039), .IN4(n28205), .Q(
        n24798) );
  NAND4X0 U28343 ( .IN1(n24801), .IN2(n24800), .IN3(n24799), .IN4(n24798), 
        .QN(s11_data_o[6]) );
  OA22X1 U28344 ( .IN1(n25055), .IN2(n28219), .IN3(n25029), .IN4(n28217), .Q(
        n24805) );
  OA22X1 U28345 ( .IN1(n25053), .IN2(n28220), .IN3(n25051), .IN4(n28221), .Q(
        n24804) );
  OA22X1 U28346 ( .IN1(n25028), .IN2(n28218), .IN3(n25045), .IN4(n28222), .Q(
        n24803) );
  OA22X1 U28347 ( .IN1(n25011), .IN2(n28224), .IN3(n25039), .IN4(n28223), .Q(
        n24802) );
  NAND4X0 U28348 ( .IN1(n24805), .IN2(n24804), .IN3(n24803), .IN4(n24802), 
        .QN(s11_data_o[7]) );
  OA22X1 U28349 ( .IN1(n25054), .IN2(n28229), .IN3(n25051), .IN4(n28235), .Q(
        n24809) );
  OA22X1 U28350 ( .IN1(n25050), .IN2(n28236), .IN3(n25045), .IN4(n28233), .Q(
        n24808) );
  OA22X1 U28351 ( .IN1(n25038), .IN2(n28230), .IN3(n25044), .IN4(n28232), .Q(
        n24807) );
  OA22X1 U28352 ( .IN1(n25011), .IN2(n28231), .IN3(n25052), .IN4(n28234), .Q(
        n24806) );
  NAND4X0 U28353 ( .IN1(n24809), .IN2(n24808), .IN3(n24807), .IN4(n24806), 
        .QN(s11_data_o[8]) );
  OA22X1 U28354 ( .IN1(n25029), .IN2(n28241), .IN3(n25056), .IN4(n28243), .Q(
        n24813) );
  OA22X1 U28355 ( .IN1(n25054), .IN2(n28245), .IN3(n25051), .IN4(n28247), .Q(
        n24812) );
  OA22X1 U28356 ( .IN1(n25053), .IN2(n28242), .IN3(n25011), .IN4(n28246), .Q(
        n24811) );
  OA22X1 U28357 ( .IN1(n25055), .IN2(n28244), .IN3(n25052), .IN4(n28248), .Q(
        n24810) );
  NAND4X0 U28358 ( .IN1(n24813), .IN2(n24812), .IN3(n24811), .IN4(n24810), 
        .QN(s11_data_o[9]) );
  OA22X1 U28359 ( .IN1(n25038), .IN2(n28258), .IN3(n25056), .IN4(n28253), .Q(
        n24817) );
  OA22X1 U28360 ( .IN1(n25052), .IN2(n28256), .IN3(n25051), .IN4(n28259), .Q(
        n24816) );
  OA22X1 U28361 ( .IN1(n25011), .IN2(n28260), .IN3(n25039), .IN4(n28255), .Q(
        n24815) );
  OA22X1 U28362 ( .IN1(n25055), .IN2(n28257), .IN3(n25050), .IN4(n28254), .Q(
        n24814) );
  NAND4X0 U28363 ( .IN1(n24817), .IN2(n24816), .IN3(n24815), .IN4(n24814), 
        .QN(s11_data_o[10]) );
  OA22X1 U28364 ( .IN1(n25054), .IN2(n28270), .IN3(n25056), .IN4(n28267), .Q(
        n24821) );
  OA22X1 U28365 ( .IN1(n25053), .IN2(n28266), .IN3(n25011), .IN4(n28265), .Q(
        n24820) );
  OA22X1 U28366 ( .IN1(n25028), .IN2(n28271), .IN3(n25050), .IN4(n28268), .Q(
        n24819) );
  OA22X1 U28367 ( .IN1(n25055), .IN2(n28272), .IN3(n25051), .IN4(n28269), .Q(
        n24818) );
  NAND4X0 U28368 ( .IN1(n24821), .IN2(n24820), .IN3(n24819), .IN4(n24818), 
        .QN(s11_data_o[11]) );
  OA22X1 U28369 ( .IN1(n25057), .IN2(n28280), .IN3(n25050), .IN4(n28283), .Q(
        n24825) );
  OA22X1 U28370 ( .IN1(n25038), .IN2(n28284), .IN3(n25039), .IN4(n28281), .Q(
        n24824) );
  OA22X1 U28371 ( .IN1(n25055), .IN2(n28278), .IN3(n25052), .IN4(n28282), .Q(
        n24823) );
  OA22X1 U28372 ( .IN1(n25045), .IN2(n28279), .IN3(n25051), .IN4(n28277), .Q(
        n24822) );
  NAND4X0 U28373 ( .IN1(n24825), .IN2(n24824), .IN3(n24823), .IN4(n24822), 
        .QN(s11_data_o[12]) );
  OA22X1 U28374 ( .IN1(n25055), .IN2(n28294), .IN3(n25056), .IN4(n28291), .Q(
        n24829) );
  OA22X1 U28375 ( .IN1(n25011), .IN2(n28296), .IN3(n25052), .IN4(n28292), .Q(
        n24828) );
  OA22X1 U28376 ( .IN1(n25053), .IN2(n28290), .IN3(n25051), .IN4(n28295), .Q(
        n24827) );
  OA22X1 U28377 ( .IN1(n25050), .IN2(n28289), .IN3(n25039), .IN4(n28293), .Q(
        n24826) );
  NAND4X0 U28378 ( .IN1(n24829), .IN2(n24828), .IN3(n24827), .IN4(n24826), 
        .QN(s11_data_o[13]) );
  OA22X1 U28379 ( .IN1(n25055), .IN2(n28304), .IN3(n25039), .IN4(n28302), .Q(
        n24833) );
  OA22X1 U28380 ( .IN1(n25057), .IN2(n28308), .IN3(n25051), .IN4(n28303), .Q(
        n24832) );
  OA22X1 U28381 ( .IN1(n25052), .IN2(n28305), .IN3(n25056), .IN4(n28301), .Q(
        n24831) );
  OA22X1 U28382 ( .IN1(n25038), .IN2(n28306), .IN3(n25050), .IN4(n28307), .Q(
        n24830) );
  NAND4X0 U28383 ( .IN1(n24833), .IN2(n24832), .IN3(n24831), .IN4(n24830), 
        .QN(s11_data_o[14]) );
  OA22X1 U28384 ( .IN1(n25055), .IN2(n28315), .IN3(n25056), .IN4(n28317), .Q(
        n24837) );
  OA22X1 U28385 ( .IN1(n25053), .IN2(n28316), .IN3(n25039), .IN4(n28318), .Q(
        n24836) );
  OA22X1 U28386 ( .IN1(n25052), .IN2(n28313), .IN3(n25051), .IN4(n28319), .Q(
        n24835) );
  OA22X1 U28387 ( .IN1(n25057), .IN2(n28314), .IN3(n25050), .IN4(n28320), .Q(
        n24834) );
  NAND4X0 U28388 ( .IN1(n24837), .IN2(n24836), .IN3(n24835), .IN4(n24834), 
        .QN(s11_data_o[15]) );
  OA22X1 U28389 ( .IN1(n25029), .IN2(n28329), .IN3(n25051), .IN4(n28327), .Q(
        n24841) );
  OA22X1 U28390 ( .IN1(n25038), .IN2(n28330), .IN3(n25056), .IN4(n28328), .Q(
        n24840) );
  OA22X1 U28391 ( .IN1(n25011), .IN2(n28331), .IN3(n25052), .IN4(n28326), .Q(
        n24839) );
  OA22X1 U28392 ( .IN1(n25044), .IN2(n28332), .IN3(n25039), .IN4(n28325), .Q(
        n24838) );
  NAND4X0 U28393 ( .IN1(n24841), .IN2(n24840), .IN3(n24839), .IN4(n24838), 
        .QN(s11_data_o[16]) );
  OA22X1 U28394 ( .IN1(n25053), .IN2(n28340), .IN3(n25044), .IN4(n28344), .Q(
        n24845) );
  OA22X1 U28395 ( .IN1(n25054), .IN2(n28339), .IN3(n25056), .IN4(n28343), .Q(
        n24844) );
  OA22X1 U28396 ( .IN1(n25028), .IN2(n28338), .IN3(n25050), .IN4(n28337), .Q(
        n24843) );
  OA22X1 U28397 ( .IN1(n25057), .IN2(n28342), .IN3(n25051), .IN4(n28341), .Q(
        n24842) );
  NAND4X0 U28398 ( .IN1(n24845), .IN2(n24844), .IN3(n24843), .IN4(n24842), 
        .QN(s11_data_o[17]) );
  OA22X1 U28399 ( .IN1(n25055), .IN2(n28356), .IN3(n25029), .IN4(n28354), .Q(
        n24849) );
  OA22X1 U28400 ( .IN1(n25038), .IN2(n28352), .IN3(n25056), .IN4(n28351), .Q(
        n24848) );
  OA22X1 U28401 ( .IN1(n25054), .IN2(n28349), .IN3(n25051), .IN4(n28353), .Q(
        n24847) );
  OA22X1 U28402 ( .IN1(n25057), .IN2(n28350), .IN3(n25028), .IN4(n28355), .Q(
        n24846) );
  NAND4X0 U28403 ( .IN1(n24849), .IN2(n24848), .IN3(n24847), .IN4(n24846), 
        .QN(s11_data_o[18]) );
  OA22X1 U28404 ( .IN1(n25053), .IN2(n28366), .IN3(n25039), .IN4(n28361), .Q(
        n24853) );
  OA22X1 U28405 ( .IN1(n25056), .IN2(n28368), .IN3(n25051), .IN4(n28367), .Q(
        n24852) );
  OA22X1 U28406 ( .IN1(n25011), .IN2(n28362), .IN3(n25050), .IN4(n28365), .Q(
        n24851) );
  OA22X1 U28407 ( .IN1(n25055), .IN2(n28364), .IN3(n25028), .IN4(n28363), .Q(
        n24850) );
  NAND4X0 U28408 ( .IN1(n24853), .IN2(n24852), .IN3(n24851), .IN4(n24850), 
        .QN(s11_data_o[19]) );
  OA22X1 U28409 ( .IN1(n25054), .IN2(n28380), .IN3(n25056), .IN4(n28379), .Q(
        n24857) );
  OA22X1 U28410 ( .IN1(n25055), .IN2(n28377), .IN3(n25057), .IN4(n28374), .Q(
        n24856) );
  OA22X1 U28411 ( .IN1(n25052), .IN2(n28373), .IN3(n25029), .IN4(n28376), .Q(
        n24855) );
  OA22X1 U28412 ( .IN1(n25053), .IN2(n28378), .IN3(n25051), .IN4(n28375), .Q(
        n24854) );
  NAND4X0 U28413 ( .IN1(n24857), .IN2(n24856), .IN3(n24855), .IN4(n24854), 
        .QN(s11_data_o[20]) );
  OA22X1 U28414 ( .IN1(n25053), .IN2(n28392), .IN3(n25051), .IN4(n28391), .Q(
        n24861) );
  OA22X1 U28415 ( .IN1(n25011), .IN2(n28390), .IN3(n25039), .IN4(n28385), .Q(
        n24860) );
  OA22X1 U28416 ( .IN1(n25028), .IN2(n28388), .IN3(n25056), .IN4(n28389), .Q(
        n24859) );
  OA22X1 U28417 ( .IN1(n25044), .IN2(n28386), .IN3(n25029), .IN4(n28387), .Q(
        n24858) );
  NAND4X0 U28418 ( .IN1(n24861), .IN2(n24860), .IN3(n24859), .IN4(n24858), 
        .QN(s11_data_o[21]) );
  OA22X1 U28419 ( .IN1(n25053), .IN2(n28400), .IN3(n25028), .IN4(n28403), .Q(
        n24865) );
  OA22X1 U28420 ( .IN1(n25057), .IN2(n28404), .IN3(n25056), .IN4(n28401), .Q(
        n24864) );
  OA22X1 U28421 ( .IN1(n25050), .IN2(n28398), .IN3(n25039), .IN4(n28399), .Q(
        n24863) );
  OA22X1 U28422 ( .IN1(n25055), .IN2(n28402), .IN3(n25051), .IN4(n28397), .Q(
        n24862) );
  NAND4X0 U28423 ( .IN1(n24865), .IN2(n24864), .IN3(n24863), .IN4(n24862), 
        .QN(s11_data_o[22]) );
  OA22X1 U28424 ( .IN1(n25053), .IN2(n28416), .IN3(n25044), .IN4(n28415), .Q(
        n24869) );
  OA22X1 U28425 ( .IN1(n25052), .IN2(n28413), .IN3(n25006), .IN4(n28411), .Q(
        n24868) );
  OA22X1 U28426 ( .IN1(n25011), .IN2(n28414), .IN3(n25039), .IN4(n28412), .Q(
        n24867) );
  OA22X1 U28427 ( .IN1(n25029), .IN2(n28410), .IN3(n25056), .IN4(n28409), .Q(
        n24866) );
  NAND4X0 U28428 ( .IN1(n24869), .IN2(n24868), .IN3(n24867), .IN4(n24866), 
        .QN(s11_data_o[23]) );
  OA22X1 U28429 ( .IN1(n25028), .IN2(n28421), .IN3(n25006), .IN4(n28423), .Q(
        n24873) );
  OA22X1 U28430 ( .IN1(n25044), .IN2(n28424), .IN3(n25050), .IN4(n28425), .Q(
        n24872) );
  OA22X1 U28431 ( .IN1(n25053), .IN2(n28426), .IN3(n25039), .IN4(n28428), .Q(
        n24871) );
  OA22X1 U28432 ( .IN1(n25057), .IN2(n28422), .IN3(n25056), .IN4(n28427), .Q(
        n24870) );
  NAND4X0 U28433 ( .IN1(n24873), .IN2(n24872), .IN3(n24871), .IN4(n24870), 
        .QN(s11_data_o[24]) );
  OA22X1 U28434 ( .IN1(n25029), .IN2(n28433), .IN3(n25006), .IN4(n28435), .Q(
        n24877) );
  OA22X1 U28435 ( .IN1(n25053), .IN2(n28438), .IN3(n25044), .IN4(n28440), .Q(
        n24876) );
  OA22X1 U28436 ( .IN1(n25052), .IN2(n28439), .IN3(n25056), .IN4(n28436), .Q(
        n24875) );
  OA22X1 U28437 ( .IN1(n25057), .IN2(n28434), .IN3(n25054), .IN4(n28437), .Q(
        n24874) );
  NAND4X0 U28438 ( .IN1(n24877), .IN2(n24876), .IN3(n24875), .IN4(n24874), 
        .QN(s11_data_o[25]) );
  OA22X1 U28439 ( .IN1(n25053), .IN2(n28452), .IN3(n25056), .IN4(n28447), .Q(
        n24881) );
  OA22X1 U28440 ( .IN1(n25055), .IN2(n28451), .IN3(n25057), .IN4(n28450), .Q(
        n24880) );
  OA22X1 U28441 ( .IN1(n25028), .IN2(n28446), .IN3(n25029), .IN4(n28449), .Q(
        n24879) );
  OA22X1 U28442 ( .IN1(n25054), .IN2(n28448), .IN3(n25006), .IN4(n28445), .Q(
        n24878) );
  NAND4X0 U28443 ( .IN1(n24881), .IN2(n24880), .IN3(n24879), .IN4(n24878), 
        .QN(s11_data_o[26]) );
  OA22X1 U28444 ( .IN1(n25053), .IN2(n28462), .IN3(n25044), .IN4(n28461), .Q(
        n24885) );
  OA22X1 U28445 ( .IN1(n25054), .IN2(n28463), .IN3(n25006), .IN4(n28459), .Q(
        n24884) );
  OA22X1 U28446 ( .IN1(n25011), .IN2(n28464), .IN3(n25050), .IN4(n28457), .Q(
        n24883) );
  OA22X1 U28447 ( .IN1(n25052), .IN2(n28458), .IN3(n25045), .IN4(n28460), .Q(
        n24882) );
  NAND4X0 U28448 ( .IN1(n24885), .IN2(n24884), .IN3(n24883), .IN4(n24882), 
        .QN(s11_data_o[27]) );
  OA22X1 U28449 ( .IN1(n25053), .IN2(n28474), .IN3(n25052), .IN4(n28470), .Q(
        n24889) );
  OA22X1 U28450 ( .IN1(n25029), .IN2(n28471), .IN3(n25045), .IN4(n28469), .Q(
        n24888) );
  OA22X1 U28451 ( .IN1(n25044), .IN2(n28476), .IN3(n25054), .IN4(n28475), .Q(
        n24887) );
  OA22X1 U28452 ( .IN1(n25057), .IN2(n28472), .IN3(n25006), .IN4(n28473), .Q(
        n24886) );
  NAND4X0 U28453 ( .IN1(n24889), .IN2(n24888), .IN3(n24887), .IN4(n24886), 
        .QN(s11_data_o[28]) );
  OA22X1 U28454 ( .IN1(n25029), .IN2(n28487), .IN3(n25045), .IN4(n28485), .Q(
        n24893) );
  OA22X1 U28455 ( .IN1(n25055), .IN2(n28482), .IN3(n25052), .IN4(n28486), .Q(
        n24892) );
  OA22X1 U28456 ( .IN1(n25053), .IN2(n28484), .IN3(n25011), .IN4(n28488), .Q(
        n24891) );
  OA22X1 U28457 ( .IN1(n25054), .IN2(n28483), .IN3(n25006), .IN4(n28481), .Q(
        n24890) );
  NAND4X0 U28458 ( .IN1(n24893), .IN2(n24892), .IN3(n24891), .IN4(n24890), 
        .QN(s11_data_o[29]) );
  OA22X1 U28459 ( .IN1(n25044), .IN2(n28498), .IN3(n25057), .IN4(n28497), .Q(
        n24897) );
  OA22X1 U28460 ( .IN1(n25053), .IN2(n28494), .IN3(n25006), .IN4(n28499), .Q(
        n24896) );
  OA22X1 U28461 ( .IN1(n25029), .IN2(n28493), .IN3(n25045), .IN4(n28500), .Q(
        n24895) );
  OA22X1 U28462 ( .IN1(n25028), .IN2(n28496), .IN3(n25039), .IN4(n28495), .Q(
        n24894) );
  NAND4X0 U28463 ( .IN1(n24897), .IN2(n24896), .IN3(n24895), .IN4(n24894), 
        .QN(s11_data_o[30]) );
  OA22X1 U28464 ( .IN1(n25029), .IN2(n28512), .IN3(n25045), .IN4(n28511), .Q(
        n24901) );
  OA22X1 U28465 ( .IN1(n25052), .IN2(n28505), .IN3(n25006), .IN4(n28507), .Q(
        n24900) );
  OA22X1 U28466 ( .IN1(n25055), .IN2(n28509), .IN3(n25011), .IN4(n28506), .Q(
        n24899) );
  OA22X1 U28467 ( .IN1(n25053), .IN2(n28510), .IN3(n25039), .IN4(n28508), .Q(
        n24898) );
  NAND4X0 U28468 ( .IN1(n24901), .IN2(n24900), .IN3(n24899), .IN4(n24898), 
        .QN(s11_data_o[31]) );
  OA22X1 U28469 ( .IN1(n25011), .IN2(n28522), .IN3(n25028), .IN4(n28524), .Q(
        n24905) );
  OA22X1 U28470 ( .IN1(n25039), .IN2(n28520), .IN3(n25006), .IN4(n28519), .Q(
        n24904) );
  OA22X1 U28471 ( .IN1(n25053), .IN2(n28518), .IN3(n25050), .IN4(n28523), .Q(
        n24903) );
  OA22X1 U28472 ( .IN1(n25044), .IN2(n28517), .IN3(n25045), .IN4(n28521), .Q(
        n24902) );
  NAND4X0 U28473 ( .IN1(n24905), .IN2(n24904), .IN3(n24903), .IN4(n24902), 
        .QN(s11_sel_o[0]) );
  OA22X1 U28474 ( .IN1(n25044), .IN2(n28532), .IN3(n25045), .IN4(n28531), .Q(
        n24909) );
  OA22X1 U28475 ( .IN1(n25053), .IN2(n28534), .IN3(n25028), .IN4(n28536), .Q(
        n24908) );
  OA22X1 U28476 ( .IN1(n25057), .IN2(n28530), .IN3(n25006), .IN4(n28529), .Q(
        n24907) );
  OA22X1 U28477 ( .IN1(n25029), .IN2(n28535), .IN3(n25054), .IN4(n28533), .Q(
        n24906) );
  NAND4X0 U28478 ( .IN1(n24909), .IN2(n24908), .IN3(n24907), .IN4(n24906), 
        .QN(s11_sel_o[1]) );
  OA22X1 U28479 ( .IN1(n25056), .IN2(n28545), .IN3(n25006), .IN4(n28541), .Q(
        n24913) );
  OA22X1 U28480 ( .IN1(n25028), .IN2(n28548), .IN3(n25039), .IN4(n28542), .Q(
        n24912) );
  OA22X1 U28481 ( .IN1(n25044), .IN2(n28546), .IN3(n25029), .IN4(n28547), .Q(
        n24911) );
  OA22X1 U28482 ( .IN1(n25038), .IN2(n28544), .IN3(n25011), .IN4(n28543), .Q(
        n24910) );
  NAND4X0 U28483 ( .IN1(n24913), .IN2(n24912), .IN3(n24911), .IN4(n24910), 
        .QN(s11_sel_o[2]) );
  OA22X1 U28484 ( .IN1(n25044), .IN2(n28554), .IN3(n25057), .IN4(n28553), .Q(
        n24917) );
  OA22X1 U28485 ( .IN1(n25052), .IN2(n28557), .IN3(n25029), .IN4(n28556), .Q(
        n24916) );
  OA22X1 U28486 ( .IN1(n25038), .IN2(n28558), .IN3(n25045), .IN4(n28559), .Q(
        n24915) );
  OA22X1 U28487 ( .IN1(n25054), .IN2(n28560), .IN3(n25006), .IN4(n28555), .Q(
        n24914) );
  NAND4X0 U28488 ( .IN1(n24917), .IN2(n24916), .IN3(n24915), .IN4(n24914), 
        .QN(s11_sel_o[3]) );
  OA22X1 U28489 ( .IN1(n25011), .IN2(n28571), .IN3(n25006), .IN4(n28569), .Q(
        n24921) );
  OA22X1 U28490 ( .IN1(n25044), .IN2(n28570), .IN3(n25054), .IN4(n28567), .Q(
        n24920) );
  OA22X1 U28491 ( .IN1(n25028), .IN2(n28566), .IN3(n25050), .IN4(n28568), .Q(
        n24919) );
  OA22X1 U28492 ( .IN1(n25038), .IN2(n28572), .IN3(n25045), .IN4(n28565), .Q(
        n24918) );
  NAND4X0 U28493 ( .IN1(n24921), .IN2(n24920), .IN3(n24919), .IN4(n24918), 
        .QN(s11_addr_o[0]) );
  OA22X1 U28494 ( .IN1(n25038), .IN2(n28580), .IN3(n25045), .IN4(n28577), .Q(
        n24925) );
  OA22X1 U28495 ( .IN1(n25044), .IN2(n28578), .IN3(n25054), .IN4(n28584), .Q(
        n24924) );
  OA22X1 U28496 ( .IN1(n25029), .IN2(n28579), .IN3(n25006), .IN4(n28583), .Q(
        n24923) );
  OA22X1 U28497 ( .IN1(n25057), .IN2(n28582), .IN3(n25052), .IN4(n28581), .Q(
        n24922) );
  NAND4X0 U28498 ( .IN1(n24925), .IN2(n24924), .IN3(n24923), .IN4(n24922), 
        .QN(s11_addr_o[1]) );
  OA22X1 U28499 ( .IN1(n28590), .IN2(n25029), .IN3(n28593), .IN4(n25039), .Q(
        n24929) );
  OA22X1 U28500 ( .IN1(n28592), .IN2(n25028), .IN3(n28589), .IN4(n25055), .Q(
        n24928) );
  OA22X1 U28501 ( .IN1(n28591), .IN2(n25038), .IN3(n28594), .IN4(n25011), .Q(
        n24927) );
  OA22X1 U28502 ( .IN1(n28596), .IN2(n25051), .IN3(n28595), .IN4(n25045), .Q(
        n24926) );
  NAND4X0 U28503 ( .IN1(n24929), .IN2(n24928), .IN3(n24927), .IN4(n24926), 
        .QN(s11_addr_o[2]) );
  OA22X1 U28504 ( .IN1(n28601), .IN2(n25053), .IN3(n28603), .IN4(n25056), .Q(
        n24933) );
  OA22X1 U28505 ( .IN1(n28608), .IN2(n25051), .IN3(n28607), .IN4(n25028), .Q(
        n24932) );
  OA22X1 U28506 ( .IN1(n28604), .IN2(n25057), .IN3(n28606), .IN4(n25050), .Q(
        n24931) );
  OA22X1 U28507 ( .IN1(n28602), .IN2(n25039), .IN3(n28605), .IN4(n25055), .Q(
        n24930) );
  NAND4X0 U28508 ( .IN1(n24933), .IN2(n24932), .IN3(n24931), .IN4(n24930), 
        .QN(s11_addr_o[3]) );
  OA22X1 U28509 ( .IN1(n28614), .IN2(n25054), .IN3(n28617), .IN4(n25038), .Q(
        n24937) );
  OA22X1 U28510 ( .IN1(n28618), .IN2(n25028), .IN3(n28616), .IN4(n25044), .Q(
        n24936) );
  OA22X1 U28511 ( .IN1(n28619), .IN2(n25051), .IN3(n28615), .IN4(n25029), .Q(
        n24935) );
  OA22X1 U28512 ( .IN1(n28620), .IN2(n25045), .IN3(n28613), .IN4(n25011), .Q(
        n24934) );
  NAND4X0 U28513 ( .IN1(n24937), .IN2(n24936), .IN3(n24935), .IN4(n24934), 
        .QN(s11_addr_o[4]) );
  OA22X1 U28514 ( .IN1(n28630), .IN2(n25044), .IN3(n28629), .IN4(n25038), .Q(
        n24941) );
  OA22X1 U28515 ( .IN1(n28628), .IN2(n25056), .IN3(n28627), .IN4(n25039), .Q(
        n24940) );
  OA22X1 U28516 ( .IN1(n28632), .IN2(n25057), .IN3(n28631), .IN4(n25050), .Q(
        n24939) );
  OA22X1 U28517 ( .IN1(n28626), .IN2(n25028), .IN3(n28625), .IN4(n25051), .Q(
        n24938) );
  NAND4X0 U28518 ( .IN1(n24941), .IN2(n24940), .IN3(n24939), .IN4(n24938), 
        .QN(s11_addr_o[5]) );
  OA22X1 U28519 ( .IN1(n25028), .IN2(n28643), .IN3(n25006), .IN4(n28639), .Q(
        n24945) );
  OA22X1 U28520 ( .IN1(n25044), .IN2(n28640), .IN3(n25056), .IN4(n28641), .Q(
        n24944) );
  OA22X1 U28521 ( .IN1(n25011), .IN2(n28644), .IN3(n25029), .IN4(n28638), .Q(
        n24943) );
  OA22X1 U28522 ( .IN1(n25038), .IN2(n28642), .IN3(n25039), .IN4(n28637), .Q(
        n24942) );
  NAND4X0 U28523 ( .IN1(n24945), .IN2(n24944), .IN3(n24943), .IN4(n24942), 
        .QN(s11_addr_o[6]) );
  OA22X1 U28524 ( .IN1(n25055), .IN2(n28652), .IN3(n25011), .IN4(n28656), .Q(
        n24949) );
  OA22X1 U28525 ( .IN1(n25028), .IN2(n28653), .IN3(n25050), .IN4(n28650), .Q(
        n24948) );
  OA22X1 U28526 ( .IN1(n25045), .IN2(n28651), .IN3(n25006), .IN4(n28655), .Q(
        n24947) );
  OA22X1 U28527 ( .IN1(n25038), .IN2(n28654), .IN3(n25039), .IN4(n28649), .Q(
        n24946) );
  NAND4X0 U28528 ( .IN1(n24949), .IN2(n24948), .IN3(n24947), .IN4(n24946), 
        .QN(s11_addr_o[7]) );
  OA22X1 U28529 ( .IN1(n25029), .IN2(n28668), .IN3(n25054), .IN4(n28662), .Q(
        n24953) );
  OA22X1 U28530 ( .IN1(n25053), .IN2(n28664), .IN3(n25006), .IN4(n28667), .Q(
        n24952) );
  OA22X1 U28531 ( .IN1(n25055), .IN2(n28663), .IN3(n25056), .IN4(n28661), .Q(
        n24951) );
  OA22X1 U28532 ( .IN1(n25057), .IN2(n28666), .IN3(n25052), .IN4(n28665), .Q(
        n24950) );
  NAND4X0 U28533 ( .IN1(n24953), .IN2(n24952), .IN3(n24951), .IN4(n24950), 
        .QN(s11_addr_o[8]) );
  OA22X1 U28534 ( .IN1(n25054), .IN2(n28678), .IN3(n25006), .IN4(n28677), .Q(
        n24957) );
  OA22X1 U28535 ( .IN1(n25028), .IN2(n28676), .IN3(n25050), .IN4(n28673), .Q(
        n24956) );
  OA22X1 U28536 ( .IN1(n25055), .IN2(n28679), .IN3(n25056), .IN4(n28675), .Q(
        n24955) );
  OA22X1 U28537 ( .IN1(n25038), .IN2(n28680), .IN3(n25011), .IN4(n28674), .Q(
        n24954) );
  NAND4X0 U28538 ( .IN1(n24957), .IN2(n24956), .IN3(n24955), .IN4(n24954), 
        .QN(s11_addr_o[9]) );
  OA22X1 U28539 ( .IN1(n25028), .IN2(n28687), .IN3(n25006), .IN4(n28689), .Q(
        n24961) );
  OA22X1 U28540 ( .IN1(n25011), .IN2(n28688), .IN3(n25029), .IN4(n28685), .Q(
        n24960) );
  OA22X1 U28541 ( .IN1(n25038), .IN2(n28692), .IN3(n25044), .IN4(n28686), .Q(
        n24959) );
  OA22X1 U28542 ( .IN1(n25039), .IN2(n28691), .IN3(n25045), .IN4(n28690), .Q(
        n24958) );
  NAND4X0 U28543 ( .IN1(n24961), .IN2(n24960), .IN3(n24959), .IN4(n24958), 
        .QN(s11_addr_o[10]) );
  OA22X1 U28544 ( .IN1(n25057), .IN2(n28697), .IN3(n25039), .IN4(n28703), .Q(
        n24965) );
  OA22X1 U28545 ( .IN1(n25053), .IN2(n28702), .IN3(n25044), .IN4(n28698), .Q(
        n24964) );
  OA22X1 U28546 ( .IN1(n25056), .IN2(n28700), .IN3(n25006), .IN4(n28699), .Q(
        n24963) );
  OA22X1 U28547 ( .IN1(n25028), .IN2(n28704), .IN3(n25050), .IN4(n28701), .Q(
        n24962) );
  NAND4X0 U28548 ( .IN1(n24965), .IN2(n24964), .IN3(n24963), .IN4(n24962), 
        .QN(s11_addr_o[11]) );
  OA22X1 U28549 ( .IN1(n25044), .IN2(n28710), .IN3(n25006), .IN4(n28713), .Q(
        n24969) );
  OA22X1 U28550 ( .IN1(n25053), .IN2(n28714), .IN3(n25056), .IN4(n28711), .Q(
        n24968) );
  OA22X1 U28551 ( .IN1(n25011), .IN2(n28712), .IN3(n25029), .IN4(n28709), .Q(
        n24967) );
  OA22X1 U28552 ( .IN1(n25028), .IN2(n28716), .IN3(n25039), .IN4(n28715), .Q(
        n24966) );
  NAND4X0 U28553 ( .IN1(n24969), .IN2(n24968), .IN3(n24967), .IN4(n24966), 
        .QN(s11_addr_o[12]) );
  OA22X1 U28554 ( .IN1(n25053), .IN2(n28722), .IN3(n25050), .IN4(n28723), .Q(
        n24973) );
  OA22X1 U28555 ( .IN1(n25054), .IN2(n28721), .IN3(n25045), .IN4(n28725), .Q(
        n24972) );
  OA22X1 U28556 ( .IN1(n25057), .IN2(n28726), .IN3(n25052), .IN4(n28724), .Q(
        n24971) );
  OA22X1 U28557 ( .IN1(n25055), .IN2(n28728), .IN3(n25006), .IN4(n28727), .Q(
        n24970) );
  NAND4X0 U28558 ( .IN1(n24973), .IN2(n24972), .IN3(n24971), .IN4(n24970), 
        .QN(s11_addr_o[13]) );
  OA22X1 U28559 ( .IN1(n25038), .IN2(n28734), .IN3(n25029), .IN4(n28740), .Q(
        n24977) );
  OA22X1 U28560 ( .IN1(n25044), .IN2(n28738), .IN3(n25045), .IN4(n28733), .Q(
        n24976) );
  OA22X1 U28561 ( .IN1(n25011), .IN2(n28736), .IN3(n25052), .IN4(n28735), .Q(
        n24975) );
  OA22X1 U28562 ( .IN1(n25039), .IN2(n28737), .IN3(n25006), .IN4(n28739), .Q(
        n24974) );
  NAND4X0 U28563 ( .IN1(n24977), .IN2(n24976), .IN3(n24975), .IN4(n24974), 
        .QN(s11_addr_o[14]) );
  OA22X1 U28564 ( .IN1(n25029), .IN2(n28747), .IN3(n25056), .IN4(n28749), .Q(
        n24981) );
  OA22X1 U28565 ( .IN1(n25054), .IN2(n28751), .IN3(n25006), .IN4(n28745), .Q(
        n24980) );
  OA22X1 U28566 ( .IN1(n25053), .IN2(n28746), .IN3(n25044), .IN4(n28748), .Q(
        n24979) );
  OA22X1 U28567 ( .IN1(n25011), .IN2(n28750), .IN3(n25052), .IN4(n28752), .Q(
        n24978) );
  NAND4X0 U28568 ( .IN1(n24981), .IN2(n24980), .IN3(n24979), .IN4(n24978), 
        .QN(s11_addr_o[15]) );
  OA22X1 U28569 ( .IN1(n25054), .IN2(n28757), .IN3(n25006), .IN4(n28763), .Q(
        n24985) );
  OA22X1 U28570 ( .IN1(n25028), .IN2(n28761), .IN3(n25045), .IN4(n28764), .Q(
        n24984) );
  OA22X1 U28571 ( .IN1(n25044), .IN2(n28762), .IN3(n25011), .IN4(n28760), .Q(
        n24983) );
  OA22X1 U28572 ( .IN1(n25053), .IN2(n28758), .IN3(n25050), .IN4(n28759), .Q(
        n24982) );
  NAND4X0 U28573 ( .IN1(n24985), .IN2(n24984), .IN3(n24983), .IN4(n24982), 
        .QN(s11_addr_o[16]) );
  OA22X1 U28574 ( .IN1(n25028), .IN2(n28773), .IN3(n25045), .IN4(n28770), .Q(
        n24989) );
  OA22X1 U28575 ( .IN1(n25038), .IN2(n28772), .IN3(n25039), .IN4(n28771), .Q(
        n24988) );
  OA22X1 U28576 ( .IN1(n25029), .IN2(n28775), .IN3(n25006), .IN4(n28769), .Q(
        n24987) );
  OA22X1 U28577 ( .IN1(n25044), .IN2(n28776), .IN3(n25011), .IN4(n28774), .Q(
        n24986) );
  NAND4X0 U28578 ( .IN1(n24989), .IN2(n24988), .IN3(n24987), .IN4(n24986), 
        .QN(s11_addr_o[17]) );
  OA22X1 U28579 ( .IN1(n25053), .IN2(n28786), .IN3(n25054), .IN4(n28783), .Q(
        n24993) );
  OA22X1 U28580 ( .IN1(n25029), .IN2(n28784), .IN3(n25006), .IN4(n28781), .Q(
        n24992) );
  OA22X1 U28581 ( .IN1(n25055), .IN2(n28788), .IN3(n25045), .IN4(n28785), .Q(
        n24991) );
  OA22X1 U28582 ( .IN1(n25057), .IN2(n28787), .IN3(n25052), .IN4(n28782), .Q(
        n24990) );
  NAND4X0 U28583 ( .IN1(n24993), .IN2(n24992), .IN3(n24991), .IN4(n24990), 
        .QN(s11_addr_o[18]) );
  OA22X1 U28584 ( .IN1(n25057), .IN2(n28798), .IN3(n25050), .IN4(n28797), .Q(
        n24997) );
  OA22X1 U28585 ( .IN1(n25055), .IN2(n28800), .IN3(n25039), .IN4(n28795), .Q(
        n24996) );
  OA22X1 U28586 ( .IN1(n25052), .IN2(n28794), .IN3(n25006), .IN4(n28799), .Q(
        n24995) );
  OA22X1 U28587 ( .IN1(n25038), .IN2(n28796), .IN3(n25056), .IN4(n28793), .Q(
        n24994) );
  NAND4X0 U28588 ( .IN1(n24997), .IN2(n24996), .IN3(n24995), .IN4(n24994), 
        .QN(s11_addr_o[19]) );
  OA22X1 U28589 ( .IN1(n25028), .IN2(n28810), .IN3(n25050), .IN4(n28806), .Q(
        n25001) );
  OA22X1 U28590 ( .IN1(n25044), .IN2(n28808), .IN3(n25056), .IN4(n28809), .Q(
        n25000) );
  OA22X1 U28591 ( .IN1(n25057), .IN2(n28807), .IN3(n25006), .IN4(n28805), .Q(
        n24999) );
  OA22X1 U28592 ( .IN1(n25053), .IN2(n28812), .IN3(n25054), .IN4(n28811), .Q(
        n24998) );
  NAND4X0 U28593 ( .IN1(n25001), .IN2(n25000), .IN3(n24999), .IN4(n24998), 
        .QN(s11_addr_o[20]) );
  OA22X1 U28594 ( .IN1(n25055), .IN2(n28824), .IN3(n25054), .IN4(n28823), .Q(
        n25005) );
  OA22X1 U28595 ( .IN1(n25028), .IN2(n28819), .IN3(n25050), .IN4(n28821), .Q(
        n25004) );
  OA22X1 U28596 ( .IN1(n25045), .IN2(n28818), .IN3(n25006), .IN4(n28817), .Q(
        n25003) );
  OA22X1 U28597 ( .IN1(n25053), .IN2(n28822), .IN3(n25011), .IN4(n28820), .Q(
        n25002) );
  NAND4X0 U28598 ( .IN1(n25005), .IN2(n25004), .IN3(n25003), .IN4(n25002), 
        .QN(s11_addr_o[21]) );
  OA22X1 U28599 ( .IN1(n25029), .IN2(n28836), .IN3(n25006), .IN4(n28829), .Q(
        n25010) );
  OA22X1 U28600 ( .IN1(n25038), .IN2(n28833), .IN3(n25045), .IN4(n28837), .Q(
        n25009) );
  OA22X1 U28601 ( .IN1(n25057), .IN2(n28831), .IN3(n25039), .IN4(n28834), .Q(
        n25008) );
  OA22X1 U28602 ( .IN1(n25044), .IN2(n28832), .IN3(n25052), .IN4(n28838), .Q(
        n25007) );
  NAND4X0 U28603 ( .IN1(n25010), .IN2(n25009), .IN3(n25008), .IN4(n25007), 
        .QN(s11_addr_o[22]) );
  OA22X1 U28604 ( .IN1(n25038), .IN2(n28848), .IN3(n25011), .IN4(n28843), .Q(
        n25015) );
  OA22X1 U28605 ( .IN1(n25029), .IN2(n28852), .IN3(n25054), .IN4(n28849), .Q(
        n25014) );
  OA22X1 U28606 ( .IN1(n25028), .IN2(n28850), .IN3(n25051), .IN4(n28851), .Q(
        n25013) );
  OA22X1 U28607 ( .IN1(n25055), .IN2(n28845), .IN3(n25056), .IN4(n28846), .Q(
        n25012) );
  NAND4X0 U28608 ( .IN1(n25015), .IN2(n25014), .IN3(n25013), .IN4(n25012), 
        .QN(s11_addr_o[23]) );
  OA22X1 U28609 ( .IN1(n28864), .IN2(n25055), .IN3(n28857), .IN4(n25052), .Q(
        n25019) );
  OA22X1 U28610 ( .IN1(n28859), .IN2(n25039), .IN3(n28863), .IN4(n25038), .Q(
        n25018) );
  OA22X1 U28611 ( .IN1(n28860), .IN2(n25051), .IN3(n28861), .IN4(n25029), .Q(
        n25017) );
  OA22X1 U28612 ( .IN1(n28858), .IN2(n25057), .IN3(n28865), .IN4(n25056), .Q(
        n25016) );
  NAND4X0 U28613 ( .IN1(n25019), .IN2(n25018), .IN3(n25017), .IN4(n25016), 
        .QN(s11_addr_o[24]) );
  OA22X1 U28614 ( .IN1(n28877), .IN2(n25055), .IN3(n28875), .IN4(n25051), .Q(
        n25023) );
  OA22X1 U28615 ( .IN1(n28871), .IN2(n25045), .IN3(n28874), .IN4(n25052), .Q(
        n25022) );
  OA22X1 U28616 ( .IN1(n28873), .IN2(n25057), .IN3(n28876), .IN4(n25054), .Q(
        n25021) );
  OA22X1 U28617 ( .IN1(n28870), .IN2(n25038), .IN3(n28872), .IN4(n25050), .Q(
        n25020) );
  NAND4X0 U28618 ( .IN1(n25023), .IN2(n25022), .IN3(n25021), .IN4(n25020), 
        .QN(s11_addr_o[25]) );
  OA22X1 U28619 ( .IN1(n28885), .IN2(n25057), .IN3(n28882), .IN4(n25052), .Q(
        n25027) );
  OA22X1 U28620 ( .IN1(n28883), .IN2(n25056), .IN3(n28887), .IN4(n25044), .Q(
        n25026) );
  OA22X1 U28621 ( .IN1(n28888), .IN2(n25054), .IN3(n28886), .IN4(n25050), .Q(
        n25025) );
  OA22X1 U28622 ( .IN1(n28889), .IN2(n25051), .IN3(n28884), .IN4(n25038), .Q(
        n25024) );
  NAND4X0 U28623 ( .IN1(n25027), .IN2(n25026), .IN3(n25025), .IN4(n25024), 
        .QN(s11_addr_o[26]) );
  OA22X1 U28624 ( .IN1(n28896), .IN2(n25039), .IN3(n28901), .IN4(n25028), .Q(
        n25033) );
  OA22X1 U28625 ( .IN1(n28895), .IN2(n25044), .IN3(n28900), .IN4(n25029), .Q(
        n25032) );
  OA22X1 U28626 ( .IN1(n28899), .IN2(n25057), .IN3(n28894), .IN4(n25038), .Q(
        n25031) );
  OA22X1 U28627 ( .IN1(n28897), .IN2(n25045), .IN3(n28898), .IN4(n25051), .Q(
        n25030) );
  NAND4X0 U28628 ( .IN1(n25033), .IN2(n25032), .IN3(n25031), .IN4(n25030), 
        .QN(s11_addr_o[27]) );
  OA22X1 U28629 ( .IN1(n28911), .IN2(n25055), .IN3(n28908), .IN4(n25052), .Q(
        n25037) );
  OA22X1 U28630 ( .IN1(n28907), .IN2(n25056), .IN3(n28906), .IN4(n25050), .Q(
        n25036) );
  OA22X1 U28631 ( .IN1(n28910), .IN2(n25054), .IN3(n28912), .IN4(n25038), .Q(
        n25035) );
  OA22X1 U28632 ( .IN1(n28909), .IN2(n25057), .IN3(n28913), .IN4(n25051), .Q(
        n25034) );
  NAND4X0 U28633 ( .IN1(n25037), .IN2(n25036), .IN3(n25035), .IN4(n25034), 
        .QN(s11_addr_o[28]) );
  OA22X1 U28634 ( .IN1(n28925), .IN2(n25038), .IN3(n28923), .IN4(n25050), .Q(
        n25043) );
  OA22X1 U28635 ( .IN1(n28920), .IN2(n25039), .IN3(n28919), .IN4(n25052), .Q(
        n25042) );
  OA22X1 U28636 ( .IN1(n28926), .IN2(n25057), .IN3(n28922), .IN4(n25045), .Q(
        n25041) );
  OA22X1 U28637 ( .IN1(n28924), .IN2(n25044), .IN3(n28921), .IN4(n25051), .Q(
        n25040) );
  NAND4X0 U28638 ( .IN1(n25043), .IN2(n25042), .IN3(n25041), .IN4(n25040), 
        .QN(s11_addr_o[29]) );
  OA22X1 U28639 ( .IN1(n28932), .IN2(n25057), .IN3(n28933), .IN4(n25051), .Q(
        n25049) );
  OA22X1 U28640 ( .IN1(n28935), .IN2(n25044), .IN3(n28940), .IN4(n25052), .Q(
        n25048) );
  OA22X1 U28641 ( .IN1(n28931), .IN2(n25053), .IN3(n28939), .IN4(n25050), .Q(
        n25047) );
  OA22X1 U28642 ( .IN1(n28937), .IN2(n25045), .IN3(n28936), .IN4(n25054), .Q(
        n25046) );
  NAND4X0 U28643 ( .IN1(n25049), .IN2(n25048), .IN3(n25047), .IN4(n25046), 
        .QN(s11_addr_o[30]) );
  OA22X1 U28644 ( .IN1(n28960), .IN2(n25051), .IN3(n28946), .IN4(n25050), .Q(
        n25061) );
  OA22X1 U28645 ( .IN1(n28950), .IN2(n25053), .IN3(n28958), .IN4(n25052), .Q(
        n25060) );
  OA22X1 U28646 ( .IN1(n28952), .IN2(n25055), .IN3(n28954), .IN4(n25054), .Q(
        n25059) );
  OA22X1 U28647 ( .IN1(n28948), .IN2(n25057), .IN3(n28956), .IN4(n25056), .Q(
        n25058) );
  NAND4X0 U28648 ( .IN1(n25061), .IN2(n25060), .IN3(n25059), .IN4(n25058), 
        .QN(s11_addr_o[31]) );
  OA22X1 U28649 ( .IN1(n29273), .IN2(n25063), .IN3(n29254), .IN4(n25062), .Q(
        n25074) );
  INVX0 U28650 ( .INP(n25064), .ZN(n25066) );
  OA22X1 U28651 ( .IN1(n29235), .IN2(n25066), .IN3(n29292), .IN4(n25065), .Q(
        n25073) );
  OA22X1 U28652 ( .IN1(n29349), .IN2(n25068), .IN3(n29311), .IN4(n25067), .Q(
        n25072) );
  OA22X1 U28653 ( .IN1(n29368), .IN2(n25070), .IN3(n29330), .IN4(n25069), .Q(
        n25071) );
  NAND4X0 U28654 ( .IN1(n25074), .IN2(n25073), .IN3(n25072), .IN4(n25071), 
        .QN(s10_stb_o) );
  INVX0 U28655 ( .INP(n29155), .ZN(n25359) );
  INVX0 U28656 ( .INP(n29146), .ZN(n25347) );
  OA22X1 U28657 ( .IN1(n25359), .IN2(n28124), .IN3(n25347), .IN4(n28121), .Q(
        n25078) );
  INVX0 U28658 ( .INP(n29148), .ZN(n25350) );
  INVX0 U28659 ( .INP(n29154), .ZN(n25357) );
  OA22X1 U28660 ( .IN1(n25350), .IN2(n28123), .IN3(n25357), .IN4(n28122), .Q(
        n25077) );
  INVX0 U28661 ( .INP(n29147), .ZN(n25361) );
  INVX0 U28662 ( .INP(n29156), .ZN(n25345) );
  OA22X1 U28663 ( .IN1(n25361), .IN2(n28126), .IN3(n25345), .IN4(n28125), .Q(
        n25076) );
  INVX0 U28664 ( .INP(n29153), .ZN(n25360) );
  OA22X1 U28665 ( .IN1(n25360), .IN2(n28128), .IN3(n25355), .IN4(n28127), .Q(
        n25075) );
  NAND4X0 U28666 ( .IN1(n25078), .IN2(n25077), .IN3(n25076), .IN4(n25075), 
        .QN(s10_we_o) );
  OA22X1 U28667 ( .IN1(n25350), .IN2(n28133), .IN3(n25347), .IN4(n28135), .Q(
        n25082) );
  INVX0 U28668 ( .INP(n29154), .ZN(n25307) );
  OA22X1 U28669 ( .IN1(n25360), .IN2(n28140), .IN3(n25307), .IN4(n28138), .Q(
        n25081) );
  OA22X1 U28670 ( .IN1(n25359), .IN2(n28134), .IN3(n25355), .IN4(n28137), .Q(
        n25080) );
  INVX0 U28671 ( .INP(n29147), .ZN(n25340) );
  OA22X1 U28672 ( .IN1(n25340), .IN2(n28139), .IN3(n25345), .IN4(n28136), .Q(
        n25079) );
  NAND4X0 U28673 ( .IN1(n25082), .IN2(n25081), .IN3(n25080), .IN4(n25079), 
        .QN(s10_data_o[0]) );
  OA22X1 U28674 ( .IN1(n25359), .IN2(n28150), .IN3(n25345), .IN4(n28152), .Q(
        n25086) );
  INVX0 U28675 ( .INP(n29153), .ZN(n25349) );
  OA22X1 U28676 ( .IN1(n25349), .IN2(n28146), .IN3(n25350), .IN4(n28148), .Q(
        n25085) );
  INVX0 U28677 ( .INP(n25355), .ZN(n29145) );
  INVX0 U28678 ( .INP(n29145), .ZN(n25346) );
  OA22X1 U28679 ( .IN1(n25346), .IN2(n28151), .IN3(n25347), .IN4(n28147), .Q(
        n25084) );
  OA22X1 U28680 ( .IN1(n25340), .IN2(n28145), .IN3(n25307), .IN4(n28149), .Q(
        n25083) );
  NAND4X0 U28681 ( .IN1(n25086), .IN2(n25085), .IN3(n25084), .IN4(n25083), 
        .QN(s10_data_o[1]) );
  OA22X1 U28682 ( .IN1(n25349), .IN2(n28164), .IN3(n25355), .IN4(n28157), .Q(
        n25090) );
  OA22X1 U28683 ( .IN1(n25361), .IN2(n28159), .IN3(n25347), .IN4(n28161), .Q(
        n25089) );
  INVX0 U28684 ( .INP(n29148), .ZN(n25356) );
  OA22X1 U28685 ( .IN1(n25356), .IN2(n28163), .IN3(n25307), .IN4(n28158), .Q(
        n25088) );
  OA22X1 U28686 ( .IN1(n25359), .IN2(n28160), .IN3(n25345), .IN4(n28162), .Q(
        n25087) );
  NAND4X0 U28687 ( .IN1(n25090), .IN2(n25089), .IN3(n25088), .IN4(n25087), 
        .QN(s10_data_o[2]) );
  OA22X1 U28688 ( .IN1(n25348), .IN2(n28172), .IN3(n25350), .IN4(n28176), .Q(
        n25094) );
  OA22X1 U28689 ( .IN1(n25346), .IN2(n28169), .IN3(n25347), .IN4(n28173), .Q(
        n25093) );
  OA22X1 U28690 ( .IN1(n25349), .IN2(n28174), .IN3(n25340), .IN4(n28170), .Q(
        n25092) );
  OA22X1 U28691 ( .IN1(n25307), .IN2(n28171), .IN3(n25345), .IN4(n28175), .Q(
        n25091) );
  NAND4X0 U28692 ( .IN1(n25094), .IN2(n25093), .IN3(n25092), .IN4(n25091), 
        .QN(s10_data_o[3]) );
  OA22X1 U28693 ( .IN1(n25359), .IN2(n28182), .IN3(n25360), .IN4(n28184), .Q(
        n25098) );
  OA22X1 U28694 ( .IN1(n25357), .IN2(n28185), .IN3(n25355), .IN4(n28187), .Q(
        n25097) );
  OA22X1 U28695 ( .IN1(n25350), .IN2(n28186), .IN3(n25345), .IN4(n28183), .Q(
        n25096) );
  OA22X1 U28696 ( .IN1(n25340), .IN2(n28188), .IN3(n25347), .IN4(n28181), .Q(
        n25095) );
  NAND4X0 U28697 ( .IN1(n25098), .IN2(n25097), .IN3(n25096), .IN4(n25095), 
        .QN(s10_data_o[4]) );
  OA22X1 U28698 ( .IN1(n25349), .IN2(n28200), .IN3(n25340), .IN4(n28193), .Q(
        n25102) );
  OA22X1 U28699 ( .IN1(n25350), .IN2(n28194), .IN3(n25307), .IN4(n28198), .Q(
        n25101) );
  OA22X1 U28700 ( .IN1(n25346), .IN2(n28195), .IN3(n25347), .IN4(n28199), .Q(
        n25100) );
  INVX0 U28701 ( .INP(n29156), .ZN(n25358) );
  OA22X1 U28702 ( .IN1(n25348), .IN2(n28196), .IN3(n25358), .IN4(n28197), .Q(
        n25099) );
  NAND4X0 U28703 ( .IN1(n25102), .IN2(n25101), .IN3(n25100), .IN4(n25099), 
        .QN(s10_data_o[5]) );
  OA22X1 U28704 ( .IN1(n25349), .IN2(n28207), .IN3(n25307), .IN4(n28211), .Q(
        n25106) );
  OA22X1 U28705 ( .IN1(n25359), .IN2(n28208), .IN3(n25347), .IN4(n28209), .Q(
        n25105) );
  OA22X1 U28706 ( .IN1(n25340), .IN2(n28212), .IN3(n25345), .IN4(n28205), .Q(
        n25104) );
  OA22X1 U28707 ( .IN1(n25356), .IN2(n28206), .IN3(n25355), .IN4(n28210), .Q(
        n25103) );
  NAND4X0 U28708 ( .IN1(n25106), .IN2(n25105), .IN3(n25104), .IN4(n25103), 
        .QN(s10_data_o[6]) );
  OA22X1 U28709 ( .IN1(n25361), .IN2(n28218), .IN3(n25355), .IN4(n28222), .Q(
        n25110) );
  OA22X1 U28710 ( .IN1(n25348), .IN2(n28220), .IN3(n25360), .IN4(n28219), .Q(
        n25109) );
  OA22X1 U28711 ( .IN1(n25345), .IN2(n28223), .IN3(n25347), .IN4(n28221), .Q(
        n25108) );
  OA22X1 U28712 ( .IN1(n25350), .IN2(n28224), .IN3(n25307), .IN4(n28217), .Q(
        n25107) );
  NAND4X0 U28713 ( .IN1(n25110), .IN2(n25109), .IN3(n25108), .IN4(n25107), 
        .QN(s10_data_o[7]) );
  OA22X1 U28714 ( .IN1(n25349), .IN2(n28232), .IN3(n25307), .IN4(n28236), .Q(
        n25114) );
  OA22X1 U28715 ( .IN1(n25359), .IN2(n28230), .IN3(n25350), .IN4(n28231), .Q(
        n25113) );
  OA22X1 U28716 ( .IN1(n25361), .IN2(n28234), .IN3(n25358), .IN4(n28229), .Q(
        n25112) );
  INVX0 U28717 ( .INP(n29146), .ZN(n25362) );
  OA22X1 U28718 ( .IN1(n25346), .IN2(n28233), .IN3(n25362), .IN4(n28235), .Q(
        n25111) );
  NAND4X0 U28719 ( .IN1(n25114), .IN2(n25113), .IN3(n25112), .IN4(n25111), 
        .QN(s10_data_o[8]) );
  OA22X1 U28720 ( .IN1(n25340), .IN2(n28248), .IN3(n25307), .IN4(n28241), .Q(
        n25118) );
  OA22X1 U28721 ( .IN1(n25349), .IN2(n28244), .IN3(n25355), .IN4(n28243), .Q(
        n25117) );
  OA22X1 U28722 ( .IN1(n25358), .IN2(n28245), .IN3(n25362), .IN4(n28247), .Q(
        n25116) );
  OA22X1 U28723 ( .IN1(n25348), .IN2(n28242), .IN3(n25350), .IN4(n28246), .Q(
        n25115) );
  NAND4X0 U28724 ( .IN1(n25118), .IN2(n25117), .IN3(n25116), .IN4(n25115), 
        .QN(s10_data_o[9]) );
  OA22X1 U28725 ( .IN1(n25356), .IN2(n28260), .IN3(n25340), .IN4(n28256), .Q(
        n25122) );
  OA22X1 U28726 ( .IN1(n25359), .IN2(n28258), .IN3(n25362), .IN4(n28259), .Q(
        n25121) );
  OA22X1 U28727 ( .IN1(n25349), .IN2(n28257), .IN3(n25345), .IN4(n28255), .Q(
        n25120) );
  OA22X1 U28728 ( .IN1(n25307), .IN2(n28254), .IN3(n25355), .IN4(n28253), .Q(
        n25119) );
  NAND4X0 U28729 ( .IN1(n25122), .IN2(n25121), .IN3(n25120), .IN4(n25119), 
        .QN(s10_data_o[10]) );
  OA22X1 U28730 ( .IN1(n25350), .IN2(n28265), .IN3(n25340), .IN4(n28271), .Q(
        n25126) );
  OA22X1 U28731 ( .IN1(n25349), .IN2(n28272), .IN3(n25358), .IN4(n28270), .Q(
        n25125) );
  OA22X1 U28732 ( .IN1(n25357), .IN2(n28268), .IN3(n25362), .IN4(n28269), .Q(
        n25124) );
  OA22X1 U28733 ( .IN1(n25348), .IN2(n28266), .IN3(n25355), .IN4(n28267), .Q(
        n25123) );
  NAND4X0 U28734 ( .IN1(n25126), .IN2(n25125), .IN3(n25124), .IN4(n25123), 
        .QN(s10_data_o[11]) );
  OA22X1 U28735 ( .IN1(n25340), .IN2(n28282), .IN3(n25362), .IN4(n28277), .Q(
        n25130) );
  OA22X1 U28736 ( .IN1(n25350), .IN2(n28280), .IN3(n25345), .IN4(n28281), .Q(
        n25129) );
  OA22X1 U28737 ( .IN1(n25307), .IN2(n28283), .IN3(n25355), .IN4(n28279), .Q(
        n25128) );
  OA22X1 U28738 ( .IN1(n25359), .IN2(n28284), .IN3(n25360), .IN4(n28278), .Q(
        n25127) );
  NAND4X0 U28739 ( .IN1(n25130), .IN2(n25129), .IN3(n25128), .IN4(n25127), 
        .QN(s10_data_o[12]) );
  OA22X1 U28740 ( .IN1(n25348), .IN2(n28290), .IN3(n25307), .IN4(n28289), .Q(
        n25134) );
  OA22X1 U28741 ( .IN1(n25349), .IN2(n28294), .IN3(n25362), .IN4(n28295), .Q(
        n25133) );
  OA22X1 U28742 ( .IN1(n25345), .IN2(n28293), .IN3(n25355), .IN4(n28291), .Q(
        n25132) );
  OA22X1 U28743 ( .IN1(n25356), .IN2(n28296), .IN3(n25340), .IN4(n28292), .Q(
        n25131) );
  NAND4X0 U28744 ( .IN1(n25134), .IN2(n25133), .IN3(n25132), .IN4(n25131), 
        .QN(s10_data_o[13]) );
  OA22X1 U28745 ( .IN1(n25359), .IN2(n28306), .IN3(n25350), .IN4(n28308), .Q(
        n25138) );
  OA22X1 U28746 ( .IN1(n25355), .IN2(n28301), .IN3(n25362), .IN4(n28303), .Q(
        n25137) );
  OA22X1 U28747 ( .IN1(n25349), .IN2(n28304), .IN3(n25345), .IN4(n28302), .Q(
        n25136) );
  OA22X1 U28748 ( .IN1(n25361), .IN2(n28305), .IN3(n25307), .IN4(n28307), .Q(
        n25135) );
  NAND4X0 U28749 ( .IN1(n25138), .IN2(n25137), .IN3(n25136), .IN4(n25135), 
        .QN(s10_data_o[14]) );
  OA22X1 U28750 ( .IN1(n25358), .IN2(n28318), .IN3(n25362), .IN4(n28319), .Q(
        n25142) );
  OA22X1 U28751 ( .IN1(n25360), .IN2(n28315), .IN3(n25361), .IN4(n28313), .Q(
        n25141) );
  OA22X1 U28752 ( .IN1(n25348), .IN2(n28316), .IN3(n25346), .IN4(n28317), .Q(
        n25140) );
  OA22X1 U28753 ( .IN1(n25350), .IN2(n28314), .IN3(n25307), .IN4(n28320), .Q(
        n25139) );
  NAND4X0 U28754 ( .IN1(n25142), .IN2(n25141), .IN3(n25140), .IN4(n25139), 
        .QN(s10_data_o[15]) );
  OA22X1 U28755 ( .IN1(n25350), .IN2(n28331), .IN3(n25307), .IN4(n28329), .Q(
        n25146) );
  OA22X1 U28756 ( .IN1(n25340), .IN2(n28326), .IN3(n25362), .IN4(n28327), .Q(
        n25145) );
  OA22X1 U28757 ( .IN1(n25345), .IN2(n28325), .IN3(n25346), .IN4(n28328), .Q(
        n25144) );
  OA22X1 U28758 ( .IN1(n25359), .IN2(n28330), .IN3(n25360), .IN4(n28332), .Q(
        n25143) );
  NAND4X0 U28759 ( .IN1(n25146), .IN2(n25145), .IN3(n25144), .IN4(n25143), 
        .QN(s10_data_o[16]) );
  OA22X1 U28760 ( .IN1(n25360), .IN2(n28344), .IN3(n25362), .IN4(n28341), .Q(
        n25150) );
  OA22X1 U28761 ( .IN1(n25348), .IN2(n28340), .IN3(n25345), .IN4(n28339), .Q(
        n25149) );
  OA22X1 U28762 ( .IN1(n25350), .IN2(n28342), .IN3(n25307), .IN4(n28337), .Q(
        n25148) );
  OA22X1 U28763 ( .IN1(n25361), .IN2(n28338), .IN3(n25346), .IN4(n28343), .Q(
        n25147) );
  NAND4X0 U28764 ( .IN1(n25150), .IN2(n25149), .IN3(n25148), .IN4(n25147), 
        .QN(s10_data_o[17]) );
  OA22X1 U28765 ( .IN1(n25348), .IN2(n28352), .IN3(n25350), .IN4(n28350), .Q(
        n25154) );
  OA22X1 U28766 ( .IN1(n25361), .IN2(n28355), .IN3(n25358), .IN4(n28349), .Q(
        n25153) );
  OA22X1 U28767 ( .IN1(n25349), .IN2(n28356), .IN3(n25362), .IN4(n28353), .Q(
        n25152) );
  OA22X1 U28768 ( .IN1(n25357), .IN2(n28354), .IN3(n25346), .IN4(n28351), .Q(
        n25151) );
  NAND4X0 U28769 ( .IN1(n25154), .IN2(n25153), .IN3(n25152), .IN4(n25151), 
        .QN(s10_data_o[18]) );
  OA22X1 U28770 ( .IN1(n25340), .IN2(n28363), .IN3(n25358), .IN4(n28361), .Q(
        n25158) );
  OA22X1 U28771 ( .IN1(n25360), .IN2(n28364), .IN3(n25350), .IN4(n28362), .Q(
        n25157) );
  OA22X1 U28772 ( .IN1(n25307), .IN2(n28365), .IN3(n25346), .IN4(n28368), .Q(
        n25156) );
  OA22X1 U28773 ( .IN1(n25348), .IN2(n28366), .IN3(n25362), .IN4(n28367), .Q(
        n25155) );
  NAND4X0 U28774 ( .IN1(n25158), .IN2(n25157), .IN3(n25156), .IN4(n25155), 
        .QN(s10_data_o[19]) );
  OA22X1 U28775 ( .IN1(n25356), .IN2(n28374), .IN3(n25358), .IN4(n28380), .Q(
        n25162) );
  OA22X1 U28776 ( .IN1(n25349), .IN2(n28377), .IN3(n25362), .IN4(n28375), .Q(
        n25161) );
  OA22X1 U28777 ( .IN1(n25348), .IN2(n28378), .IN3(n25361), .IN4(n28373), .Q(
        n25160) );
  OA22X1 U28778 ( .IN1(n25357), .IN2(n28376), .IN3(n25346), .IN4(n28379), .Q(
        n25159) );
  NAND4X0 U28779 ( .IN1(n25162), .IN2(n25161), .IN3(n25160), .IN4(n25159), 
        .QN(s10_data_o[20]) );
  OA22X1 U28780 ( .IN1(n25348), .IN2(n28392), .IN3(n25360), .IN4(n28386), .Q(
        n25166) );
  OA22X1 U28781 ( .IN1(n25358), .IN2(n28385), .IN3(n25346), .IN4(n28389), .Q(
        n25165) );
  OA22X1 U28782 ( .IN1(n25350), .IN2(n28390), .IN3(n25307), .IN4(n28387), .Q(
        n25164) );
  OA22X1 U28783 ( .IN1(n25340), .IN2(n28388), .IN3(n25362), .IN4(n28391), .Q(
        n25163) );
  NAND4X0 U28784 ( .IN1(n25166), .IN2(n25165), .IN3(n25164), .IN4(n25163), 
        .QN(s10_data_o[21]) );
  OA22X1 U28785 ( .IN1(n25345), .IN2(n28399), .IN3(n25362), .IN4(n28397), .Q(
        n25170) );
  OA22X1 U28786 ( .IN1(n25348), .IN2(n28400), .IN3(n25361), .IN4(n28403), .Q(
        n25169) );
  OA22X1 U28787 ( .IN1(n25349), .IN2(n28402), .IN3(n25356), .IN4(n28404), .Q(
        n25168) );
  OA22X1 U28788 ( .IN1(n25357), .IN2(n28398), .IN3(n25346), .IN4(n28401), .Q(
        n25167) );
  NAND4X0 U28789 ( .IN1(n25170), .IN2(n25169), .IN3(n25168), .IN4(n25167), 
        .QN(s10_data_o[22]) );
  OA22X1 U28790 ( .IN1(n25348), .IN2(n28416), .IN3(n25350), .IN4(n28414), .Q(
        n25174) );
  OA22X1 U28791 ( .IN1(n25360), .IN2(n28415), .IN3(n25340), .IN4(n28413), .Q(
        n25173) );
  OA22X1 U28792 ( .IN1(n25358), .IN2(n28412), .IN3(n25346), .IN4(n28409), .Q(
        n25172) );
  OA22X1 U28793 ( .IN1(n25357), .IN2(n28410), .IN3(n25362), .IN4(n28411), .Q(
        n25171) );
  NAND4X0 U28794 ( .IN1(n25174), .IN2(n25173), .IN3(n25172), .IN4(n25171), 
        .QN(s10_data_o[23]) );
  OA22X1 U28795 ( .IN1(n25348), .IN2(n28426), .IN3(n25360), .IN4(n28424), .Q(
        n25178) );
  OA22X1 U28796 ( .IN1(n25345), .IN2(n28428), .IN3(n25362), .IN4(n28423), .Q(
        n25177) );
  OA22X1 U28797 ( .IN1(n25361), .IN2(n28421), .IN3(n25307), .IN4(n28425), .Q(
        n25176) );
  OA22X1 U28798 ( .IN1(n25356), .IN2(n28422), .IN3(n25346), .IN4(n28427), .Q(
        n25175) );
  NAND4X0 U28799 ( .IN1(n25178), .IN2(n25177), .IN3(n25176), .IN4(n25175), 
        .QN(s10_data_o[24]) );
  OA22X1 U28800 ( .IN1(n25361), .IN2(n28439), .IN3(n25307), .IN4(n28433), .Q(
        n25182) );
  OA22X1 U28801 ( .IN1(n25360), .IN2(n28440), .IN3(n25350), .IN4(n28434), .Q(
        n25181) );
  OA22X1 U28802 ( .IN1(n25348), .IN2(n28438), .IN3(n25346), .IN4(n28436), .Q(
        n25180) );
  OA22X1 U28803 ( .IN1(n25358), .IN2(n28437), .IN3(n25362), .IN4(n28435), .Q(
        n25179) );
  NAND4X0 U28804 ( .IN1(n25182), .IN2(n25181), .IN3(n25180), .IN4(n25179), 
        .QN(s10_data_o[25]) );
  OA22X1 U28805 ( .IN1(n25349), .IN2(n28451), .IN3(n25307), .IN4(n28449), .Q(
        n25186) );
  OA22X1 U28806 ( .IN1(n25356), .IN2(n28450), .IN3(n25346), .IN4(n28447), .Q(
        n25185) );
  OA22X1 U28807 ( .IN1(n25361), .IN2(n28446), .IN3(n25345), .IN4(n28448), .Q(
        n25184) );
  OA22X1 U28808 ( .IN1(n25348), .IN2(n28452), .IN3(n25347), .IN4(n28445), .Q(
        n25183) );
  NAND4X0 U28809 ( .IN1(n25186), .IN2(n25185), .IN3(n25184), .IN4(n25183), 
        .QN(s10_data_o[26]) );
  OA22X1 U28810 ( .IN1(n25345), .IN2(n28463), .IN3(n25346), .IN4(n28460), .Q(
        n25190) );
  OA22X1 U28811 ( .IN1(n25356), .IN2(n28464), .IN3(n25340), .IN4(n28458), .Q(
        n25189) );
  OA22X1 U28812 ( .IN1(n25360), .IN2(n28461), .IN3(n25307), .IN4(n28457), .Q(
        n25188) );
  OA22X1 U28813 ( .IN1(n25348), .IN2(n28462), .IN3(n25362), .IN4(n28459), .Q(
        n25187) );
  NAND4X0 U28814 ( .IN1(n25190), .IN2(n25189), .IN3(n25188), .IN4(n25187), 
        .QN(s10_data_o[27]) );
  OA22X1 U28815 ( .IN1(n25350), .IN2(n28472), .IN3(n25357), .IN4(n28471), .Q(
        n25194) );
  OA22X1 U28816 ( .IN1(n25348), .IN2(n28474), .IN3(n25347), .IN4(n28473), .Q(
        n25193) );
  OA22X1 U28817 ( .IN1(n25361), .IN2(n28470), .IN3(n25358), .IN4(n28475), .Q(
        n25192) );
  OA22X1 U28818 ( .IN1(n25360), .IN2(n28476), .IN3(n25346), .IN4(n28469), .Q(
        n25191) );
  NAND4X0 U28819 ( .IN1(n25194), .IN2(n25193), .IN3(n25192), .IN4(n25191), 
        .QN(s10_data_o[28]) );
  OA22X1 U28820 ( .IN1(n25358), .IN2(n28483), .IN3(n25347), .IN4(n28481), .Q(
        n25198) );
  OA22X1 U28821 ( .IN1(n25356), .IN2(n28488), .IN3(n25346), .IN4(n28485), .Q(
        n25197) );
  OA22X1 U28822 ( .IN1(n25361), .IN2(n28486), .IN3(n25357), .IN4(n28487), .Q(
        n25196) );
  OA22X1 U28823 ( .IN1(n25348), .IN2(n28484), .IN3(n25360), .IN4(n28482), .Q(
        n25195) );
  NAND4X0 U28824 ( .IN1(n25198), .IN2(n25197), .IN3(n25196), .IN4(n25195), 
        .QN(s10_data_o[29]) );
  OA22X1 U28825 ( .IN1(n25358), .IN2(n28495), .IN3(n25346), .IN4(n28500), .Q(
        n25202) );
  OA22X1 U28826 ( .IN1(n25348), .IN2(n28494), .IN3(n25307), .IN4(n28493), .Q(
        n25201) );
  OA22X1 U28827 ( .IN1(n25350), .IN2(n28497), .IN3(n25340), .IN4(n28496), .Q(
        n25200) );
  OA22X1 U28828 ( .IN1(n25360), .IN2(n28498), .IN3(n25362), .IN4(n28499), .Q(
        n25199) );
  NAND4X0 U28829 ( .IN1(n25202), .IN2(n25201), .IN3(n25200), .IN4(n25199), 
        .QN(s10_data_o[30]) );
  OA22X1 U28830 ( .IN1(n25358), .IN2(n28508), .IN3(n25355), .IN4(n28511), .Q(
        n25206) );
  OA22X1 U28831 ( .IN1(n25359), .IN2(n28510), .IN3(n25350), .IN4(n28506), .Q(
        n25205) );
  OA22X1 U28832 ( .IN1(n25361), .IN2(n28505), .IN3(n25362), .IN4(n28507), .Q(
        n25204) );
  OA22X1 U28833 ( .IN1(n25360), .IN2(n28509), .IN3(n25307), .IN4(n28512), .Q(
        n25203) );
  NAND4X0 U28834 ( .IN1(n25206), .IN2(n25205), .IN3(n25204), .IN4(n25203), 
        .QN(s10_data_o[31]) );
  OA22X1 U28835 ( .IN1(n25359), .IN2(n28518), .IN3(n25345), .IN4(n28520), .Q(
        n25210) );
  OA22X1 U28836 ( .IN1(n25355), .IN2(n28521), .IN3(n25347), .IN4(n28519), .Q(
        n25209) );
  OA22X1 U28837 ( .IN1(n25361), .IN2(n28524), .IN3(n25357), .IN4(n28523), .Q(
        n25208) );
  OA22X1 U28838 ( .IN1(n25349), .IN2(n28517), .IN3(n25350), .IN4(n28522), .Q(
        n25207) );
  NAND4X0 U28839 ( .IN1(n25210), .IN2(n25209), .IN3(n25208), .IN4(n25207), 
        .QN(s10_sel_o[0]) );
  OA22X1 U28840 ( .IN1(n25359), .IN2(n28534), .IN3(n25350), .IN4(n28530), .Q(
        n25214) );
  OA22X1 U28841 ( .IN1(n25357), .IN2(n28535), .IN3(n25362), .IN4(n28529), .Q(
        n25213) );
  OA22X1 U28842 ( .IN1(n25361), .IN2(n28536), .IN3(n25345), .IN4(n28533), .Q(
        n25212) );
  OA22X1 U28843 ( .IN1(n25360), .IN2(n28532), .IN3(n25355), .IN4(n28531), .Q(
        n25211) );
  NAND4X0 U28844 ( .IN1(n25214), .IN2(n25213), .IN3(n25212), .IN4(n25211), 
        .QN(s10_sel_o[1]) );
  OA22X1 U28845 ( .IN1(n25358), .IN2(n28542), .IN3(n25355), .IN4(n28545), .Q(
        n25218) );
  OA22X1 U28846 ( .IN1(n25356), .IN2(n28543), .IN3(n25307), .IN4(n28547), .Q(
        n25217) );
  OA22X1 U28847 ( .IN1(n25359), .IN2(n28544), .IN3(n25340), .IN4(n28548), .Q(
        n25216) );
  OA22X1 U28848 ( .IN1(n25349), .IN2(n28546), .IN3(n25347), .IN4(n28541), .Q(
        n25215) );
  NAND4X0 U28849 ( .IN1(n25218), .IN2(n25217), .IN3(n25216), .IN4(n25215), 
        .QN(s10_sel_o[2]) );
  OA22X1 U28850 ( .IN1(n25359), .IN2(n28558), .IN3(n25355), .IN4(n28559), .Q(
        n25222) );
  OA22X1 U28851 ( .IN1(n25357), .IN2(n28556), .IN3(n25347), .IN4(n28555), .Q(
        n25221) );
  OA22X1 U28852 ( .IN1(n25361), .IN2(n28557), .IN3(n25358), .IN4(n28560), .Q(
        n25220) );
  OA22X1 U28853 ( .IN1(n25360), .IN2(n28554), .IN3(n25356), .IN4(n28553), .Q(
        n25219) );
  NAND4X0 U28854 ( .IN1(n25222), .IN2(n25221), .IN3(n25220), .IN4(n25219), 
        .QN(s10_sel_o[3]) );
  OA22X1 U28855 ( .IN1(n25356), .IN2(n28571), .IN3(n25358), .IN4(n28567), .Q(
        n25226) );
  OA22X1 U28856 ( .IN1(n25361), .IN2(n28566), .IN3(n25355), .IN4(n28565), .Q(
        n25225) );
  OA22X1 U28857 ( .IN1(n25360), .IN2(n28570), .IN3(n25362), .IN4(n28569), .Q(
        n25224) );
  OA22X1 U28858 ( .IN1(n25348), .IN2(n28572), .IN3(n25357), .IN4(n28568), .Q(
        n25223) );
  NAND4X0 U28859 ( .IN1(n25226), .IN2(n25225), .IN3(n25224), .IN4(n25223), 
        .QN(s10_addr_o[0]) );
  OA22X1 U28860 ( .IN1(n25349), .IN2(n28578), .IN3(n25350), .IN4(n28582), .Q(
        n25230) );
  OA22X1 U28861 ( .IN1(n25359), .IN2(n28580), .IN3(n25345), .IN4(n28584), .Q(
        n25229) );
  OA22X1 U28862 ( .IN1(n25355), .IN2(n28577), .IN3(n25362), .IN4(n28583), .Q(
        n25228) );
  OA22X1 U28863 ( .IN1(n25361), .IN2(n28581), .IN3(n25307), .IN4(n28579), .Q(
        n25227) );
  NAND4X0 U28864 ( .IN1(n25230), .IN2(n25229), .IN3(n25228), .IN4(n25227), 
        .QN(s10_addr_o[1]) );
  OA22X1 U28865 ( .IN1(n28592), .IN2(n25340), .IN3(n28593), .IN4(n25345), .Q(
        n25234) );
  OA22X1 U28866 ( .IN1(n28591), .IN2(n25359), .IN3(n28589), .IN4(n25349), .Q(
        n25233) );
  OA22X1 U28867 ( .IN1(n28594), .IN2(n25350), .IN3(n28595), .IN4(n25355), .Q(
        n25232) );
  OA22X1 U28868 ( .IN1(n28596), .IN2(n25347), .IN3(n28590), .IN4(n25307), .Q(
        n25231) );
  NAND4X0 U28869 ( .IN1(n25234), .IN2(n25233), .IN3(n25232), .IN4(n25231), 
        .QN(s10_addr_o[2]) );
  OA22X1 U28870 ( .IN1(n28602), .IN2(n25358), .IN3(n28604), .IN4(n25356), .Q(
        n25238) );
  OA22X1 U28871 ( .IN1(n28606), .IN2(n25307), .IN3(n28605), .IN4(n25349), .Q(
        n25237) );
  OA22X1 U28872 ( .IN1(n28608), .IN2(n25362), .IN3(n28607), .IN4(n25340), .Q(
        n25236) );
  OA22X1 U28873 ( .IN1(n28601), .IN2(n25359), .IN3(n28603), .IN4(n25355), .Q(
        n25235) );
  NAND4X0 U28874 ( .IN1(n25238), .IN2(n25237), .IN3(n25236), .IN4(n25235), 
        .QN(s10_addr_o[3]) );
  OA22X1 U28875 ( .IN1(n28620), .IN2(n25346), .IN3(n28614), .IN4(n25345), .Q(
        n25242) );
  OA22X1 U28876 ( .IN1(n28619), .IN2(n25347), .IN3(n28617), .IN4(n25359), .Q(
        n25241) );
  OA22X1 U28877 ( .IN1(n28616), .IN2(n25349), .IN3(n28615), .IN4(n25357), .Q(
        n25240) );
  OA22X1 U28878 ( .IN1(n28618), .IN2(n25361), .IN3(n28613), .IN4(n25350), .Q(
        n25239) );
  NAND4X0 U28879 ( .IN1(n25242), .IN2(n25241), .IN3(n25240), .IN4(n25239), 
        .QN(s10_addr_o[4]) );
  OA22X1 U28880 ( .IN1(n28632), .IN2(n25356), .IN3(n28629), .IN4(n25359), .Q(
        n25246) );
  OA22X1 U28881 ( .IN1(n28626), .IN2(n25340), .IN3(n28625), .IN4(n25347), .Q(
        n25245) );
  OA22X1 U28882 ( .IN1(n28631), .IN2(n25357), .IN3(n28630), .IN4(n25349), .Q(
        n25244) );
  OA22X1 U28883 ( .IN1(n28628), .IN2(n25346), .IN3(n28627), .IN4(n25345), .Q(
        n25243) );
  NAND4X0 U28884 ( .IN1(n25246), .IN2(n25245), .IN3(n25244), .IN4(n25243), 
        .QN(s10_addr_o[5]) );
  OA22X1 U28885 ( .IN1(n25348), .IN2(n28642), .IN3(n25360), .IN4(n28640), .Q(
        n25250) );
  OA22X1 U28886 ( .IN1(n25357), .IN2(n28638), .IN3(n25347), .IN4(n28639), .Q(
        n25249) );
  OA22X1 U28887 ( .IN1(n25356), .IN2(n28644), .IN3(n25358), .IN4(n28637), .Q(
        n25248) );
  OA22X1 U28888 ( .IN1(n25340), .IN2(n28643), .IN3(n25355), .IN4(n28641), .Q(
        n25247) );
  NAND4X0 U28889 ( .IN1(n25250), .IN2(n25249), .IN3(n25248), .IN4(n25247), 
        .QN(s10_addr_o[6]) );
  OA22X1 U28890 ( .IN1(n25356), .IN2(n28656), .IN3(n25355), .IN4(n28651), .Q(
        n25254) );
  OA22X1 U28891 ( .IN1(n25349), .IN2(n28652), .IN3(n25347), .IN4(n28655), .Q(
        n25253) );
  OA22X1 U28892 ( .IN1(n25359), .IN2(n28654), .IN3(n25357), .IN4(n28650), .Q(
        n25252) );
  OA22X1 U28893 ( .IN1(n25361), .IN2(n28653), .IN3(n25345), .IN4(n28649), .Q(
        n25251) );
  NAND4X0 U28894 ( .IN1(n25254), .IN2(n25253), .IN3(n25252), .IN4(n25251), 
        .QN(s10_addr_o[7]) );
  OA22X1 U28895 ( .IN1(n25359), .IN2(n28664), .IN3(n25347), .IN4(n28667), .Q(
        n25258) );
  OA22X1 U28896 ( .IN1(n25356), .IN2(n28666), .IN3(n25345), .IN4(n28662), .Q(
        n25257) );
  OA22X1 U28897 ( .IN1(n25360), .IN2(n28663), .IN3(n25355), .IN4(n28661), .Q(
        n25256) );
  OA22X1 U28898 ( .IN1(n25361), .IN2(n28665), .IN3(n25307), .IN4(n28668), .Q(
        n25255) );
  NAND4X0 U28899 ( .IN1(n25258), .IN2(n25257), .IN3(n25256), .IN4(n25255), 
        .QN(s10_addr_o[8]) );
  OA22X1 U28900 ( .IN1(n25359), .IN2(n28680), .IN3(n25358), .IN4(n28678), .Q(
        n25262) );
  OA22X1 U28901 ( .IN1(n25361), .IN2(n28676), .IN3(n25355), .IN4(n28675), .Q(
        n25261) );
  OA22X1 U28902 ( .IN1(n25360), .IN2(n28679), .IN3(n25356), .IN4(n28674), .Q(
        n25260) );
  OA22X1 U28903 ( .IN1(n25307), .IN2(n28673), .IN3(n25347), .IN4(n28677), .Q(
        n25259) );
  NAND4X0 U28904 ( .IN1(n25262), .IN2(n25261), .IN3(n25260), .IN4(n25259), 
        .QN(s10_addr_o[9]) );
  OA22X1 U28905 ( .IN1(n25349), .IN2(n28686), .IN3(n25355), .IN4(n28690), .Q(
        n25266) );
  OA22X1 U28906 ( .IN1(n25356), .IN2(n28688), .IN3(n25340), .IN4(n28687), .Q(
        n25265) );
  OA22X1 U28907 ( .IN1(n25348), .IN2(n28692), .IN3(n25307), .IN4(n28685), .Q(
        n25264) );
  OA22X1 U28908 ( .IN1(n25358), .IN2(n28691), .IN3(n25347), .IN4(n28689), .Q(
        n25263) );
  NAND4X0 U28909 ( .IN1(n25266), .IN2(n25265), .IN3(n25264), .IN4(n25263), 
        .QN(s10_addr_o[10]) );
  OA22X1 U28910 ( .IN1(n25356), .IN2(n28697), .IN3(n25355), .IN4(n28700), .Q(
        n25270) );
  OA22X1 U28911 ( .IN1(n25340), .IN2(n28704), .IN3(n25347), .IN4(n28699), .Q(
        n25269) );
  OA22X1 U28912 ( .IN1(n25348), .IN2(n28702), .IN3(n25360), .IN4(n28698), .Q(
        n25268) );
  OA22X1 U28913 ( .IN1(n25357), .IN2(n28701), .IN3(n25358), .IN4(n28703), .Q(
        n25267) );
  NAND4X0 U28914 ( .IN1(n25270), .IN2(n25269), .IN3(n25268), .IN4(n25267), 
        .QN(s10_addr_o[11]) );
  OA22X1 U28915 ( .IN1(n25349), .IN2(n28710), .IN3(n25357), .IN4(n28709), .Q(
        n25274) );
  OA22X1 U28916 ( .IN1(n25356), .IN2(n28712), .IN3(n25340), .IN4(n28716), .Q(
        n25273) );
  OA22X1 U28917 ( .IN1(n25358), .IN2(n28715), .IN3(n25347), .IN4(n28713), .Q(
        n25272) );
  OA22X1 U28918 ( .IN1(n25348), .IN2(n28714), .IN3(n25355), .IN4(n28711), .Q(
        n25271) );
  NAND4X0 U28919 ( .IN1(n25274), .IN2(n25273), .IN3(n25272), .IN4(n25271), 
        .QN(s10_addr_o[12]) );
  OA22X1 U28920 ( .IN1(n25356), .IN2(n28726), .IN3(n25347), .IN4(n28727), .Q(
        n25278) );
  OA22X1 U28921 ( .IN1(n25361), .IN2(n28724), .IN3(n25345), .IN4(n28721), .Q(
        n25277) );
  OA22X1 U28922 ( .IN1(n25359), .IN2(n28722), .IN3(n25360), .IN4(n28728), .Q(
        n25276) );
  OA22X1 U28923 ( .IN1(n25357), .IN2(n28723), .IN3(n25355), .IN4(n28725), .Q(
        n25275) );
  NAND4X0 U28924 ( .IN1(n25278), .IN2(n25277), .IN3(n25276), .IN4(n25275), 
        .QN(s10_addr_o[13]) );
  OA22X1 U28925 ( .IN1(n25340), .IN2(n28735), .IN3(n25355), .IN4(n28733), .Q(
        n25282) );
  OA22X1 U28926 ( .IN1(n25348), .IN2(n28734), .IN3(n25360), .IN4(n28738), .Q(
        n25281) );
  OA22X1 U28927 ( .IN1(n25356), .IN2(n28736), .IN3(n25357), .IN4(n28740), .Q(
        n25280) );
  OA22X1 U28928 ( .IN1(n25358), .IN2(n28737), .IN3(n25347), .IN4(n28739), .Q(
        n25279) );
  NAND4X0 U28929 ( .IN1(n25282), .IN2(n25281), .IN3(n25280), .IN4(n25279), 
        .QN(s10_addr_o[14]) );
  OA22X1 U28930 ( .IN1(n25348), .IN2(n28746), .IN3(n25360), .IN4(n28748), .Q(
        n25286) );
  OA22X1 U28931 ( .IN1(n25361), .IN2(n28752), .IN3(n25307), .IN4(n28747), .Q(
        n25285) );
  OA22X1 U28932 ( .IN1(n25356), .IN2(n28750), .IN3(n25355), .IN4(n28749), .Q(
        n25284) );
  OA22X1 U28933 ( .IN1(n25358), .IN2(n28751), .IN3(n25362), .IN4(n28745), .Q(
        n25283) );
  NAND4X0 U28934 ( .IN1(n25286), .IN2(n25285), .IN3(n25284), .IN4(n25283), 
        .QN(s10_addr_o[15]) );
  OA22X1 U28935 ( .IN1(n25357), .IN2(n28759), .IN3(n25355), .IN4(n28764), .Q(
        n25290) );
  OA22X1 U28936 ( .IN1(n25356), .IN2(n28760), .IN3(n25347), .IN4(n28763), .Q(
        n25289) );
  OA22X1 U28937 ( .IN1(n25349), .IN2(n28762), .IN3(n25340), .IN4(n28761), .Q(
        n25288) );
  OA22X1 U28938 ( .IN1(n25359), .IN2(n28758), .IN3(n25358), .IN4(n28757), .Q(
        n25287) );
  NAND4X0 U28939 ( .IN1(n25290), .IN2(n25289), .IN3(n25288), .IN4(n25287), 
        .QN(s10_addr_o[16]) );
  OA22X1 U28940 ( .IN1(n25356), .IN2(n28774), .IN3(n25345), .IN4(n28771), .Q(
        n25294) );
  OA22X1 U28941 ( .IN1(n25348), .IN2(n28772), .IN3(n25355), .IN4(n28770), .Q(
        n25293) );
  OA22X1 U28942 ( .IN1(n25361), .IN2(n28773), .IN3(n25347), .IN4(n28769), .Q(
        n25292) );
  OA22X1 U28943 ( .IN1(n25360), .IN2(n28776), .IN3(n25357), .IN4(n28775), .Q(
        n25291) );
  NAND4X0 U28944 ( .IN1(n25294), .IN2(n25293), .IN3(n25292), .IN4(n25291), 
        .QN(s10_addr_o[17]) );
  OA22X1 U28945 ( .IN1(n25307), .IN2(n28784), .IN3(n25362), .IN4(n28781), .Q(
        n25298) );
  OA22X1 U28946 ( .IN1(n25358), .IN2(n28783), .IN3(n25355), .IN4(n28785), .Q(
        n25297) );
  OA22X1 U28947 ( .IN1(n25359), .IN2(n28786), .IN3(n25340), .IN4(n28782), .Q(
        n25296) );
  OA22X1 U28948 ( .IN1(n25349), .IN2(n28788), .IN3(n25350), .IN4(n28787), .Q(
        n25295) );
  NAND4X0 U28949 ( .IN1(n25298), .IN2(n25297), .IN3(n25296), .IN4(n25295), 
        .QN(s10_addr_o[18]) );
  OA22X1 U28950 ( .IN1(n25360), .IN2(n28800), .IN3(n25362), .IN4(n28799), .Q(
        n25302) );
  OA22X1 U28951 ( .IN1(n25348), .IN2(n28796), .IN3(n25340), .IN4(n28794), .Q(
        n25301) );
  OA22X1 U28952 ( .IN1(n25357), .IN2(n28797), .IN3(n25345), .IN4(n28795), .Q(
        n25300) );
  OA22X1 U28953 ( .IN1(n25356), .IN2(n28798), .IN3(n25355), .IN4(n28793), .Q(
        n25299) );
  NAND4X0 U28954 ( .IN1(n25302), .IN2(n25301), .IN3(n25300), .IN4(n25299), 
        .QN(s10_addr_o[19]) );
  OA22X1 U28955 ( .IN1(n25356), .IN2(n28807), .IN3(n25355), .IN4(n28809), .Q(
        n25306) );
  OA22X1 U28956 ( .IN1(n25358), .IN2(n28811), .IN3(n25347), .IN4(n28805), .Q(
        n25305) );
  OA22X1 U28957 ( .IN1(n25340), .IN2(n28810), .IN3(n25307), .IN4(n28806), .Q(
        n25304) );
  OA22X1 U28958 ( .IN1(n25359), .IN2(n28812), .IN3(n25360), .IN4(n28808), .Q(
        n25303) );
  NAND4X0 U28959 ( .IN1(n25306), .IN2(n25305), .IN3(n25304), .IN4(n25303), 
        .QN(s10_addr_o[20]) );
  OA22X1 U28960 ( .IN1(n25359), .IN2(n28822), .IN3(n25307), .IN4(n28821), .Q(
        n25311) );
  OA22X1 U28961 ( .IN1(n25350), .IN2(n28820), .IN3(n25347), .IN4(n28817), .Q(
        n25310) );
  OA22X1 U28962 ( .IN1(n25349), .IN2(n28824), .IN3(n25355), .IN4(n28818), .Q(
        n25309) );
  OA22X1 U28963 ( .IN1(n25361), .IN2(n28819), .IN3(n25345), .IN4(n28823), .Q(
        n25308) );
  NAND4X0 U28964 ( .IN1(n25311), .IN2(n25310), .IN3(n25309), .IN4(n25308), 
        .QN(s10_addr_o[21]) );
  OA22X1 U28965 ( .IN1(n25348), .IN2(n28833), .IN3(n25357), .IN4(n28836), .Q(
        n25315) );
  OA22X1 U28966 ( .IN1(n25355), .IN2(n28837), .IN3(n25362), .IN4(n28829), .Q(
        n25314) );
  OA22X1 U28967 ( .IN1(n25356), .IN2(n28831), .IN3(n25345), .IN4(n28834), .Q(
        n25313) );
  OA22X1 U28968 ( .IN1(n25360), .IN2(n28832), .IN3(n25340), .IN4(n28838), .Q(
        n25312) );
  NAND4X0 U28969 ( .IN1(n25315), .IN2(n25314), .IN3(n25313), .IN4(n25312), 
        .QN(s10_addr_o[22]) );
  OA22X1 U28970 ( .IN1(n25361), .IN2(n28850), .IN3(n25345), .IN4(n28849), .Q(
        n25319) );
  OA22X1 U28971 ( .IN1(n25348), .IN2(n28848), .IN3(n25350), .IN4(n28843), .Q(
        n25318) );
  OA22X1 U28972 ( .IN1(n25349), .IN2(n28845), .IN3(n25357), .IN4(n28852), .Q(
        n25317) );
  OA22X1 U28973 ( .IN1(n25355), .IN2(n28846), .IN3(n25347), .IN4(n28851), .Q(
        n25316) );
  NAND4X0 U28974 ( .IN1(n25319), .IN2(n25318), .IN3(n25317), .IN4(n25316), 
        .QN(s10_addr_o[23]) );
  OA22X1 U28975 ( .IN1(n28858), .IN2(n25350), .IN3(n28863), .IN4(n25359), .Q(
        n25323) );
  OA22X1 U28976 ( .IN1(n28857), .IN2(n25361), .IN3(n28861), .IN4(n25357), .Q(
        n25322) );
  OA22X1 U28977 ( .IN1(n28860), .IN2(n25362), .IN3(n28859), .IN4(n25345), .Q(
        n25321) );
  OA22X1 U28978 ( .IN1(n28865), .IN2(n25346), .IN3(n28864), .IN4(n25349), .Q(
        n25320) );
  NAND4X0 U28979 ( .IN1(n25323), .IN2(n25322), .IN3(n25321), .IN4(n25320), 
        .QN(s10_addr_o[24]) );
  OA22X1 U28980 ( .IN1(n28875), .IN2(n25347), .IN3(n28874), .IN4(n25340), .Q(
        n25327) );
  OA22X1 U28981 ( .IN1(n28877), .IN2(n25360), .IN3(n28876), .IN4(n25345), .Q(
        n25326) );
  OA22X1 U28982 ( .IN1(n28871), .IN2(n25346), .IN3(n28872), .IN4(n25357), .Q(
        n25325) );
  OA22X1 U28983 ( .IN1(n28873), .IN2(n25356), .IN3(n28870), .IN4(n25359), .Q(
        n25324) );
  NAND4X0 U28984 ( .IN1(n25327), .IN2(n25326), .IN3(n25325), .IN4(n25324), 
        .QN(s10_addr_o[25]) );
  OA22X1 U28985 ( .IN1(n28889), .IN2(n25362), .IN3(n28882), .IN4(n25340), .Q(
        n25331) );
  OA22X1 U28986 ( .IN1(n28883), .IN2(n25346), .IN3(n28888), .IN4(n25345), .Q(
        n25330) );
  OA22X1 U28987 ( .IN1(n28887), .IN2(n25349), .IN3(n28886), .IN4(n25357), .Q(
        n25329) );
  OA22X1 U28988 ( .IN1(n28885), .IN2(n25350), .IN3(n28884), .IN4(n25359), .Q(
        n25328) );
  NAND4X0 U28989 ( .IN1(n25331), .IN2(n25330), .IN3(n25329), .IN4(n25328), 
        .QN(s10_addr_o[26]) );
  OA22X1 U28990 ( .IN1(n28895), .IN2(n25360), .IN3(n28900), .IN4(n25357), .Q(
        n25335) );
  OA22X1 U28991 ( .IN1(n28898), .IN2(n25347), .IN3(n28901), .IN4(n25361), .Q(
        n25334) );
  OA22X1 U28992 ( .IN1(n28897), .IN2(n25346), .IN3(n28894), .IN4(n25359), .Q(
        n25333) );
  OA22X1 U28993 ( .IN1(n28899), .IN2(n25356), .IN3(n28896), .IN4(n25358), .Q(
        n25332) );
  NAND4X0 U28994 ( .IN1(n25335), .IN2(n25334), .IN3(n25333), .IN4(n25332), 
        .QN(s10_addr_o[27]) );
  OA22X1 U28995 ( .IN1(n28910), .IN2(n25358), .IN3(n28912), .IN4(n25359), .Q(
        n25339) );
  OA22X1 U28996 ( .IN1(n28909), .IN2(n25350), .IN3(n28906), .IN4(n25357), .Q(
        n25338) );
  OA22X1 U28997 ( .IN1(n28907), .IN2(n25346), .IN3(n28913), .IN4(n25362), .Q(
        n25337) );
  OA22X1 U28998 ( .IN1(n28911), .IN2(n25349), .IN3(n28908), .IN4(n25340), .Q(
        n25336) );
  NAND4X0 U28999 ( .IN1(n25339), .IN2(n25338), .IN3(n25337), .IN4(n25336), 
        .QN(s10_addr_o[28]) );
  OA22X1 U29000 ( .IN1(n28920), .IN2(n25358), .IN3(n28923), .IN4(n25357), .Q(
        n25344) );
  OA22X1 U29001 ( .IN1(n28926), .IN2(n25356), .IN3(n28924), .IN4(n25349), .Q(
        n25343) );
  OA22X1 U29002 ( .IN1(n28921), .IN2(n25362), .IN3(n28919), .IN4(n25340), .Q(
        n25342) );
  OA22X1 U29003 ( .IN1(n28922), .IN2(n25346), .IN3(n28925), .IN4(n25359), .Q(
        n25341) );
  NAND4X0 U29004 ( .IN1(n25344), .IN2(n25343), .IN3(n25342), .IN4(n25341), 
        .QN(s10_addr_o[29]) );
  OA22X1 U29005 ( .IN1(n28937), .IN2(n25346), .IN3(n28936), .IN4(n25345), .Q(
        n25354) );
  OA22X1 U29006 ( .IN1(n28933), .IN2(n25347), .IN3(n28939), .IN4(n25357), .Q(
        n25353) );
  OA22X1 U29007 ( .IN1(n28931), .IN2(n25348), .IN3(n28940), .IN4(n25361), .Q(
        n25352) );
  OA22X1 U29008 ( .IN1(n28932), .IN2(n25350), .IN3(n28935), .IN4(n25349), .Q(
        n25351) );
  NAND4X0 U29009 ( .IN1(n25354), .IN2(n25353), .IN3(n25352), .IN4(n25351), 
        .QN(s10_addr_o[30]) );
  OA22X1 U29010 ( .IN1(n28948), .IN2(n25356), .IN3(n28956), .IN4(n25355), .Q(
        n25366) );
  OA22X1 U29011 ( .IN1(n28954), .IN2(n25358), .IN3(n28946), .IN4(n25357), .Q(
        n25365) );
  OA22X1 U29012 ( .IN1(n28952), .IN2(n25360), .IN3(n28950), .IN4(n25359), .Q(
        n25364) );
  OA22X1 U29013 ( .IN1(n28960), .IN2(n25362), .IN3(n28958), .IN4(n25361), .Q(
        n25363) );
  NAND4X0 U29014 ( .IN1(n25366), .IN2(n25365), .IN3(n25364), .IN4(n25363), 
        .QN(s10_addr_o[31]) );
  OA22X1 U29015 ( .IN1(n29368), .IN2(n25368), .IN3(n29311), .IN4(n25367), .Q(
        n25378) );
  OA22X1 U29016 ( .IN1(n29330), .IN2(n25370), .IN3(n29292), .IN4(n25369), .Q(
        n25377) );
  OA22X1 U29017 ( .IN1(n29273), .IN2(n25372), .IN3(n29254), .IN4(n25371), .Q(
        n25376) );
  OA22X1 U29018 ( .IN1(n29349), .IN2(n25374), .IN3(n29235), .IN4(n25373), .Q(
        n25375) );
  NAND4X0 U29019 ( .IN1(n25378), .IN2(n25377), .IN3(n25376), .IN4(n25375), 
        .QN(s9_stb_o) );
  INVX0 U29020 ( .INP(n29130), .ZN(n25652) );
  INVX0 U29021 ( .INP(n29128), .ZN(n25665) );
  OA22X1 U29022 ( .IN1(n25652), .IN2(n28124), .IN3(n25665), .IN4(n28122), .Q(
        n25382) );
  INVX0 U29023 ( .INP(n29127), .ZN(n25641) );
  INVX0 U29024 ( .INP(n29138), .ZN(n25662) );
  OA22X1 U29025 ( .IN1(n25641), .IN2(n28126), .IN3(n25662), .IN4(n28127), .Q(
        n25381) );
  INVX0 U29026 ( .INP(n29137), .ZN(n25659) );
  INVX0 U29027 ( .INP(n25619), .ZN(n29129) );
  INVX0 U29028 ( .INP(n29129), .ZN(n25664) );
  OA22X1 U29029 ( .IN1(n25659), .IN2(n28128), .IN3(n25664), .IN4(n28121), .Q(
        n25380) );
  INVX0 U29030 ( .INP(n29135), .ZN(n25654) );
  INVX0 U29031 ( .INP(n29136), .ZN(n25653) );
  OA22X1 U29032 ( .IN1(n25654), .IN2(n28123), .IN3(n25653), .IN4(n28125), .Q(
        n25379) );
  NAND4X0 U29033 ( .IN1(n25382), .IN2(n25381), .IN3(n25380), .IN4(n25379), 
        .QN(s9_we_o) );
  OA22X1 U29034 ( .IN1(n25652), .IN2(n28134), .IN3(n25662), .IN4(n28137), .Q(
        n25386) );
  INVX0 U29035 ( .INP(n29135), .ZN(n25660) );
  OA22X1 U29036 ( .IN1(n25660), .IN2(n28133), .IN3(n25665), .IN4(n28138), .Q(
        n25385) );
  INVX0 U29037 ( .INP(n29127), .ZN(n25661) );
  OA22X1 U29038 ( .IN1(n25659), .IN2(n28140), .IN3(n25661), .IN4(n28139), .Q(
        n25384) );
  INVX0 U29039 ( .INP(n29136), .ZN(n25663) );
  OA22X1 U29040 ( .IN1(n25663), .IN2(n28136), .IN3(n25619), .IN4(n28135), .Q(
        n25383) );
  NAND4X0 U29041 ( .IN1(n25386), .IN2(n25385), .IN3(n25384), .IN4(n25383), 
        .QN(s9_data_o[0]) );
  OA22X1 U29042 ( .IN1(n25662), .IN2(n28151), .IN3(n25619), .IN4(n28147), .Q(
        n25390) );
  OA22X1 U29043 ( .IN1(n25659), .IN2(n28146), .IN3(n25661), .IN4(n28145), .Q(
        n25389) );
  OA22X1 U29044 ( .IN1(n25654), .IN2(n28148), .IN3(n25663), .IN4(n28152), .Q(
        n25388) );
  OA22X1 U29045 ( .IN1(n25652), .IN2(n28150), .IN3(n25665), .IN4(n28149), .Q(
        n25387) );
  NAND4X0 U29046 ( .IN1(n25390), .IN2(n25389), .IN3(n25388), .IN4(n25387), 
        .QN(s9_data_o[1]) );
  OA22X1 U29047 ( .IN1(n25641), .IN2(n28159), .IN3(n25619), .IN4(n28161), .Q(
        n25394) );
  OA22X1 U29048 ( .IN1(n25659), .IN2(n28164), .IN3(n25665), .IN4(n28158), .Q(
        n25393) );
  OA22X1 U29049 ( .IN1(n25653), .IN2(n28162), .IN3(n25662), .IN4(n28157), .Q(
        n25392) );
  INVX0 U29050 ( .INP(n29130), .ZN(n25666) );
  OA22X1 U29051 ( .IN1(n25666), .IN2(n28160), .IN3(n25654), .IN4(n28163), .Q(
        n25391) );
  NAND4X0 U29052 ( .IN1(n25394), .IN2(n25393), .IN3(n25392), .IN4(n25391), 
        .QN(s9_data_o[2]) );
  OA22X1 U29053 ( .IN1(n25641), .IN2(n28170), .IN3(n25653), .IN4(n28175), .Q(
        n25398) );
  INVX0 U29054 ( .INP(n29128), .ZN(n25651) );
  OA22X1 U29055 ( .IN1(n25651), .IN2(n28171), .IN3(n25619), .IN4(n28173), .Q(
        n25397) );
  OA22X1 U29056 ( .IN1(n25652), .IN2(n28172), .IN3(n25659), .IN4(n28174), .Q(
        n25396) );
  OA22X1 U29057 ( .IN1(n25654), .IN2(n28176), .IN3(n25662), .IN4(n28169), .Q(
        n25395) );
  NAND4X0 U29058 ( .IN1(n25398), .IN2(n25397), .IN3(n25396), .IN4(n25395), 
        .QN(s9_data_o[3]) );
  OA22X1 U29059 ( .IN1(n25660), .IN2(n28186), .IN3(n25653), .IN4(n28183), .Q(
        n25402) );
  OA22X1 U29060 ( .IN1(n25661), .IN2(n28188), .IN3(n25662), .IN4(n28187), .Q(
        n25401) );
  OA22X1 U29061 ( .IN1(n25652), .IN2(n28182), .IN3(n25659), .IN4(n28184), .Q(
        n25400) );
  OA22X1 U29062 ( .IN1(n25665), .IN2(n28185), .IN3(n25619), .IN4(n28181), .Q(
        n25399) );
  NAND4X0 U29063 ( .IN1(n25402), .IN2(n25401), .IN3(n25400), .IN4(n25399), 
        .QN(s9_data_o[4]) );
  INVX0 U29064 ( .INP(n29137), .ZN(n25640) );
  OA22X1 U29065 ( .IN1(n25640), .IN2(n28200), .IN3(n25653), .IN4(n28197), .Q(
        n25406) );
  OA22X1 U29066 ( .IN1(n25651), .IN2(n28198), .IN3(n25619), .IN4(n28199), .Q(
        n25405) );
  OA22X1 U29067 ( .IN1(n25641), .IN2(n28193), .IN3(n25662), .IN4(n28195), .Q(
        n25404) );
  OA22X1 U29068 ( .IN1(n25652), .IN2(n28196), .IN3(n25654), .IN4(n28194), .Q(
        n25403) );
  NAND4X0 U29069 ( .IN1(n25406), .IN2(n25405), .IN3(n25404), .IN4(n25403), 
        .QN(s9_data_o[5]) );
  OA22X1 U29070 ( .IN1(n25659), .IN2(n28207), .IN3(n25661), .IN4(n28212), .Q(
        n25410) );
  OA22X1 U29071 ( .IN1(n25652), .IN2(n28208), .IN3(n25654), .IN4(n28206), .Q(
        n25409) );
  INVX0 U29072 ( .INP(n29138), .ZN(n25650) );
  OA22X1 U29073 ( .IN1(n25650), .IN2(n28210), .IN3(n25619), .IN4(n28209), .Q(
        n25408) );
  OA22X1 U29074 ( .IN1(n25665), .IN2(n28211), .IN3(n25653), .IN4(n28205), .Q(
        n25407) );
  NAND4X0 U29075 ( .IN1(n25410), .IN2(n25409), .IN3(n25408), .IN4(n25407), 
        .QN(s9_data_o[6]) );
  OA22X1 U29076 ( .IN1(n25661), .IN2(n28218), .IN3(n25619), .IN4(n28221), .Q(
        n25414) );
  OA22X1 U29077 ( .IN1(n25640), .IN2(n28219), .IN3(n25653), .IN4(n28223), .Q(
        n25413) );
  OA22X1 U29078 ( .IN1(n25666), .IN2(n28220), .IN3(n25665), .IN4(n28217), .Q(
        n25412) );
  OA22X1 U29079 ( .IN1(n25660), .IN2(n28224), .IN3(n25662), .IN4(n28222), .Q(
        n25411) );
  NAND4X0 U29080 ( .IN1(n25414), .IN2(n25413), .IN3(n25412), .IN4(n25411), 
        .QN(s9_data_o[7]) );
  OA22X1 U29081 ( .IN1(n25662), .IN2(n28233), .IN3(n25664), .IN4(n28235), .Q(
        n25418) );
  OA22X1 U29082 ( .IN1(n25659), .IN2(n28232), .IN3(n25654), .IN4(n28231), .Q(
        n25417) );
  OA22X1 U29083 ( .IN1(n25661), .IN2(n28234), .IN3(n25653), .IN4(n28229), .Q(
        n25416) );
  OA22X1 U29084 ( .IN1(n25666), .IN2(n28230), .IN3(n25665), .IN4(n28236), .Q(
        n25415) );
  NAND4X0 U29085 ( .IN1(n25418), .IN2(n25417), .IN3(n25416), .IN4(n25415), 
        .QN(s9_data_o[8]) );
  OA22X1 U29086 ( .IN1(n25654), .IN2(n28246), .IN3(n25664), .IN4(n28247), .Q(
        n25422) );
  OA22X1 U29087 ( .IN1(n25651), .IN2(n28241), .IN3(n25653), .IN4(n28245), .Q(
        n25421) );
  OA22X1 U29088 ( .IN1(n25652), .IN2(n28242), .IN3(n25659), .IN4(n28244), .Q(
        n25420) );
  OA22X1 U29089 ( .IN1(n25641), .IN2(n28248), .IN3(n25662), .IN4(n28243), .Q(
        n25419) );
  NAND4X0 U29090 ( .IN1(n25422), .IN2(n25421), .IN3(n25420), .IN4(n25419), 
        .QN(s9_data_o[9]) );
  OA22X1 U29091 ( .IN1(n25659), .IN2(n28257), .IN3(n25654), .IN4(n28260), .Q(
        n25426) );
  OA22X1 U29092 ( .IN1(n25666), .IN2(n28258), .IN3(n25661), .IN4(n28256), .Q(
        n25425) );
  OA22X1 U29093 ( .IN1(n25665), .IN2(n28254), .IN3(n25662), .IN4(n28253), .Q(
        n25424) );
  OA22X1 U29094 ( .IN1(n25663), .IN2(n28255), .IN3(n25664), .IN4(n28259), .Q(
        n25423) );
  NAND4X0 U29095 ( .IN1(n25426), .IN2(n25425), .IN3(n25424), .IN4(n25423), 
        .QN(s9_data_o[10]) );
  OA22X1 U29096 ( .IN1(n25640), .IN2(n28272), .IN3(n25661), .IN4(n28271), .Q(
        n25430) );
  OA22X1 U29097 ( .IN1(n25651), .IN2(n28268), .IN3(n25653), .IN4(n28270), .Q(
        n25429) );
  OA22X1 U29098 ( .IN1(n25654), .IN2(n28265), .IN3(n25664), .IN4(n28269), .Q(
        n25428) );
  OA22X1 U29099 ( .IN1(n25652), .IN2(n28266), .IN3(n25662), .IN4(n28267), .Q(
        n25427) );
  NAND4X0 U29100 ( .IN1(n25430), .IN2(n25429), .IN3(n25428), .IN4(n25427), 
        .QN(s9_data_o[11]) );
  OA22X1 U29101 ( .IN1(n25660), .IN2(n28280), .IN3(n25653), .IN4(n28281), .Q(
        n25434) );
  OA22X1 U29102 ( .IN1(n25641), .IN2(n28282), .IN3(n25664), .IN4(n28277), .Q(
        n25433) );
  OA22X1 U29103 ( .IN1(n25640), .IN2(n28278), .IN3(n25665), .IN4(n28283), .Q(
        n25432) );
  OA22X1 U29104 ( .IN1(n25652), .IN2(n28284), .IN3(n25650), .IN4(n28279), .Q(
        n25431) );
  NAND4X0 U29105 ( .IN1(n25434), .IN2(n25433), .IN3(n25432), .IN4(n25431), 
        .QN(s9_data_o[12]) );
  OA22X1 U29106 ( .IN1(n25666), .IN2(n28290), .IN3(n25661), .IN4(n28292), .Q(
        n25438) );
  OA22X1 U29107 ( .IN1(n25663), .IN2(n28293), .IN3(n25650), .IN4(n28291), .Q(
        n25437) );
  OA22X1 U29108 ( .IN1(n25660), .IN2(n28296), .IN3(n25665), .IN4(n28289), .Q(
        n25436) );
  OA22X1 U29109 ( .IN1(n25640), .IN2(n28294), .IN3(n25664), .IN4(n28295), .Q(
        n25435) );
  NAND4X0 U29110 ( .IN1(n25438), .IN2(n25437), .IN3(n25436), .IN4(n25435), 
        .QN(s9_data_o[13]) );
  OA22X1 U29111 ( .IN1(n25652), .IN2(n28306), .IN3(n25650), .IN4(n28301), .Q(
        n25442) );
  OA22X1 U29112 ( .IN1(n25661), .IN2(n28305), .IN3(n25653), .IN4(n28302), .Q(
        n25441) );
  OA22X1 U29113 ( .IN1(n25654), .IN2(n28308), .IN3(n25651), .IN4(n28307), .Q(
        n25440) );
  OA22X1 U29114 ( .IN1(n25640), .IN2(n28304), .IN3(n25664), .IN4(n28303), .Q(
        n25439) );
  NAND4X0 U29115 ( .IN1(n25442), .IN2(n25441), .IN3(n25440), .IN4(n25439), 
        .QN(s9_data_o[14]) );
  OA22X1 U29116 ( .IN1(n25659), .IN2(n28315), .IN3(n25665), .IN4(n28320), .Q(
        n25446) );
  OA22X1 U29117 ( .IN1(n25666), .IN2(n28316), .IN3(n25664), .IN4(n28319), .Q(
        n25445) );
  OA22X1 U29118 ( .IN1(n25661), .IN2(n28313), .IN3(n25650), .IN4(n28317), .Q(
        n25444) );
  OA22X1 U29119 ( .IN1(n25654), .IN2(n28314), .IN3(n25653), .IN4(n28318), .Q(
        n25443) );
  NAND4X0 U29120 ( .IN1(n25446), .IN2(n25445), .IN3(n25444), .IN4(n25443), 
        .QN(s9_data_o[15]) );
  OA22X1 U29121 ( .IN1(n25641), .IN2(n28326), .IN3(n25664), .IN4(n28327), .Q(
        n25450) );
  OA22X1 U29122 ( .IN1(n25652), .IN2(n28330), .IN3(n25653), .IN4(n28325), .Q(
        n25449) );
  OA22X1 U29123 ( .IN1(n25640), .IN2(n28332), .IN3(n25654), .IN4(n28331), .Q(
        n25448) );
  OA22X1 U29124 ( .IN1(n25665), .IN2(n28329), .IN3(n25650), .IN4(n28328), .Q(
        n25447) );
  NAND4X0 U29125 ( .IN1(n25450), .IN2(n25449), .IN3(n25448), .IN4(n25447), 
        .QN(s9_data_o[16]) );
  OA22X1 U29126 ( .IN1(n25654), .IN2(n28342), .IN3(n25653), .IN4(n28339), .Q(
        n25454) );
  OA22X1 U29127 ( .IN1(n25659), .IN2(n28344), .IN3(n25651), .IN4(n28337), .Q(
        n25453) );
  OA22X1 U29128 ( .IN1(n25652), .IN2(n28340), .IN3(n25641), .IN4(n28338), .Q(
        n25452) );
  OA22X1 U29129 ( .IN1(n25662), .IN2(n28343), .IN3(n25664), .IN4(n28341), .Q(
        n25451) );
  NAND4X0 U29130 ( .IN1(n25454), .IN2(n25453), .IN3(n25452), .IN4(n25451), 
        .QN(s9_data_o[17]) );
  OA22X1 U29131 ( .IN1(n25650), .IN2(n28351), .IN3(n25664), .IN4(n28353), .Q(
        n25458) );
  OA22X1 U29132 ( .IN1(n25654), .IN2(n28350), .IN3(n25651), .IN4(n28354), .Q(
        n25457) );
  OA22X1 U29133 ( .IN1(n25666), .IN2(n28352), .IN3(n25653), .IN4(n28349), .Q(
        n25456) );
  OA22X1 U29134 ( .IN1(n25659), .IN2(n28356), .IN3(n25641), .IN4(n28355), .Q(
        n25455) );
  NAND4X0 U29135 ( .IN1(n25458), .IN2(n25457), .IN3(n25456), .IN4(n25455), 
        .QN(s9_data_o[18]) );
  OA22X1 U29136 ( .IN1(n25652), .IN2(n28366), .IN3(n25665), .IN4(n28365), .Q(
        n25462) );
  OA22X1 U29137 ( .IN1(n25640), .IN2(n28364), .IN3(n25653), .IN4(n28361), .Q(
        n25461) );
  OA22X1 U29138 ( .IN1(n25662), .IN2(n28368), .IN3(n25664), .IN4(n28367), .Q(
        n25460) );
  OA22X1 U29139 ( .IN1(n25654), .IN2(n28362), .IN3(n25661), .IN4(n28363), .Q(
        n25459) );
  NAND4X0 U29140 ( .IN1(n25462), .IN2(n25461), .IN3(n25460), .IN4(n25459), 
        .QN(s9_data_o[19]) );
  OA22X1 U29141 ( .IN1(n25662), .IN2(n28379), .IN3(n25664), .IN4(n28375), .Q(
        n25466) );
  OA22X1 U29142 ( .IN1(n25666), .IN2(n28378), .IN3(n25659), .IN4(n28377), .Q(
        n25465) );
  OA22X1 U29143 ( .IN1(n25661), .IN2(n28373), .IN3(n25653), .IN4(n28380), .Q(
        n25464) );
  OA22X1 U29144 ( .IN1(n25660), .IN2(n28374), .IN3(n25665), .IN4(n28376), .Q(
        n25463) );
  NAND4X0 U29145 ( .IN1(n25466), .IN2(n25465), .IN3(n25464), .IN4(n25463), 
        .QN(s9_data_o[20]) );
  OA22X1 U29146 ( .IN1(n25640), .IN2(n28386), .IN3(n25651), .IN4(n28387), .Q(
        n25470) );
  OA22X1 U29147 ( .IN1(n25663), .IN2(n28385), .IN3(n25650), .IN4(n28389), .Q(
        n25469) );
  OA22X1 U29148 ( .IN1(n25652), .IN2(n28392), .IN3(n25664), .IN4(n28391), .Q(
        n25468) );
  OA22X1 U29149 ( .IN1(n25654), .IN2(n28390), .IN3(n25661), .IN4(n28388), .Q(
        n25467) );
  NAND4X0 U29150 ( .IN1(n25470), .IN2(n25469), .IN3(n25468), .IN4(n25467), 
        .QN(s9_data_o[21]) );
  OA22X1 U29151 ( .IN1(n25652), .IN2(n28400), .IN3(n25661), .IN4(n28403), .Q(
        n25474) );
  OA22X1 U29152 ( .IN1(n25659), .IN2(n28402), .IN3(n25665), .IN4(n28398), .Q(
        n25473) );
  OA22X1 U29153 ( .IN1(n25660), .IN2(n28404), .IN3(n25664), .IN4(n28397), .Q(
        n25472) );
  OA22X1 U29154 ( .IN1(n25663), .IN2(n28399), .IN3(n25650), .IN4(n28401), .Q(
        n25471) );
  NAND4X0 U29155 ( .IN1(n25474), .IN2(n25473), .IN3(n25472), .IN4(n25471), 
        .QN(s9_data_o[22]) );
  OA22X1 U29156 ( .IN1(n25660), .IN2(n28414), .IN3(n25663), .IN4(n28412), .Q(
        n25478) );
  OA22X1 U29157 ( .IN1(n25640), .IN2(n28415), .IN3(n25641), .IN4(n28413), .Q(
        n25477) );
  OA22X1 U29158 ( .IN1(n25662), .IN2(n28409), .IN3(n25664), .IN4(n28411), .Q(
        n25476) );
  OA22X1 U29159 ( .IN1(n25652), .IN2(n28416), .IN3(n25651), .IN4(n28410), .Q(
        n25475) );
  NAND4X0 U29160 ( .IN1(n25478), .IN2(n25477), .IN3(n25476), .IN4(n25475), 
        .QN(s9_data_o[23]) );
  OA22X1 U29161 ( .IN1(n25662), .IN2(n28427), .IN3(n25619), .IN4(n28423), .Q(
        n25482) );
  OA22X1 U29162 ( .IN1(n25641), .IN2(n28421), .IN3(n25663), .IN4(n28428), .Q(
        n25481) );
  OA22X1 U29163 ( .IN1(n25659), .IN2(n28424), .IN3(n25654), .IN4(n28422), .Q(
        n25480) );
  OA22X1 U29164 ( .IN1(n25666), .IN2(n28426), .IN3(n25651), .IN4(n28425), .Q(
        n25479) );
  NAND4X0 U29165 ( .IN1(n25482), .IN2(n25481), .IN3(n25480), .IN4(n25479), 
        .QN(s9_data_o[24]) );
  OA22X1 U29166 ( .IN1(n25661), .IN2(n28439), .IN3(n25653), .IN4(n28437), .Q(
        n25486) );
  OA22X1 U29167 ( .IN1(n25666), .IN2(n28438), .IN3(n25654), .IN4(n28434), .Q(
        n25485) );
  OA22X1 U29168 ( .IN1(n25659), .IN2(n28440), .IN3(n25619), .IN4(n28435), .Q(
        n25484) );
  OA22X1 U29169 ( .IN1(n25651), .IN2(n28433), .IN3(n25650), .IN4(n28436), .Q(
        n25483) );
  NAND4X0 U29170 ( .IN1(n25486), .IN2(n25485), .IN3(n25484), .IN4(n25483), 
        .QN(s9_data_o[25]) );
  OA22X1 U29171 ( .IN1(n25663), .IN2(n28448), .IN3(n25619), .IN4(n28445), .Q(
        n25490) );
  OA22X1 U29172 ( .IN1(n25666), .IN2(n28452), .IN3(n25641), .IN4(n28446), .Q(
        n25489) );
  OA22X1 U29173 ( .IN1(n25640), .IN2(n28451), .IN3(n25665), .IN4(n28449), .Q(
        n25488) );
  OA22X1 U29174 ( .IN1(n25654), .IN2(n28450), .IN3(n25650), .IN4(n28447), .Q(
        n25487) );
  NAND4X0 U29175 ( .IN1(n25490), .IN2(n25489), .IN3(n25488), .IN4(n25487), 
        .QN(s9_data_o[26]) );
  OA22X1 U29176 ( .IN1(n25652), .IN2(n28462), .IN3(n25661), .IN4(n28458), .Q(
        n25494) );
  OA22X1 U29177 ( .IN1(n25654), .IN2(n28464), .IN3(n25665), .IN4(n28457), .Q(
        n25493) );
  OA22X1 U29178 ( .IN1(n25662), .IN2(n28460), .IN3(n25619), .IN4(n28459), .Q(
        n25492) );
  OA22X1 U29179 ( .IN1(n25659), .IN2(n28461), .IN3(n25663), .IN4(n28463), .Q(
        n25491) );
  NAND4X0 U29180 ( .IN1(n25494), .IN2(n25493), .IN3(n25492), .IN4(n25491), 
        .QN(s9_data_o[27]) );
  OA22X1 U29181 ( .IN1(n25666), .IN2(n28474), .IN3(n25665), .IN4(n28471), .Q(
        n25498) );
  OA22X1 U29182 ( .IN1(n25640), .IN2(n28476), .IN3(n25641), .IN4(n28470), .Q(
        n25497) );
  OA22X1 U29183 ( .IN1(n25660), .IN2(n28472), .IN3(n25650), .IN4(n28469), .Q(
        n25496) );
  OA22X1 U29184 ( .IN1(n25663), .IN2(n28475), .IN3(n25619), .IN4(n28473), .Q(
        n25495) );
  NAND4X0 U29185 ( .IN1(n25498), .IN2(n25497), .IN3(n25496), .IN4(n25495), 
        .QN(s9_data_o[28]) );
  OA22X1 U29186 ( .IN1(n25641), .IN2(n28486), .IN3(n25650), .IN4(n28485), .Q(
        n25502) );
  OA22X1 U29187 ( .IN1(n25652), .IN2(n28484), .IN3(n25651), .IN4(n28487), .Q(
        n25501) );
  OA22X1 U29188 ( .IN1(n25659), .IN2(n28482), .IN3(n25619), .IN4(n28481), .Q(
        n25500) );
  OA22X1 U29189 ( .IN1(n25654), .IN2(n28488), .IN3(n25663), .IN4(n28483), .Q(
        n25499) );
  NAND4X0 U29190 ( .IN1(n25502), .IN2(n25501), .IN3(n25500), .IN4(n25499), 
        .QN(s9_data_o[29]) );
  OA22X1 U29191 ( .IN1(n25660), .IN2(n28497), .IN3(n25641), .IN4(n28496), .Q(
        n25506) );
  OA22X1 U29192 ( .IN1(n25640), .IN2(n28498), .IN3(n25653), .IN4(n28495), .Q(
        n25505) );
  OA22X1 U29193 ( .IN1(n25651), .IN2(n28493), .IN3(n25650), .IN4(n28500), .Q(
        n25504) );
  OA22X1 U29194 ( .IN1(n25666), .IN2(n28494), .IN3(n25619), .IN4(n28499), .Q(
        n25503) );
  NAND4X0 U29195 ( .IN1(n25506), .IN2(n25505), .IN3(n25504), .IN4(n25503), 
        .QN(s9_data_o[30]) );
  OA22X1 U29196 ( .IN1(n25660), .IN2(n28506), .IN3(n25650), .IN4(n28511), .Q(
        n25510) );
  OA22X1 U29197 ( .IN1(n25659), .IN2(n28509), .IN3(n25653), .IN4(n28508), .Q(
        n25509) );
  OA22X1 U29198 ( .IN1(n25661), .IN2(n28505), .IN3(n25619), .IN4(n28507), .Q(
        n25508) );
  OA22X1 U29199 ( .IN1(n25666), .IN2(n28510), .IN3(n25651), .IN4(n28512), .Q(
        n25507) );
  NAND4X0 U29200 ( .IN1(n25510), .IN2(n25509), .IN3(n25508), .IN4(n25507), 
        .QN(s9_data_o[31]) );
  OA22X1 U29201 ( .IN1(n25651), .IN2(n28523), .IN3(n25663), .IN4(n28520), .Q(
        n25514) );
  OA22X1 U29202 ( .IN1(n25641), .IN2(n28524), .IN3(n25619), .IN4(n28519), .Q(
        n25513) );
  OA22X1 U29203 ( .IN1(n25666), .IN2(n28518), .IN3(n25650), .IN4(n28521), .Q(
        n25512) );
  OA22X1 U29204 ( .IN1(n25640), .IN2(n28517), .IN3(n25654), .IN4(n28522), .Q(
        n25511) );
  NAND4X0 U29205 ( .IN1(n25514), .IN2(n25513), .IN3(n25512), .IN4(n25511), 
        .QN(s9_sel_o[0]) );
  OA22X1 U29206 ( .IN1(n25660), .IN2(n28530), .IN3(n25661), .IN4(n28536), .Q(
        n25518) );
  OA22X1 U29207 ( .IN1(n25651), .IN2(n28535), .IN3(n25663), .IN4(n28533), .Q(
        n25517) );
  OA22X1 U29208 ( .IN1(n25666), .IN2(n28534), .IN3(n25619), .IN4(n28529), .Q(
        n25516) );
  OA22X1 U29209 ( .IN1(n25659), .IN2(n28532), .IN3(n25650), .IN4(n28531), .Q(
        n25515) );
  NAND4X0 U29210 ( .IN1(n25518), .IN2(n25517), .IN3(n25516), .IN4(n25515), 
        .QN(s9_sel_o[1]) );
  OA22X1 U29211 ( .IN1(n25661), .IN2(n28548), .IN3(n25665), .IN4(n28547), .Q(
        n25522) );
  OA22X1 U29212 ( .IN1(n25666), .IN2(n28544), .IN3(n25659), .IN4(n28546), .Q(
        n25521) );
  OA22X1 U29213 ( .IN1(n25660), .IN2(n28543), .IN3(n25653), .IN4(n28542), .Q(
        n25520) );
  OA22X1 U29214 ( .IN1(n25662), .IN2(n28545), .IN3(n25619), .IN4(n28541), .Q(
        n25519) );
  NAND4X0 U29215 ( .IN1(n25522), .IN2(n25521), .IN3(n25520), .IN4(n25519), 
        .QN(s9_sel_o[2]) );
  OA22X1 U29216 ( .IN1(n25666), .IN2(n28558), .IN3(n25619), .IN4(n28555), .Q(
        n25526) );
  OA22X1 U29217 ( .IN1(n25660), .IN2(n28553), .IN3(n25661), .IN4(n28557), .Q(
        n25525) );
  OA22X1 U29218 ( .IN1(n25640), .IN2(n28554), .IN3(n25665), .IN4(n28556), .Q(
        n25524) );
  OA22X1 U29219 ( .IN1(n25663), .IN2(n28560), .IN3(n25650), .IN4(n28559), .Q(
        n25523) );
  NAND4X0 U29220 ( .IN1(n25526), .IN2(n25525), .IN3(n25524), .IN4(n25523), 
        .QN(s9_sel_o[3]) );
  OA22X1 U29221 ( .IN1(n25666), .IN2(n28572), .IN3(n25659), .IN4(n28570), .Q(
        n25530) );
  OA22X1 U29222 ( .IN1(n25641), .IN2(n28566), .IN3(n25619), .IN4(n28569), .Q(
        n25529) );
  OA22X1 U29223 ( .IN1(n25663), .IN2(n28567), .IN3(n25650), .IN4(n28565), .Q(
        n25528) );
  OA22X1 U29224 ( .IN1(n25660), .IN2(n28571), .IN3(n25651), .IN4(n28568), .Q(
        n25527) );
  NAND4X0 U29225 ( .IN1(n25530), .IN2(n25529), .IN3(n25528), .IN4(n25527), 
        .QN(s9_addr_o[0]) );
  OA22X1 U29226 ( .IN1(n25660), .IN2(n28582), .IN3(n25619), .IN4(n28583), .Q(
        n25534) );
  OA22X1 U29227 ( .IN1(n25661), .IN2(n28581), .IN3(n25663), .IN4(n28584), .Q(
        n25533) );
  OA22X1 U29228 ( .IN1(n25651), .IN2(n28579), .IN3(n25650), .IN4(n28577), .Q(
        n25532) );
  OA22X1 U29229 ( .IN1(n25666), .IN2(n28580), .IN3(n25659), .IN4(n28578), .Q(
        n25531) );
  NAND4X0 U29230 ( .IN1(n25534), .IN2(n25533), .IN3(n25532), .IN4(n25531), 
        .QN(s9_addr_o[1]) );
  OA22X1 U29231 ( .IN1(n28594), .IN2(n25660), .IN3(n28589), .IN4(n25640), .Q(
        n25538) );
  OA22X1 U29232 ( .IN1(n28596), .IN2(n25664), .IN3(n28590), .IN4(n25665), .Q(
        n25537) );
  OA22X1 U29233 ( .IN1(n28591), .IN2(n25652), .IN3(n28595), .IN4(n25650), .Q(
        n25536) );
  OA22X1 U29234 ( .IN1(n28592), .IN2(n25641), .IN3(n28593), .IN4(n25653), .Q(
        n25535) );
  NAND4X0 U29235 ( .IN1(n25538), .IN2(n25537), .IN3(n25536), .IN4(n25535), 
        .QN(s9_addr_o[2]) );
  OA22X1 U29236 ( .IN1(n28605), .IN2(n25640), .IN3(n28608), .IN4(n25664), .Q(
        n25542) );
  OA22X1 U29237 ( .IN1(n28606), .IN2(n25665), .IN3(n28603), .IN4(n25650), .Q(
        n25541) );
  OA22X1 U29238 ( .IN1(n28602), .IN2(n25653), .IN3(n28607), .IN4(n25661), .Q(
        n25540) );
  OA22X1 U29239 ( .IN1(n28604), .IN2(n25654), .IN3(n28601), .IN4(n25652), .Q(
        n25539) );
  NAND4X0 U29240 ( .IN1(n25542), .IN2(n25541), .IN3(n25540), .IN4(n25539), 
        .QN(s9_addr_o[3]) );
  OA22X1 U29241 ( .IN1(n28614), .IN2(n25663), .IN3(n28613), .IN4(n25660), .Q(
        n25546) );
  OA22X1 U29242 ( .IN1(n28618), .IN2(n25641), .IN3(n28617), .IN4(n25652), .Q(
        n25545) );
  OA22X1 U29243 ( .IN1(n28616), .IN2(n25640), .IN3(n28620), .IN4(n25650), .Q(
        n25544) );
  OA22X1 U29244 ( .IN1(n28619), .IN2(n25664), .IN3(n28615), .IN4(n25665), .Q(
        n25543) );
  NAND4X0 U29245 ( .IN1(n25546), .IN2(n25545), .IN3(n25544), .IN4(n25543), 
        .QN(s9_addr_o[4]) );
  OA22X1 U29246 ( .IN1(n28627), .IN2(n25653), .IN3(n28631), .IN4(n25665), .Q(
        n25550) );
  OA22X1 U29247 ( .IN1(n28626), .IN2(n25641), .IN3(n28630), .IN4(n25659), .Q(
        n25549) );
  OA22X1 U29248 ( .IN1(n28632), .IN2(n25660), .IN3(n28625), .IN4(n25664), .Q(
        n25548) );
  OA22X1 U29249 ( .IN1(n28628), .IN2(n25650), .IN3(n28629), .IN4(n25652), .Q(
        n25547) );
  NAND4X0 U29250 ( .IN1(n25550), .IN2(n25549), .IN3(n25548), .IN4(n25547), 
        .QN(s9_addr_o[5]) );
  OA22X1 U29251 ( .IN1(n25663), .IN2(n28637), .IN3(n25619), .IN4(n28639), .Q(
        n25554) );
  OA22X1 U29252 ( .IN1(n25651), .IN2(n28638), .IN3(n25662), .IN4(n28641), .Q(
        n25553) );
  OA22X1 U29253 ( .IN1(n25659), .IN2(n28640), .IN3(n25654), .IN4(n28644), .Q(
        n25552) );
  OA22X1 U29254 ( .IN1(n25666), .IN2(n28642), .IN3(n25661), .IN4(n28643), .Q(
        n25551) );
  NAND4X0 U29255 ( .IN1(n25554), .IN2(n25553), .IN3(n25552), .IN4(n25551), 
        .QN(s9_addr_o[6]) );
  OA22X1 U29256 ( .IN1(n25660), .IN2(n28656), .IN3(n25650), .IN4(n28651), .Q(
        n25558) );
  OA22X1 U29257 ( .IN1(n25666), .IN2(n28654), .IN3(n25653), .IN4(n28649), .Q(
        n25557) );
  OA22X1 U29258 ( .IN1(n25640), .IN2(n28652), .IN3(n25651), .IN4(n28650), .Q(
        n25556) );
  OA22X1 U29259 ( .IN1(n25641), .IN2(n28653), .IN3(n25619), .IN4(n28655), .Q(
        n25555) );
  NAND4X0 U29260 ( .IN1(n25558), .IN2(n25557), .IN3(n25556), .IN4(n25555), 
        .QN(s9_addr_o[7]) );
  OA22X1 U29261 ( .IN1(n25666), .IN2(n28664), .IN3(n25661), .IN4(n28665), .Q(
        n25562) );
  OA22X1 U29262 ( .IN1(n25651), .IN2(n28668), .IN3(n25662), .IN4(n28661), .Q(
        n25561) );
  OA22X1 U29263 ( .IN1(n25659), .IN2(n28663), .IN3(n25654), .IN4(n28666), .Q(
        n25560) );
  OA22X1 U29264 ( .IN1(n25653), .IN2(n28662), .IN3(n25619), .IN4(n28667), .Q(
        n25559) );
  NAND4X0 U29265 ( .IN1(n25562), .IN2(n25561), .IN3(n25560), .IN4(n25559), 
        .QN(s9_addr_o[8]) );
  OA22X1 U29266 ( .IN1(n25651), .IN2(n28673), .IN3(n25662), .IN4(n28675), .Q(
        n25566) );
  OA22X1 U29267 ( .IN1(n25661), .IN2(n28676), .IN3(n25663), .IN4(n28678), .Q(
        n25565) );
  OA22X1 U29268 ( .IN1(n25660), .IN2(n28674), .IN3(n25619), .IN4(n28677), .Q(
        n25564) );
  OA22X1 U29269 ( .IN1(n25666), .IN2(n28680), .IN3(n25659), .IN4(n28679), .Q(
        n25563) );
  NAND4X0 U29270 ( .IN1(n25566), .IN2(n25565), .IN3(n25564), .IN4(n25563), 
        .QN(s9_addr_o[9]) );
  OA22X1 U29271 ( .IN1(n25666), .IN2(n28692), .IN3(n25654), .IN4(n28688), .Q(
        n25570) );
  OA22X1 U29272 ( .IN1(n25651), .IN2(n28685), .IN3(n25653), .IN4(n28691), .Q(
        n25569) );
  OA22X1 U29273 ( .IN1(n25641), .IN2(n28687), .IN3(n25619), .IN4(n28689), .Q(
        n25568) );
  OA22X1 U29274 ( .IN1(n25640), .IN2(n28686), .IN3(n25650), .IN4(n28690), .Q(
        n25567) );
  NAND4X0 U29275 ( .IN1(n25570), .IN2(n25569), .IN3(n25568), .IN4(n25567), 
        .QN(s9_addr_o[10]) );
  OA22X1 U29276 ( .IN1(n25666), .IN2(n28702), .IN3(n25665), .IN4(n28701), .Q(
        n25574) );
  OA22X1 U29277 ( .IN1(n25641), .IN2(n28704), .IN3(n25653), .IN4(n28703), .Q(
        n25573) );
  OA22X1 U29278 ( .IN1(n25659), .IN2(n28698), .IN3(n25650), .IN4(n28700), .Q(
        n25572) );
  OA22X1 U29279 ( .IN1(n25660), .IN2(n28697), .IN3(n25619), .IN4(n28699), .Q(
        n25571) );
  NAND4X0 U29280 ( .IN1(n25574), .IN2(n25573), .IN3(n25572), .IN4(n25571), 
        .QN(s9_addr_o[11]) );
  OA22X1 U29281 ( .IN1(n25641), .IN2(n28716), .IN3(n25663), .IN4(n28715), .Q(
        n25578) );
  OA22X1 U29282 ( .IN1(n25660), .IN2(n28712), .IN3(n25665), .IN4(n28709), .Q(
        n25577) );
  OA22X1 U29283 ( .IN1(n25666), .IN2(n28714), .IN3(n25659), .IN4(n28710), .Q(
        n25576) );
  OA22X1 U29284 ( .IN1(n25662), .IN2(n28711), .IN3(n25619), .IN4(n28713), .Q(
        n25575) );
  NAND4X0 U29285 ( .IN1(n25578), .IN2(n25577), .IN3(n25576), .IN4(n25575), 
        .QN(s9_addr_o[12]) );
  OA22X1 U29286 ( .IN1(n25652), .IN2(n28722), .IN3(n25619), .IN4(n28727), .Q(
        n25582) );
  OA22X1 U29287 ( .IN1(n25651), .IN2(n28723), .IN3(n25663), .IN4(n28721), .Q(
        n25581) );
  OA22X1 U29288 ( .IN1(n25640), .IN2(n28728), .IN3(n25654), .IN4(n28726), .Q(
        n25580) );
  OA22X1 U29289 ( .IN1(n25641), .IN2(n28724), .IN3(n25662), .IN4(n28725), .Q(
        n25579) );
  NAND4X0 U29290 ( .IN1(n25582), .IN2(n25581), .IN3(n25580), .IN4(n25579), 
        .QN(s9_addr_o[13]) );
  OA22X1 U29291 ( .IN1(n25665), .IN2(n28740), .IN3(n25650), .IN4(n28733), .Q(
        n25586) );
  OA22X1 U29292 ( .IN1(n25641), .IN2(n28735), .IN3(n25653), .IN4(n28737), .Q(
        n25585) );
  OA22X1 U29293 ( .IN1(n25640), .IN2(n28738), .IN3(n25654), .IN4(n28736), .Q(
        n25584) );
  OA22X1 U29294 ( .IN1(n25666), .IN2(n28734), .IN3(n25619), .IN4(n28739), .Q(
        n25583) );
  NAND4X0 U29295 ( .IN1(n25586), .IN2(n25585), .IN3(n25584), .IN4(n25583), 
        .QN(s9_addr_o[14]) );
  OA22X1 U29296 ( .IN1(n25651), .IN2(n28747), .IN3(n25663), .IN4(n28751), .Q(
        n25590) );
  OA22X1 U29297 ( .IN1(n25640), .IN2(n28748), .IN3(n25619), .IN4(n28745), .Q(
        n25589) );
  OA22X1 U29298 ( .IN1(n25666), .IN2(n28746), .IN3(n25661), .IN4(n28752), .Q(
        n25588) );
  OA22X1 U29299 ( .IN1(n25660), .IN2(n28750), .IN3(n25662), .IN4(n28749), .Q(
        n25587) );
  NAND4X0 U29300 ( .IN1(n25590), .IN2(n25589), .IN3(n25588), .IN4(n25587), 
        .QN(s9_addr_o[15]) );
  OA22X1 U29301 ( .IN1(n25641), .IN2(n28761), .IN3(n25662), .IN4(n28764), .Q(
        n25594) );
  OA22X1 U29302 ( .IN1(n25652), .IN2(n28758), .IN3(n25654), .IN4(n28760), .Q(
        n25593) );
  OA22X1 U29303 ( .IN1(n25640), .IN2(n28762), .IN3(n25651), .IN4(n28759), .Q(
        n25592) );
  OA22X1 U29304 ( .IN1(n25663), .IN2(n28757), .IN3(n25619), .IN4(n28763), .Q(
        n25591) );
  NAND4X0 U29305 ( .IN1(n25594), .IN2(n25593), .IN3(n25592), .IN4(n25591), 
        .QN(s9_addr_o[16]) );
  OA22X1 U29306 ( .IN1(n25666), .IN2(n28772), .IN3(n25659), .IN4(n28776), .Q(
        n25598) );
  OA22X1 U29307 ( .IN1(n25641), .IN2(n28773), .IN3(n25665), .IN4(n28775), .Q(
        n25597) );
  OA22X1 U29308 ( .IN1(n25660), .IN2(n28774), .IN3(n25653), .IN4(n28771), .Q(
        n25596) );
  OA22X1 U29309 ( .IN1(n25650), .IN2(n28770), .IN3(n25619), .IN4(n28769), .Q(
        n25595) );
  NAND4X0 U29310 ( .IN1(n25598), .IN2(n25597), .IN3(n25596), .IN4(n25595), 
        .QN(s9_addr_o[17]) );
  OA22X1 U29311 ( .IN1(n25651), .IN2(n28784), .IN3(n25650), .IN4(n28785), .Q(
        n25602) );
  OA22X1 U29312 ( .IN1(n25661), .IN2(n28782), .IN3(n25619), .IN4(n28781), .Q(
        n25601) );
  OA22X1 U29313 ( .IN1(n25640), .IN2(n28788), .IN3(n25654), .IN4(n28787), .Q(
        n25600) );
  OA22X1 U29314 ( .IN1(n25652), .IN2(n28786), .IN3(n25653), .IN4(n28783), .Q(
        n25599) );
  NAND4X0 U29315 ( .IN1(n25602), .IN2(n25601), .IN3(n25600), .IN4(n25599), 
        .QN(s9_addr_o[18]) );
  OA22X1 U29316 ( .IN1(n25660), .IN2(n28798), .IN3(n25619), .IN4(n28799), .Q(
        n25606) );
  OA22X1 U29317 ( .IN1(n25640), .IN2(n28800), .IN3(n25661), .IN4(n28794), .Q(
        n25605) );
  OA22X1 U29318 ( .IN1(n25665), .IN2(n28797), .IN3(n25650), .IN4(n28793), .Q(
        n25604) );
  OA22X1 U29319 ( .IN1(n25666), .IN2(n28796), .IN3(n25663), .IN4(n28795), .Q(
        n25603) );
  NAND4X0 U29320 ( .IN1(n25606), .IN2(n25605), .IN3(n25604), .IN4(n25603), 
        .QN(s9_addr_o[19]) );
  OA22X1 U29321 ( .IN1(n25652), .IN2(n28812), .IN3(n25619), .IN4(n28805), .Q(
        n25610) );
  OA22X1 U29322 ( .IN1(n25641), .IN2(n28810), .IN3(n25651), .IN4(n28806), .Q(
        n25609) );
  OA22X1 U29323 ( .IN1(n25663), .IN2(n28811), .IN3(n25662), .IN4(n28809), .Q(
        n25608) );
  OA22X1 U29324 ( .IN1(n25640), .IN2(n28808), .IN3(n25654), .IN4(n28807), .Q(
        n25607) );
  NAND4X0 U29325 ( .IN1(n25610), .IN2(n25609), .IN3(n25608), .IN4(n25607), 
        .QN(s9_addr_o[20]) );
  OA22X1 U29326 ( .IN1(n25651), .IN2(n28821), .IN3(n25662), .IN4(n28818), .Q(
        n25614) );
  OA22X1 U29327 ( .IN1(n25666), .IN2(n28822), .IN3(n25661), .IN4(n28819), .Q(
        n25613) );
  OA22X1 U29328 ( .IN1(n25640), .IN2(n28824), .IN3(n25619), .IN4(n28817), .Q(
        n25612) );
  OA22X1 U29329 ( .IN1(n25660), .IN2(n28820), .IN3(n25663), .IN4(n28823), .Q(
        n25611) );
  NAND4X0 U29330 ( .IN1(n25614), .IN2(n25613), .IN3(n25612), .IN4(n25611), 
        .QN(s9_addr_o[21]) );
  OA22X1 U29331 ( .IN1(n25640), .IN2(n28832), .IN3(n25661), .IN4(n28838), .Q(
        n25618) );
  OA22X1 U29332 ( .IN1(n25660), .IN2(n28831), .IN3(n25651), .IN4(n28836), .Q(
        n25617) );
  OA22X1 U29333 ( .IN1(n25652), .IN2(n28833), .IN3(n25662), .IN4(n28837), .Q(
        n25616) );
  OA22X1 U29334 ( .IN1(n25663), .IN2(n28834), .IN3(n25619), .IN4(n28829), .Q(
        n25615) );
  NAND4X0 U29335 ( .IN1(n25618), .IN2(n25617), .IN3(n25616), .IN4(n25615), 
        .QN(s9_addr_o[22]) );
  OA22X1 U29336 ( .IN1(n25666), .IN2(n28848), .IN3(n25659), .IN4(n28845), .Q(
        n25623) );
  OA22X1 U29337 ( .IN1(n25660), .IN2(n28843), .IN3(n25665), .IN4(n28852), .Q(
        n25622) );
  OA22X1 U29338 ( .IN1(n25641), .IN2(n28850), .IN3(n25662), .IN4(n28846), .Q(
        n25621) );
  OA22X1 U29339 ( .IN1(n25653), .IN2(n28849), .IN3(n25619), .IN4(n28851), .Q(
        n25620) );
  NAND4X0 U29340 ( .IN1(n25623), .IN2(n25622), .IN3(n25621), .IN4(n25620), 
        .QN(s9_addr_o[23]) );
  OA22X1 U29341 ( .IN1(n28859), .IN2(n25663), .IN3(n28857), .IN4(n25661), .Q(
        n25627) );
  OA22X1 U29342 ( .IN1(n28858), .IN2(n25654), .IN3(n28864), .IN4(n25640), .Q(
        n25626) );
  OA22X1 U29343 ( .IN1(n28860), .IN2(n25664), .IN3(n28861), .IN4(n25665), .Q(
        n25625) );
  OA22X1 U29344 ( .IN1(n28865), .IN2(n25662), .IN3(n28863), .IN4(n25652), .Q(
        n25624) );
  NAND4X0 U29345 ( .IN1(n25627), .IN2(n25626), .IN3(n25625), .IN4(n25624), 
        .QN(s9_addr_o[24]) );
  OA22X1 U29346 ( .IN1(n28871), .IN2(n25650), .IN3(n28876), .IN4(n25663), .Q(
        n25631) );
  OA22X1 U29347 ( .IN1(n28875), .IN2(n25664), .IN3(n28870), .IN4(n25652), .Q(
        n25630) );
  OA22X1 U29348 ( .IN1(n28873), .IN2(n25660), .IN3(n28877), .IN4(n25640), .Q(
        n25629) );
  OA22X1 U29349 ( .IN1(n28874), .IN2(n25641), .IN3(n28872), .IN4(n25665), .Q(
        n25628) );
  NAND4X0 U29350 ( .IN1(n25631), .IN2(n25630), .IN3(n25629), .IN4(n25628), 
        .QN(s9_addr_o[25]) );
  OA22X1 U29351 ( .IN1(n28885), .IN2(n25654), .IN3(n28883), .IN4(n25650), .Q(
        n25635) );
  OA22X1 U29352 ( .IN1(n28889), .IN2(n25664), .IN3(n28884), .IN4(n25652), .Q(
        n25634) );
  OA22X1 U29353 ( .IN1(n28882), .IN2(n25641), .IN3(n28886), .IN4(n25651), .Q(
        n25633) );
  OA22X1 U29354 ( .IN1(n28887), .IN2(n25640), .IN3(n28888), .IN4(n25663), .Q(
        n25632) );
  NAND4X0 U29355 ( .IN1(n25635), .IN2(n25634), .IN3(n25633), .IN4(n25632), 
        .QN(s9_addr_o[26]) );
  OA22X1 U29356 ( .IN1(n28897), .IN2(n25662), .IN3(n28895), .IN4(n25640), .Q(
        n25639) );
  OA22X1 U29357 ( .IN1(n28898), .IN2(n25664), .IN3(n28901), .IN4(n25661), .Q(
        n25638) );
  OA22X1 U29358 ( .IN1(n28896), .IN2(n25653), .IN3(n28894), .IN4(n25652), .Q(
        n25637) );
  OA22X1 U29359 ( .IN1(n28899), .IN2(n25660), .IN3(n28900), .IN4(n25665), .Q(
        n25636) );
  NAND4X0 U29360 ( .IN1(n25639), .IN2(n25638), .IN3(n25637), .IN4(n25636), 
        .QN(s9_addr_o[27]) );
  OA22X1 U29361 ( .IN1(n28911), .IN2(n25640), .IN3(n28912), .IN4(n25652), .Q(
        n25645) );
  OA22X1 U29362 ( .IN1(n28909), .IN2(n25654), .IN3(n28908), .IN4(n25641), .Q(
        n25644) );
  OA22X1 U29363 ( .IN1(n28913), .IN2(n25664), .IN3(n28910), .IN4(n25663), .Q(
        n25643) );
  OA22X1 U29364 ( .IN1(n28907), .IN2(n25650), .IN3(n28906), .IN4(n25651), .Q(
        n25642) );
  NAND4X0 U29365 ( .IN1(n25645), .IN2(n25644), .IN3(n25643), .IN4(n25642), 
        .QN(s9_addr_o[28]) );
  OA22X1 U29366 ( .IN1(n28922), .IN2(n25662), .IN3(n28924), .IN4(n25659), .Q(
        n25649) );
  OA22X1 U29367 ( .IN1(n28926), .IN2(n25660), .IN3(n28925), .IN4(n25652), .Q(
        n25648) );
  OA22X1 U29368 ( .IN1(n28920), .IN2(n25663), .IN3(n28923), .IN4(n25651), .Q(
        n25647) );
  OA22X1 U29369 ( .IN1(n28921), .IN2(n25664), .IN3(n28919), .IN4(n25661), .Q(
        n25646) );
  NAND4X0 U29370 ( .IN1(n25649), .IN2(n25648), .IN3(n25647), .IN4(n25646), 
        .QN(s9_addr_o[29]) );
  OA22X1 U29371 ( .IN1(n28937), .IN2(n25650), .IN3(n28940), .IN4(n25661), .Q(
        n25658) );
  OA22X1 U29372 ( .IN1(n28933), .IN2(n25664), .IN3(n28939), .IN4(n25651), .Q(
        n25657) );
  OA22X1 U29373 ( .IN1(n28936), .IN2(n25653), .IN3(n28931), .IN4(n25652), .Q(
        n25656) );
  OA22X1 U29374 ( .IN1(n28932), .IN2(n25654), .IN3(n28935), .IN4(n25659), .Q(
        n25655) );
  NAND4X0 U29375 ( .IN1(n25658), .IN2(n25657), .IN3(n25656), .IN4(n25655), 
        .QN(s9_addr_o[30]) );
  OA22X1 U29376 ( .IN1(n28948), .IN2(n25660), .IN3(n28952), .IN4(n25659), .Q(
        n25670) );
  OA22X1 U29377 ( .IN1(n28956), .IN2(n25662), .IN3(n28958), .IN4(n25661), .Q(
        n25669) );
  OA22X1 U29378 ( .IN1(n28960), .IN2(n25664), .IN3(n28954), .IN4(n25663), .Q(
        n25668) );
  OA22X1 U29379 ( .IN1(n28950), .IN2(n25666), .IN3(n28946), .IN4(n25665), .Q(
        n25667) );
  NAND4X0 U29380 ( .IN1(n25670), .IN2(n25669), .IN3(n25668), .IN4(n25667), 
        .QN(s9_addr_o[31]) );
  OA22X1 U29381 ( .IN1(n29235), .IN2(n25672), .IN3(n29292), .IN4(n25671), .Q(
        n25682) );
  OA22X1 U29382 ( .IN1(n29368), .IN2(n25674), .IN3(n29311), .IN4(n25673), .Q(
        n25681) );
  OA22X1 U29383 ( .IN1(n29273), .IN2(n25676), .IN3(n29349), .IN4(n25675), .Q(
        n25680) );
  OA22X1 U29384 ( .IN1(n29254), .IN2(n25678), .IN3(n29330), .IN4(n25677), .Q(
        n25679) );
  NAND4X0 U29385 ( .IN1(n25682), .IN2(n25681), .IN3(n25680), .IN4(n25679), 
        .QN(s8_stb_o) );
  INVX0 U29386 ( .INP(n29119), .ZN(n25932) );
  OA22X1 U29387 ( .IN1(n25932), .IN2(n28126), .IN3(n25969), .IN4(n28122), .Q(
        n25686) );
  INVX0 U29388 ( .INP(n29112), .ZN(n25956) );
  INVX0 U29389 ( .INP(n29111), .ZN(n25964) );
  OA22X1 U29390 ( .IN1(n25956), .IN2(n28123), .IN3(n25964), .IN4(n28121), .Q(
        n25685) );
  INVX0 U29391 ( .INP(n29120), .ZN(n25965) );
  OA22X1 U29392 ( .IN1(n25965), .IN2(n28124), .IN3(n25967), .IN4(n28125), .Q(
        n25684) );
  INVX0 U29393 ( .INP(n29117), .ZN(n25968) );
  INVX0 U29394 ( .INP(n29109), .ZN(n25966) );
  OA22X1 U29395 ( .IN1(n25968), .IN2(n28128), .IN3(n25966), .IN4(n28127), .Q(
        n25683) );
  NAND4X0 U29396 ( .IN1(n25686), .IN2(n25685), .IN3(n25684), .IN4(n25683), 
        .QN(s8_we_o) );
  INVX0 U29397 ( .INP(n29112), .ZN(n25970) );
  INVX0 U29398 ( .INP(n29119), .ZN(n25963) );
  OA22X1 U29399 ( .IN1(n25970), .IN2(n28133), .IN3(n25963), .IN4(n28139), .Q(
        n25690) );
  INVX0 U29400 ( .INP(n29117), .ZN(n25955) );
  OA22X1 U29401 ( .IN1(n25965), .IN2(n28134), .IN3(n25955), .IN4(n28140), .Q(
        n25689) );
  INVX0 U29402 ( .INP(n25969), .ZN(n29110) );
  INVX0 U29403 ( .INP(n29110), .ZN(n25915) );
  INVX0 U29404 ( .INP(n29111), .ZN(n25957) );
  OA22X1 U29405 ( .IN1(n25915), .IN2(n28138), .IN3(n25957), .IN4(n28135), .Q(
        n25688) );
  INVX0 U29406 ( .INP(n25967), .ZN(n29118) );
  INVX0 U29407 ( .INP(n29118), .ZN(n25950) );
  INVX0 U29408 ( .INP(n29109), .ZN(n25958) );
  OA22X1 U29409 ( .IN1(n25950), .IN2(n28136), .IN3(n25958), .IN4(n28137), .Q(
        n25687) );
  NAND4X0 U29410 ( .IN1(n25690), .IN2(n25689), .IN3(n25688), .IN4(n25687), 
        .QN(s8_data_o[0]) );
  OA22X1 U29411 ( .IN1(n25956), .IN2(n28148), .IN3(n25969), .IN4(n28149), .Q(
        n25694) );
  OA22X1 U29412 ( .IN1(n25965), .IN2(n28150), .IN3(n25967), .IN4(n28152), .Q(
        n25693) );
  OA22X1 U29413 ( .IN1(n25955), .IN2(n28146), .IN3(n25963), .IN4(n28145), .Q(
        n25692) );
  OA22X1 U29414 ( .IN1(n25958), .IN2(n28151), .IN3(n25957), .IN4(n28147), .Q(
        n25691) );
  NAND4X0 U29415 ( .IN1(n25694), .IN2(n25693), .IN3(n25692), .IN4(n25691), 
        .QN(s8_data_o[1]) );
  OA22X1 U29416 ( .IN1(n25968), .IN2(n28164), .IN3(n25963), .IN4(n28159), .Q(
        n25698) );
  OA22X1 U29417 ( .IN1(n25915), .IN2(n28158), .IN3(n25967), .IN4(n28162), .Q(
        n25697) );
  OA22X1 U29418 ( .IN1(n25966), .IN2(n28157), .IN3(n25957), .IN4(n28161), .Q(
        n25696) );
  OA22X1 U29419 ( .IN1(n25965), .IN2(n28160), .IN3(n25956), .IN4(n28163), .Q(
        n25695) );
  NAND4X0 U29420 ( .IN1(n25698), .IN2(n25697), .IN3(n25696), .IN4(n25695), 
        .QN(s8_data_o[2]) );
  OA22X1 U29421 ( .IN1(n25965), .IN2(n28172), .IN3(n25957), .IN4(n28173), .Q(
        n25702) );
  OA22X1 U29422 ( .IN1(n25956), .IN2(n28176), .IN3(n25966), .IN4(n28169), .Q(
        n25701) );
  OA22X1 U29423 ( .IN1(n25955), .IN2(n28174), .IN3(n25963), .IN4(n28170), .Q(
        n25700) );
  OA22X1 U29424 ( .IN1(n25915), .IN2(n28171), .IN3(n25967), .IN4(n28175), .Q(
        n25699) );
  NAND4X0 U29425 ( .IN1(n25702), .IN2(n25701), .IN3(n25700), .IN4(n25699), 
        .QN(s8_data_o[3]) );
  INVX0 U29426 ( .INP(n29120), .ZN(n25945) );
  OA22X1 U29427 ( .IN1(n25945), .IN2(n28182), .IN3(n25957), .IN4(n28181), .Q(
        n25706) );
  OA22X1 U29428 ( .IN1(n25932), .IN2(n28188), .IN3(n25967), .IN4(n28183), .Q(
        n25705) );
  OA22X1 U29429 ( .IN1(n25970), .IN2(n28186), .IN3(n25969), .IN4(n28185), .Q(
        n25704) );
  OA22X1 U29430 ( .IN1(n25968), .IN2(n28184), .IN3(n25966), .IN4(n28187), .Q(
        n25703) );
  NAND4X0 U29431 ( .IN1(n25706), .IN2(n25705), .IN3(n25704), .IN4(n25703), 
        .QN(s8_data_o[4]) );
  OA22X1 U29432 ( .IN1(n25968), .IN2(n28200), .IN3(n25967), .IN4(n28197), .Q(
        n25710) );
  OA22X1 U29433 ( .IN1(n25965), .IN2(n28196), .IN3(n25966), .IN4(n28195), .Q(
        n25709) );
  OA22X1 U29434 ( .IN1(n25970), .IN2(n28194), .IN3(n25969), .IN4(n28198), .Q(
        n25708) );
  OA22X1 U29435 ( .IN1(n25932), .IN2(n28193), .IN3(n25957), .IN4(n28199), .Q(
        n25707) );
  NAND4X0 U29436 ( .IN1(n25710), .IN2(n25709), .IN3(n25708), .IN4(n25707), 
        .QN(s8_data_o[5]) );
  OA22X1 U29437 ( .IN1(n25958), .IN2(n28210), .IN3(n25957), .IN4(n28209), .Q(
        n25714) );
  OA22X1 U29438 ( .IN1(n25965), .IN2(n28208), .IN3(n25967), .IN4(n28205), .Q(
        n25713) );
  OA22X1 U29439 ( .IN1(n25955), .IN2(n28207), .IN3(n25956), .IN4(n28206), .Q(
        n25712) );
  OA22X1 U29440 ( .IN1(n25963), .IN2(n28212), .IN3(n25969), .IN4(n28211), .Q(
        n25711) );
  NAND4X0 U29441 ( .IN1(n25714), .IN2(n25713), .IN3(n25712), .IN4(n25711), 
        .QN(s8_data_o[6]) );
  OA22X1 U29442 ( .IN1(n25963), .IN2(n28218), .IN3(n25967), .IN4(n28223), .Q(
        n25718) );
  OA22X1 U29443 ( .IN1(n25915), .IN2(n28217), .IN3(n25966), .IN4(n28222), .Q(
        n25717) );
  OA22X1 U29444 ( .IN1(n25965), .IN2(n28220), .IN3(n25956), .IN4(n28224), .Q(
        n25716) );
  OA22X1 U29445 ( .IN1(n25955), .IN2(n28219), .IN3(n25964), .IN4(n28221), .Q(
        n25715) );
  NAND4X0 U29446 ( .IN1(n25718), .IN2(n25717), .IN3(n25716), .IN4(n25715), 
        .QN(s8_data_o[7]) );
  OA22X1 U29447 ( .IN1(n25956), .IN2(n28231), .IN3(n25967), .IN4(n28229), .Q(
        n25722) );
  OA22X1 U29448 ( .IN1(n25932), .IN2(n28234), .IN3(n25969), .IN4(n28236), .Q(
        n25721) );
  OA22X1 U29449 ( .IN1(n25945), .IN2(n28230), .IN3(n25966), .IN4(n28233), .Q(
        n25720) );
  OA22X1 U29450 ( .IN1(n25968), .IN2(n28232), .IN3(n25964), .IN4(n28235), .Q(
        n25719) );
  NAND4X0 U29451 ( .IN1(n25722), .IN2(n25721), .IN3(n25720), .IN4(n25719), 
        .QN(s8_data_o[8]) );
  OA22X1 U29452 ( .IN1(n25963), .IN2(n28248), .IN3(n25969), .IN4(n28241), .Q(
        n25726) );
  OA22X1 U29453 ( .IN1(n25956), .IN2(n28246), .IN3(n25966), .IN4(n28243), .Q(
        n25725) );
  OA22X1 U29454 ( .IN1(n25945), .IN2(n28242), .IN3(n25955), .IN4(n28244), .Q(
        n25724) );
  OA22X1 U29455 ( .IN1(n25950), .IN2(n28245), .IN3(n25964), .IN4(n28247), .Q(
        n25723) );
  NAND4X0 U29456 ( .IN1(n25726), .IN2(n25725), .IN3(n25724), .IN4(n25723), 
        .QN(s8_data_o[9]) );
  OA22X1 U29457 ( .IN1(n25970), .IN2(n28260), .IN3(n25969), .IN4(n28254), .Q(
        n25730) );
  OA22X1 U29458 ( .IN1(n25965), .IN2(n28258), .IN3(n25964), .IN4(n28259), .Q(
        n25729) );
  OA22X1 U29459 ( .IN1(n25932), .IN2(n28256), .IN3(n25967), .IN4(n28255), .Q(
        n25728) );
  OA22X1 U29460 ( .IN1(n25955), .IN2(n28257), .IN3(n25966), .IN4(n28253), .Q(
        n25727) );
  NAND4X0 U29461 ( .IN1(n25730), .IN2(n25729), .IN3(n25728), .IN4(n25727), 
        .QN(s8_data_o[10]) );
  OA22X1 U29462 ( .IN1(n25955), .IN2(n28272), .IN3(n25969), .IN4(n28268), .Q(
        n25734) );
  OA22X1 U29463 ( .IN1(n25945), .IN2(n28266), .IN3(n25966), .IN4(n28267), .Q(
        n25733) );
  OA22X1 U29464 ( .IN1(n25950), .IN2(n28270), .IN3(n25964), .IN4(n28269), .Q(
        n25732) );
  OA22X1 U29465 ( .IN1(n25956), .IN2(n28265), .IN3(n25932), .IN4(n28271), .Q(
        n25731) );
  NAND4X0 U29466 ( .IN1(n25734), .IN2(n25733), .IN3(n25732), .IN4(n25731), 
        .QN(s8_data_o[11]) );
  OA22X1 U29467 ( .IN1(n25950), .IN2(n28281), .IN3(n25964), .IN4(n28277), .Q(
        n25738) );
  OA22X1 U29468 ( .IN1(n25968), .IN2(n28278), .IN3(n25969), .IN4(n28283), .Q(
        n25737) );
  OA22X1 U29469 ( .IN1(n25956), .IN2(n28280), .IN3(n25966), .IN4(n28279), .Q(
        n25736) );
  OA22X1 U29470 ( .IN1(n25965), .IN2(n28284), .IN3(n25963), .IN4(n28282), .Q(
        n25735) );
  NAND4X0 U29471 ( .IN1(n25738), .IN2(n25737), .IN3(n25736), .IN4(n25735), 
        .QN(s8_data_o[12]) );
  OA22X1 U29472 ( .IN1(n25965), .IN2(n28290), .IN3(n25955), .IN4(n28294), .Q(
        n25742) );
  OA22X1 U29473 ( .IN1(n25956), .IN2(n28296), .IN3(n25915), .IN4(n28289), .Q(
        n25741) );
  OA22X1 U29474 ( .IN1(n25950), .IN2(n28293), .IN3(n25964), .IN4(n28295), .Q(
        n25740) );
  OA22X1 U29475 ( .IN1(n25932), .IN2(n28292), .IN3(n25958), .IN4(n28291), .Q(
        n25739) );
  NAND4X0 U29476 ( .IN1(n25742), .IN2(n25741), .IN3(n25740), .IN4(n25739), 
        .QN(s8_data_o[13]) );
  OA22X1 U29477 ( .IN1(n25945), .IN2(n28306), .IN3(n25956), .IN4(n28308), .Q(
        n25746) );
  OA22X1 U29478 ( .IN1(n25968), .IN2(n28304), .IN3(n25950), .IN4(n28302), .Q(
        n25745) );
  OA22X1 U29479 ( .IN1(n25915), .IN2(n28307), .IN3(n25964), .IN4(n28303), .Q(
        n25744) );
  OA22X1 U29480 ( .IN1(n25932), .IN2(n28305), .IN3(n25958), .IN4(n28301), .Q(
        n25743) );
  NAND4X0 U29481 ( .IN1(n25746), .IN2(n25745), .IN3(n25744), .IN4(n25743), 
        .QN(s8_data_o[14]) );
  OA22X1 U29482 ( .IN1(n25965), .IN2(n28316), .IN3(n25963), .IN4(n28313), .Q(
        n25750) );
  OA22X1 U29483 ( .IN1(n25955), .IN2(n28315), .IN3(n25958), .IN4(n28317), .Q(
        n25749) );
  OA22X1 U29484 ( .IN1(n25956), .IN2(n28314), .IN3(n25915), .IN4(n28320), .Q(
        n25748) );
  OA22X1 U29485 ( .IN1(n25950), .IN2(n28318), .IN3(n25964), .IN4(n28319), .Q(
        n25747) );
  NAND4X0 U29486 ( .IN1(n25750), .IN2(n25749), .IN3(n25748), .IN4(n25747), 
        .QN(s8_data_o[15]) );
  OA22X1 U29487 ( .IN1(n25963), .IN2(n28326), .IN3(n25950), .IN4(n28325), .Q(
        n25754) );
  OA22X1 U29488 ( .IN1(n25970), .IN2(n28331), .IN3(n25964), .IN4(n28327), .Q(
        n25753) );
  OA22X1 U29489 ( .IN1(n25945), .IN2(n28330), .IN3(n25955), .IN4(n28332), .Q(
        n25752) );
  OA22X1 U29490 ( .IN1(n25915), .IN2(n28329), .IN3(n25958), .IN4(n28328), .Q(
        n25751) );
  NAND4X0 U29491 ( .IN1(n25754), .IN2(n25753), .IN3(n25752), .IN4(n25751), 
        .QN(s8_data_o[16]) );
  OA22X1 U29492 ( .IN1(n25955), .IN2(n28344), .IN3(n25915), .IN4(n28337), .Q(
        n25758) );
  OA22X1 U29493 ( .IN1(n25963), .IN2(n28338), .IN3(n25964), .IN4(n28341), .Q(
        n25757) );
  OA22X1 U29494 ( .IN1(n25965), .IN2(n28340), .IN3(n25950), .IN4(n28339), .Q(
        n25756) );
  OA22X1 U29495 ( .IN1(n25956), .IN2(n28342), .IN3(n25958), .IN4(n28343), .Q(
        n25755) );
  NAND4X0 U29496 ( .IN1(n25758), .IN2(n25757), .IN3(n25756), .IN4(n25755), 
        .QN(s8_data_o[17]) );
  OA22X1 U29497 ( .IN1(n25970), .IN2(n28350), .IN3(n25932), .IN4(n28355), .Q(
        n25762) );
  OA22X1 U29498 ( .IN1(n25955), .IN2(n28356), .IN3(n25958), .IN4(n28351), .Q(
        n25761) );
  OA22X1 U29499 ( .IN1(n25915), .IN2(n28354), .IN3(n25964), .IN4(n28353), .Q(
        n25760) );
  OA22X1 U29500 ( .IN1(n25965), .IN2(n28352), .IN3(n25950), .IN4(n28349), .Q(
        n25759) );
  NAND4X0 U29501 ( .IN1(n25762), .IN2(n25761), .IN3(n25760), .IN4(n25759), 
        .QN(s8_data_o[18]) );
  OA22X1 U29502 ( .IN1(n25967), .IN2(n28361), .IN3(n25958), .IN4(n28368), .Q(
        n25766) );
  OA22X1 U29503 ( .IN1(n25968), .IN2(n28364), .IN3(n25915), .IN4(n28365), .Q(
        n25765) );
  OA22X1 U29504 ( .IN1(n25945), .IN2(n28366), .IN3(n25964), .IN4(n28367), .Q(
        n25764) );
  OA22X1 U29505 ( .IN1(n25970), .IN2(n28362), .IN3(n25963), .IN4(n28363), .Q(
        n25763) );
  NAND4X0 U29506 ( .IN1(n25766), .IN2(n25765), .IN3(n25764), .IN4(n25763), 
        .QN(s8_data_o[19]) );
  OA22X1 U29507 ( .IN1(n25967), .IN2(n28380), .IN3(n25964), .IN4(n28375), .Q(
        n25770) );
  OA22X1 U29508 ( .IN1(n25969), .IN2(n28376), .IN3(n25958), .IN4(n28379), .Q(
        n25769) );
  OA22X1 U29509 ( .IN1(n25965), .IN2(n28378), .IN3(n25963), .IN4(n28373), .Q(
        n25768) );
  OA22X1 U29510 ( .IN1(n25955), .IN2(n28377), .IN3(n25956), .IN4(n28374), .Q(
        n25767) );
  NAND4X0 U29511 ( .IN1(n25770), .IN2(n25769), .IN3(n25768), .IN4(n25767), 
        .QN(s8_data_o[20]) );
  OA22X1 U29512 ( .IN1(n25956), .IN2(n28390), .IN3(n25958), .IN4(n28389), .Q(
        n25774) );
  OA22X1 U29513 ( .IN1(n25932), .IN2(n28388), .IN3(n25950), .IN4(n28385), .Q(
        n25773) );
  OA22X1 U29514 ( .IN1(n25945), .IN2(n28392), .IN3(n25964), .IN4(n28391), .Q(
        n25772) );
  OA22X1 U29515 ( .IN1(n25968), .IN2(n28386), .IN3(n25915), .IN4(n28387), .Q(
        n25771) );
  NAND4X0 U29516 ( .IN1(n25774), .IN2(n25773), .IN3(n25772), .IN4(n25771), 
        .QN(s8_data_o[21]) );
  OA22X1 U29517 ( .IN1(n25965), .IN2(n28400), .IN3(n25964), .IN4(n28397), .Q(
        n25778) );
  OA22X1 U29518 ( .IN1(n25970), .IN2(n28404), .IN3(n25963), .IN4(n28403), .Q(
        n25777) );
  OA22X1 U29519 ( .IN1(n25969), .IN2(n28398), .IN3(n25958), .IN4(n28401), .Q(
        n25776) );
  OA22X1 U29520 ( .IN1(n25968), .IN2(n28402), .IN3(n25950), .IN4(n28399), .Q(
        n25775) );
  NAND4X0 U29521 ( .IN1(n25778), .IN2(n25777), .IN3(n25776), .IN4(n25775), 
        .QN(s8_data_o[22]) );
  OA22X1 U29522 ( .IN1(n25945), .IN2(n28416), .IN3(n25932), .IN4(n28413), .Q(
        n25782) );
  OA22X1 U29523 ( .IN1(n25915), .IN2(n28410), .IN3(n25958), .IN4(n28409), .Q(
        n25781) );
  OA22X1 U29524 ( .IN1(n25970), .IN2(n28414), .IN3(n25957), .IN4(n28411), .Q(
        n25780) );
  OA22X1 U29525 ( .IN1(n25955), .IN2(n28415), .IN3(n25950), .IN4(n28412), .Q(
        n25779) );
  NAND4X0 U29526 ( .IN1(n25782), .IN2(n25781), .IN3(n25780), .IN4(n25779), 
        .QN(s8_data_o[23]) );
  OA22X1 U29527 ( .IN1(n25965), .IN2(n28426), .IN3(n25963), .IN4(n28421), .Q(
        n25786) );
  OA22X1 U29528 ( .IN1(n25967), .IN2(n28428), .IN3(n25958), .IN4(n28427), .Q(
        n25785) );
  OA22X1 U29529 ( .IN1(n25956), .IN2(n28422), .IN3(n25915), .IN4(n28425), .Q(
        n25784) );
  OA22X1 U29530 ( .IN1(n25955), .IN2(n28424), .IN3(n25964), .IN4(n28423), .Q(
        n25783) );
  NAND4X0 U29531 ( .IN1(n25786), .IN2(n25785), .IN3(n25784), .IN4(n25783), 
        .QN(s8_data_o[24]) );
  OA22X1 U29532 ( .IN1(n25932), .IN2(n28439), .IN3(n25957), .IN4(n28435), .Q(
        n25790) );
  OA22X1 U29533 ( .IN1(n25969), .IN2(n28433), .IN3(n25950), .IN4(n28437), .Q(
        n25789) );
  OA22X1 U29534 ( .IN1(n25945), .IN2(n28438), .IN3(n25955), .IN4(n28440), .Q(
        n25788) );
  OA22X1 U29535 ( .IN1(n25956), .IN2(n28434), .IN3(n25958), .IN4(n28436), .Q(
        n25787) );
  NAND4X0 U29536 ( .IN1(n25790), .IN2(n25789), .IN3(n25788), .IN4(n25787), 
        .QN(s8_data_o[25]) );
  OA22X1 U29537 ( .IN1(n25968), .IN2(n28451), .IN3(n25915), .IN4(n28449), .Q(
        n25794) );
  OA22X1 U29538 ( .IN1(n25932), .IN2(n28446), .IN3(n25950), .IN4(n28448), .Q(
        n25793) );
  OA22X1 U29539 ( .IN1(n25966), .IN2(n28447), .IN3(n25957), .IN4(n28445), .Q(
        n25792) );
  OA22X1 U29540 ( .IN1(n25945), .IN2(n28452), .IN3(n25956), .IN4(n28450), .Q(
        n25791) );
  NAND4X0 U29541 ( .IN1(n25794), .IN2(n25793), .IN3(n25792), .IN4(n25791), 
        .QN(s8_data_o[26]) );
  OA22X1 U29542 ( .IN1(n25945), .IN2(n28462), .IN3(n25955), .IN4(n28461), .Q(
        n25798) );
  OA22X1 U29543 ( .IN1(n25970), .IN2(n28464), .IN3(n25958), .IN4(n28460), .Q(
        n25797) );
  OA22X1 U29544 ( .IN1(n25915), .IN2(n28457), .IN3(n25964), .IN4(n28459), .Q(
        n25796) );
  OA22X1 U29545 ( .IN1(n25932), .IN2(n28458), .IN3(n25950), .IN4(n28463), .Q(
        n25795) );
  NAND4X0 U29546 ( .IN1(n25798), .IN2(n25797), .IN3(n25796), .IN4(n25795), 
        .QN(s8_data_o[27]) );
  OA22X1 U29547 ( .IN1(n25965), .IN2(n28474), .IN3(n25950), .IN4(n28475), .Q(
        n25802) );
  OA22X1 U29548 ( .IN1(n25969), .IN2(n28471), .IN3(n25964), .IN4(n28473), .Q(
        n25801) );
  OA22X1 U29549 ( .IN1(n25968), .IN2(n28476), .IN3(n25958), .IN4(n28469), .Q(
        n25800) );
  OA22X1 U29550 ( .IN1(n25956), .IN2(n28472), .IN3(n25932), .IN4(n28470), .Q(
        n25799) );
  NAND4X0 U29551 ( .IN1(n25802), .IN2(n25801), .IN3(n25800), .IN4(n25799), 
        .QN(s8_data_o[28]) );
  OA22X1 U29552 ( .IN1(n25955), .IN2(n28482), .IN3(n25956), .IN4(n28488), .Q(
        n25806) );
  OA22X1 U29553 ( .IN1(n25967), .IN2(n28483), .IN3(n25958), .IN4(n28485), .Q(
        n25805) );
  OA22X1 U29554 ( .IN1(n25932), .IN2(n28486), .IN3(n25915), .IN4(n28487), .Q(
        n25804) );
  OA22X1 U29555 ( .IN1(n25945), .IN2(n28484), .IN3(n25957), .IN4(n28481), .Q(
        n25803) );
  NAND4X0 U29556 ( .IN1(n25806), .IN2(n25805), .IN3(n25804), .IN4(n25803), 
        .QN(s8_data_o[29]) );
  OA22X1 U29557 ( .IN1(n25965), .IN2(n28494), .IN3(n25963), .IN4(n28496), .Q(
        n25810) );
  OA22X1 U29558 ( .IN1(n25968), .IN2(n28498), .IN3(n25964), .IN4(n28499), .Q(
        n25809) );
  OA22X1 U29559 ( .IN1(n25967), .IN2(n28495), .IN3(n25958), .IN4(n28500), .Q(
        n25808) );
  OA22X1 U29560 ( .IN1(n25970), .IN2(n28497), .IN3(n25915), .IN4(n28493), .Q(
        n25807) );
  NAND4X0 U29561 ( .IN1(n25810), .IN2(n25809), .IN3(n25808), .IN4(n25807), 
        .QN(s8_data_o[30]) );
  OA22X1 U29562 ( .IN1(n25945), .IN2(n28510), .IN3(n25956), .IN4(n28506), .Q(
        n25814) );
  OA22X1 U29563 ( .IN1(n25932), .IN2(n28505), .IN3(n25950), .IN4(n28508), .Q(
        n25813) );
  OA22X1 U29564 ( .IN1(n25969), .IN2(n28512), .IN3(n25957), .IN4(n28507), .Q(
        n25812) );
  OA22X1 U29565 ( .IN1(n25968), .IN2(n28509), .IN3(n25958), .IN4(n28511), .Q(
        n25811) );
  NAND4X0 U29566 ( .IN1(n25814), .IN2(n25813), .IN3(n25812), .IN4(n25811), 
        .QN(s8_data_o[31]) );
  OA22X1 U29567 ( .IN1(n25945), .IN2(n28518), .IN3(n25966), .IN4(n28521), .Q(
        n25818) );
  OA22X1 U29568 ( .IN1(n25970), .IN2(n28522), .IN3(n25957), .IN4(n28519), .Q(
        n25817) );
  OA22X1 U29569 ( .IN1(n25955), .IN2(n28517), .IN3(n25915), .IN4(n28523), .Q(
        n25816) );
  OA22X1 U29570 ( .IN1(n25932), .IN2(n28524), .IN3(n25950), .IN4(n28520), .Q(
        n25815) );
  NAND4X0 U29571 ( .IN1(n25818), .IN2(n25817), .IN3(n25816), .IN4(n25815), 
        .QN(s8_sel_o[0]) );
  OA22X1 U29572 ( .IN1(n25945), .IN2(n28534), .IN3(n25950), .IN4(n28533), .Q(
        n25822) );
  OA22X1 U29573 ( .IN1(n25932), .IN2(n28536), .IN3(n25958), .IN4(n28531), .Q(
        n25821) );
  OA22X1 U29574 ( .IN1(n25970), .IN2(n28530), .IN3(n25964), .IN4(n28529), .Q(
        n25820) );
  OA22X1 U29575 ( .IN1(n25968), .IN2(n28532), .IN3(n25915), .IN4(n28535), .Q(
        n25819) );
  NAND4X0 U29576 ( .IN1(n25822), .IN2(n25821), .IN3(n25820), .IN4(n25819), 
        .QN(s8_sel_o[1]) );
  OA22X1 U29577 ( .IN1(n25915), .IN2(n28547), .IN3(n25966), .IN4(n28545), .Q(
        n25826) );
  OA22X1 U29578 ( .IN1(n25968), .IN2(n28546), .IN3(n25963), .IN4(n28548), .Q(
        n25825) );
  OA22X1 U29579 ( .IN1(n25945), .IN2(n28544), .IN3(n25950), .IN4(n28542), .Q(
        n25824) );
  OA22X1 U29580 ( .IN1(n25970), .IN2(n28543), .IN3(n25964), .IN4(n28541), .Q(
        n25823) );
  NAND4X0 U29581 ( .IN1(n25826), .IN2(n25825), .IN3(n25824), .IN4(n25823), 
        .QN(s8_sel_o[2]) );
  OA22X1 U29582 ( .IN1(n25970), .IN2(n28553), .IN3(n25966), .IN4(n28559), .Q(
        n25830) );
  OA22X1 U29583 ( .IN1(n25945), .IN2(n28558), .IN3(n25955), .IN4(n28554), .Q(
        n25829) );
  OA22X1 U29584 ( .IN1(n25932), .IN2(n28557), .IN3(n25950), .IN4(n28560), .Q(
        n25828) );
  OA22X1 U29585 ( .IN1(n25969), .IN2(n28556), .IN3(n25957), .IN4(n28555), .Q(
        n25827) );
  NAND4X0 U29586 ( .IN1(n25830), .IN2(n25829), .IN3(n25828), .IN4(n25827), 
        .QN(s8_sel_o[3]) );
  OA22X1 U29587 ( .IN1(n25932), .IN2(n28566), .IN3(n25967), .IN4(n28567), .Q(
        n25834) );
  OA22X1 U29588 ( .IN1(n25945), .IN2(n28572), .IN3(n25958), .IN4(n28565), .Q(
        n25833) );
  OA22X1 U29589 ( .IN1(n25970), .IN2(n28571), .IN3(n25915), .IN4(n28568), .Q(
        n25832) );
  OA22X1 U29590 ( .IN1(n25968), .IN2(n28570), .IN3(n25964), .IN4(n28569), .Q(
        n25831) );
  NAND4X0 U29591 ( .IN1(n25834), .IN2(n25833), .IN3(n25832), .IN4(n25831), 
        .QN(s8_addr_o[0]) );
  OA22X1 U29592 ( .IN1(n25968), .IN2(n28578), .IN3(n25958), .IN4(n28577), .Q(
        n25838) );
  OA22X1 U29593 ( .IN1(n25932), .IN2(n28581), .IN3(n25915), .IN4(n28579), .Q(
        n25837) );
  OA22X1 U29594 ( .IN1(n25945), .IN2(n28580), .IN3(n25967), .IN4(n28584), .Q(
        n25836) );
  OA22X1 U29595 ( .IN1(n25970), .IN2(n28582), .IN3(n25957), .IN4(n28583), .Q(
        n25835) );
  NAND4X0 U29596 ( .IN1(n25838), .IN2(n25837), .IN3(n25836), .IN4(n25835), 
        .QN(s8_addr_o[1]) );
  OA22X1 U29597 ( .IN1(n28592), .IN2(n25932), .IN3(n28595), .IN4(n25966), .Q(
        n25842) );
  OA22X1 U29598 ( .IN1(n28594), .IN2(n25970), .IN3(n28590), .IN4(n25969), .Q(
        n25841) );
  OA22X1 U29599 ( .IN1(n28596), .IN2(n25964), .IN3(n28589), .IN4(n25955), .Q(
        n25840) );
  OA22X1 U29600 ( .IN1(n28591), .IN2(n25965), .IN3(n28593), .IN4(n25967), .Q(
        n25839) );
  NAND4X0 U29601 ( .IN1(n25842), .IN2(n25841), .IN3(n25840), .IN4(n25839), 
        .QN(s8_addr_o[2]) );
  OA22X1 U29602 ( .IN1(n28603), .IN2(n25958), .IN3(n28607), .IN4(n25963), .Q(
        n25846) );
  OA22X1 U29603 ( .IN1(n28602), .IN2(n25950), .IN3(n28608), .IN4(n25957), .Q(
        n25845) );
  OA22X1 U29604 ( .IN1(n28604), .IN2(n25956), .IN3(n28605), .IN4(n25955), .Q(
        n25844) );
  OA22X1 U29605 ( .IN1(n28606), .IN2(n25915), .IN3(n28601), .IN4(n25965), .Q(
        n25843) );
  NAND4X0 U29606 ( .IN1(n25846), .IN2(n25845), .IN3(n25844), .IN4(n25843), 
        .QN(s8_addr_o[3]) );
  OA22X1 U29607 ( .IN1(n28616), .IN2(n25955), .IN3(n28619), .IN4(n25964), .Q(
        n25850) );
  OA22X1 U29608 ( .IN1(n28618), .IN2(n25963), .IN3(n28615), .IN4(n25969), .Q(
        n25849) );
  OA22X1 U29609 ( .IN1(n28620), .IN2(n25966), .IN3(n28613), .IN4(n25956), .Q(
        n25848) );
  OA22X1 U29610 ( .IN1(n28614), .IN2(n25950), .IN3(n28617), .IN4(n25965), .Q(
        n25847) );
  NAND4X0 U29611 ( .IN1(n25850), .IN2(n25849), .IN3(n25848), .IN4(n25847), 
        .QN(s8_addr_o[4]) );
  OA22X1 U29612 ( .IN1(n28632), .IN2(n25970), .IN3(n28628), .IN4(n25966), .Q(
        n25854) );
  OA22X1 U29613 ( .IN1(n28626), .IN2(n25932), .IN3(n28629), .IN4(n25965), .Q(
        n25853) );
  OA22X1 U29614 ( .IN1(n28627), .IN2(n25950), .IN3(n28625), .IN4(n25957), .Q(
        n25852) );
  OA22X1 U29615 ( .IN1(n28631), .IN2(n25915), .IN3(n28630), .IN4(n25955), .Q(
        n25851) );
  NAND4X0 U29616 ( .IN1(n25854), .IN2(n25853), .IN3(n25852), .IN4(n25851), 
        .QN(s8_addr_o[5]) );
  OA22X1 U29617 ( .IN1(n25945), .IN2(n28642), .IN3(n25966), .IN4(n28641), .Q(
        n25858) );
  OA22X1 U29618 ( .IN1(n25968), .IN2(n28640), .IN3(n25967), .IN4(n28637), .Q(
        n25857) );
  OA22X1 U29619 ( .IN1(n25970), .IN2(n28644), .IN3(n25915), .IN4(n28638), .Q(
        n25856) );
  OA22X1 U29620 ( .IN1(n25963), .IN2(n28643), .IN3(n25957), .IN4(n28639), .Q(
        n25855) );
  NAND4X0 U29621 ( .IN1(n25858), .IN2(n25857), .IN3(n25856), .IN4(n25855), 
        .QN(s8_addr_o[6]) );
  OA22X1 U29622 ( .IN1(n25945), .IN2(n28654), .IN3(n25915), .IN4(n28650), .Q(
        n25862) );
  OA22X1 U29623 ( .IN1(n25932), .IN2(n28653), .IN3(n25957), .IN4(n28655), .Q(
        n25861) );
  OA22X1 U29624 ( .IN1(n25970), .IN2(n28656), .IN3(n25967), .IN4(n28649), .Q(
        n25860) );
  OA22X1 U29625 ( .IN1(n25968), .IN2(n28652), .IN3(n25958), .IN4(n28651), .Q(
        n25859) );
  NAND4X0 U29626 ( .IN1(n25862), .IN2(n25861), .IN3(n25860), .IN4(n25859), 
        .QN(s8_addr_o[7]) );
  OA22X1 U29627 ( .IN1(n25970), .IN2(n28666), .IN3(n25969), .IN4(n28668), .Q(
        n25866) );
  OA22X1 U29628 ( .IN1(n25968), .IN2(n28663), .IN3(n25963), .IN4(n28665), .Q(
        n25865) );
  OA22X1 U29629 ( .IN1(n25967), .IN2(n28662), .IN3(n25957), .IN4(n28667), .Q(
        n25864) );
  OA22X1 U29630 ( .IN1(n25945), .IN2(n28664), .IN3(n25966), .IN4(n28661), .Q(
        n25863) );
  NAND4X0 U29631 ( .IN1(n25866), .IN2(n25865), .IN3(n25864), .IN4(n25863), 
        .QN(s8_addr_o[8]) );
  OA22X1 U29632 ( .IN1(n25968), .IN2(n28679), .IN3(n25969), .IN4(n28673), .Q(
        n25870) );
  OA22X1 U29633 ( .IN1(n25966), .IN2(n28675), .IN3(n25957), .IN4(n28677), .Q(
        n25869) );
  OA22X1 U29634 ( .IN1(n25970), .IN2(n28674), .IN3(n25967), .IN4(n28678), .Q(
        n25868) );
  OA22X1 U29635 ( .IN1(n25945), .IN2(n28680), .IN3(n25932), .IN4(n28676), .Q(
        n25867) );
  NAND4X0 U29636 ( .IN1(n25870), .IN2(n25869), .IN3(n25868), .IN4(n25867), 
        .QN(s8_addr_o[9]) );
  OA22X1 U29637 ( .IN1(n25970), .IN2(n28688), .IN3(n25966), .IN4(n28690), .Q(
        n25874) );
  OA22X1 U29638 ( .IN1(n25968), .IN2(n28686), .IN3(n25967), .IN4(n28691), .Q(
        n25873) );
  OA22X1 U29639 ( .IN1(n25945), .IN2(n28692), .IN3(n25963), .IN4(n28687), .Q(
        n25872) );
  OA22X1 U29640 ( .IN1(n25969), .IN2(n28685), .IN3(n25957), .IN4(n28689), .Q(
        n25871) );
  NAND4X0 U29641 ( .IN1(n25874), .IN2(n25873), .IN3(n25872), .IN4(n25871), 
        .QN(s8_addr_o[10]) );
  OA22X1 U29642 ( .IN1(n25945), .IN2(n28702), .IN3(n25958), .IN4(n28700), .Q(
        n25878) );
  OA22X1 U29643 ( .IN1(n25970), .IN2(n28697), .IN3(n25963), .IN4(n28704), .Q(
        n25877) );
  OA22X1 U29644 ( .IN1(n25967), .IN2(n28703), .IN3(n25957), .IN4(n28699), .Q(
        n25876) );
  OA22X1 U29645 ( .IN1(n25968), .IN2(n28698), .IN3(n25969), .IN4(n28701), .Q(
        n25875) );
  NAND4X0 U29646 ( .IN1(n25878), .IN2(n25877), .IN3(n25876), .IN4(n25875), 
        .QN(s8_addr_o[11]) );
  OA22X1 U29647 ( .IN1(n25968), .IN2(n28710), .IN3(n25967), .IN4(n28715), .Q(
        n25882) );
  OA22X1 U29648 ( .IN1(n25945), .IN2(n28714), .IN3(n25957), .IN4(n28713), .Q(
        n25881) );
  OA22X1 U29649 ( .IN1(n25970), .IN2(n28712), .IN3(n25963), .IN4(n28716), .Q(
        n25880) );
  OA22X1 U29650 ( .IN1(n25969), .IN2(n28709), .IN3(n25958), .IN4(n28711), .Q(
        n25879) );
  NAND4X0 U29651 ( .IN1(n25882), .IN2(n25881), .IN3(n25880), .IN4(n25879), 
        .QN(s8_addr_o[12]) );
  OA22X1 U29652 ( .IN1(n25968), .IN2(n28728), .IN3(n25967), .IN4(n28721), .Q(
        n25886) );
  OA22X1 U29653 ( .IN1(n25963), .IN2(n28724), .IN3(n25966), .IN4(n28725), .Q(
        n25885) );
  OA22X1 U29654 ( .IN1(n25945), .IN2(n28722), .IN3(n25957), .IN4(n28727), .Q(
        n25884) );
  OA22X1 U29655 ( .IN1(n25970), .IN2(n28726), .IN3(n25969), .IN4(n28723), .Q(
        n25883) );
  NAND4X0 U29656 ( .IN1(n25886), .IN2(n25885), .IN3(n25884), .IN4(n25883), 
        .QN(s8_addr_o[13]) );
  OA22X1 U29657 ( .IN1(n25969), .IN2(n28740), .IN3(n25957), .IN4(n28739), .Q(
        n25890) );
  OA22X1 U29658 ( .IN1(n25965), .IN2(n28734), .IN3(n25956), .IN4(n28736), .Q(
        n25889) );
  OA22X1 U29659 ( .IN1(n25968), .IN2(n28738), .IN3(n25967), .IN4(n28737), .Q(
        n25888) );
  OA22X1 U29660 ( .IN1(n25932), .IN2(n28735), .IN3(n25958), .IN4(n28733), .Q(
        n25887) );
  NAND4X0 U29661 ( .IN1(n25890), .IN2(n25889), .IN3(n25888), .IN4(n25887), 
        .QN(s8_addr_o[14]) );
  OA22X1 U29662 ( .IN1(n25966), .IN2(n28749), .IN3(n25957), .IN4(n28745), .Q(
        n25894) );
  OA22X1 U29663 ( .IN1(n25932), .IN2(n28752), .IN3(n25967), .IN4(n28751), .Q(
        n25893) );
  OA22X1 U29664 ( .IN1(n25945), .IN2(n28746), .IN3(n25955), .IN4(n28748), .Q(
        n25892) );
  OA22X1 U29665 ( .IN1(n25956), .IN2(n28750), .IN3(n25915), .IN4(n28747), .Q(
        n25891) );
  NAND4X0 U29666 ( .IN1(n25894), .IN2(n25893), .IN3(n25892), .IN4(n25891), 
        .QN(s8_addr_o[15]) );
  OA22X1 U29667 ( .IN1(n25932), .IN2(n28761), .IN3(n25967), .IN4(n28757), .Q(
        n25898) );
  OA22X1 U29668 ( .IN1(n25968), .IN2(n28762), .IN3(n25956), .IN4(n28760), .Q(
        n25897) );
  OA22X1 U29669 ( .IN1(n25945), .IN2(n28758), .IN3(n25964), .IN4(n28763), .Q(
        n25896) );
  OA22X1 U29670 ( .IN1(n25915), .IN2(n28759), .IN3(n25966), .IN4(n28764), .Q(
        n25895) );
  NAND4X0 U29671 ( .IN1(n25898), .IN2(n25897), .IN3(n25896), .IN4(n25895), 
        .QN(s8_addr_o[16]) );
  OA22X1 U29672 ( .IN1(n25963), .IN2(n28773), .IN3(n25966), .IN4(n28770), .Q(
        n25902) );
  OA22X1 U29673 ( .IN1(n25967), .IN2(n28771), .IN3(n25957), .IN4(n28769), .Q(
        n25901) );
  OA22X1 U29674 ( .IN1(n25965), .IN2(n28772), .IN3(n25969), .IN4(n28775), .Q(
        n25900) );
  OA22X1 U29675 ( .IN1(n25955), .IN2(n28776), .IN3(n25956), .IN4(n28774), .Q(
        n25899) );
  NAND4X0 U29676 ( .IN1(n25902), .IN2(n25901), .IN3(n25900), .IN4(n25899), 
        .QN(s8_addr_o[17]) );
  OA22X1 U29677 ( .IN1(n25968), .IN2(n28788), .IN3(n25958), .IN4(n28785), .Q(
        n25906) );
  OA22X1 U29678 ( .IN1(n25932), .IN2(n28782), .IN3(n25964), .IN4(n28781), .Q(
        n25905) );
  OA22X1 U29679 ( .IN1(n25945), .IN2(n28786), .IN3(n25956), .IN4(n28787), .Q(
        n25904) );
  OA22X1 U29680 ( .IN1(n25969), .IN2(n28784), .IN3(n25967), .IN4(n28783), .Q(
        n25903) );
  NAND4X0 U29681 ( .IN1(n25906), .IN2(n25905), .IN3(n25904), .IN4(n25903), 
        .QN(s8_addr_o[18]) );
  OA22X1 U29682 ( .IN1(n25970), .IN2(n28798), .IN3(n25963), .IN4(n28794), .Q(
        n25910) );
  OA22X1 U29683 ( .IN1(n25965), .IN2(n28796), .IN3(n25969), .IN4(n28797), .Q(
        n25909) );
  OA22X1 U29684 ( .IN1(n25955), .IN2(n28800), .IN3(n25967), .IN4(n28795), .Q(
        n25908) );
  OA22X1 U29685 ( .IN1(n25966), .IN2(n28793), .IN3(n25957), .IN4(n28799), .Q(
        n25907) );
  NAND4X0 U29686 ( .IN1(n25910), .IN2(n25909), .IN3(n25908), .IN4(n25907), 
        .QN(s8_addr_o[19]) );
  OA22X1 U29687 ( .IN1(n25932), .IN2(n28810), .IN3(n25969), .IN4(n28806), .Q(
        n25914) );
  OA22X1 U29688 ( .IN1(n25945), .IN2(n28812), .IN3(n25967), .IN4(n28811), .Q(
        n25913) );
  OA22X1 U29689 ( .IN1(n25968), .IN2(n28808), .IN3(n25958), .IN4(n28809), .Q(
        n25912) );
  OA22X1 U29690 ( .IN1(n25970), .IN2(n28807), .IN3(n25964), .IN4(n28805), .Q(
        n25911) );
  NAND4X0 U29691 ( .IN1(n25914), .IN2(n25913), .IN3(n25912), .IN4(n25911), 
        .QN(s8_addr_o[20]) );
  OA22X1 U29692 ( .IN1(n25965), .IN2(n28822), .IN3(n25963), .IN4(n28819), .Q(
        n25919) );
  OA22X1 U29693 ( .IN1(n25950), .IN2(n28823), .IN3(n25966), .IN4(n28818), .Q(
        n25918) );
  OA22X1 U29694 ( .IN1(n25955), .IN2(n28824), .IN3(n25956), .IN4(n28820), .Q(
        n25917) );
  OA22X1 U29695 ( .IN1(n25915), .IN2(n28821), .IN3(n25957), .IN4(n28817), .Q(
        n25916) );
  NAND4X0 U29696 ( .IN1(n25919), .IN2(n25918), .IN3(n25917), .IN4(n25916), 
        .QN(s8_addr_o[21]) );
  OA22X1 U29697 ( .IN1(n25945), .IN2(n28833), .IN3(n25964), .IN4(n28829), .Q(
        n25923) );
  OA22X1 U29698 ( .IN1(n25963), .IN2(n28838), .IN3(n25969), .IN4(n28836), .Q(
        n25922) );
  OA22X1 U29699 ( .IN1(n25968), .IN2(n28832), .IN3(n25956), .IN4(n28831), .Q(
        n25921) );
  OA22X1 U29700 ( .IN1(n25950), .IN2(n28834), .IN3(n25966), .IN4(n28837), .Q(
        n25920) );
  NAND4X0 U29701 ( .IN1(n25923), .IN2(n25922), .IN3(n25921), .IN4(n25920), 
        .QN(s8_addr_o[22]) );
  OA22X1 U29702 ( .IN1(n25955), .IN2(n28845), .IN3(n25969), .IN4(n28852), .Q(
        n25927) );
  OA22X1 U29703 ( .IN1(n25932), .IN2(n28850), .IN3(n25967), .IN4(n28849), .Q(
        n25926) );
  OA22X1 U29704 ( .IN1(n25965), .IN2(n28848), .IN3(n25956), .IN4(n28843), .Q(
        n25925) );
  OA22X1 U29705 ( .IN1(n25966), .IN2(n28846), .IN3(n25957), .IN4(n28851), .Q(
        n25924) );
  NAND4X0 U29706 ( .IN1(n25927), .IN2(n25926), .IN3(n25925), .IN4(n25924), 
        .QN(s8_addr_o[23]) );
  OA22X1 U29707 ( .IN1(n28859), .IN2(n25950), .IN3(n28863), .IN4(n25965), .Q(
        n25931) );
  OA22X1 U29708 ( .IN1(n28860), .IN2(n25957), .IN3(n28857), .IN4(n25963), .Q(
        n25930) );
  OA22X1 U29709 ( .IN1(n28865), .IN2(n25958), .IN3(n28864), .IN4(n25955), .Q(
        n25929) );
  OA22X1 U29710 ( .IN1(n28858), .IN2(n25956), .IN3(n28861), .IN4(n25969), .Q(
        n25928) );
  NAND4X0 U29711 ( .IN1(n25931), .IN2(n25930), .IN3(n25929), .IN4(n25928), 
        .QN(s8_addr_o[24]) );
  OA22X1 U29712 ( .IN1(n28873), .IN2(n25970), .IN3(n28872), .IN4(n25969), .Q(
        n25936) );
  OA22X1 U29713 ( .IN1(n28871), .IN2(n25966), .IN3(n28870), .IN4(n25965), .Q(
        n25935) );
  OA22X1 U29714 ( .IN1(n28875), .IN2(n25964), .IN3(n28874), .IN4(n25932), .Q(
        n25934) );
  OA22X1 U29715 ( .IN1(n28877), .IN2(n25968), .IN3(n28876), .IN4(n25967), .Q(
        n25933) );
  NAND4X0 U29716 ( .IN1(n25936), .IN2(n25935), .IN3(n25934), .IN4(n25933), 
        .QN(s8_addr_o[25]) );
  OA22X1 U29717 ( .IN1(n28885), .IN2(n25956), .IN3(n28884), .IN4(n25965), .Q(
        n25940) );
  OA22X1 U29718 ( .IN1(n28887), .IN2(n25955), .IN3(n28882), .IN4(n25963), .Q(
        n25939) );
  OA22X1 U29719 ( .IN1(n28883), .IN2(n25958), .IN3(n28886), .IN4(n25969), .Q(
        n25938) );
  OA22X1 U29720 ( .IN1(n28889), .IN2(n25957), .IN3(n28888), .IN4(n25967), .Q(
        n25937) );
  NAND4X0 U29721 ( .IN1(n25940), .IN2(n25939), .IN3(n25938), .IN4(n25937), 
        .QN(s8_addr_o[26]) );
  OA22X1 U29722 ( .IN1(n28899), .IN2(n25970), .IN3(n28896), .IN4(n25967), .Q(
        n25944) );
  OA22X1 U29723 ( .IN1(n28897), .IN2(n25966), .IN3(n28898), .IN4(n25964), .Q(
        n25943) );
  OA22X1 U29724 ( .IN1(n28895), .IN2(n25968), .IN3(n28894), .IN4(n25965), .Q(
        n25942) );
  OA22X1 U29725 ( .IN1(n28901), .IN2(n25963), .IN3(n28900), .IN4(n25969), .Q(
        n25941) );
  NAND4X0 U29726 ( .IN1(n25944), .IN2(n25943), .IN3(n25942), .IN4(n25941), 
        .QN(s8_addr_o[27]) );
  OA22X1 U29727 ( .IN1(n28912), .IN2(n25945), .IN3(n28908), .IN4(n25963), .Q(
        n25949) );
  OA22X1 U29728 ( .IN1(n28909), .IN2(n25956), .IN3(n28911), .IN4(n25955), .Q(
        n25948) );
  OA22X1 U29729 ( .IN1(n28913), .IN2(n25964), .IN3(n28910), .IN4(n25967), .Q(
        n25947) );
  OA22X1 U29730 ( .IN1(n28907), .IN2(n25958), .IN3(n28906), .IN4(n25969), .Q(
        n25946) );
  NAND4X0 U29731 ( .IN1(n25949), .IN2(n25948), .IN3(n25947), .IN4(n25946), 
        .QN(s8_addr_o[28]) );
  OA22X1 U29732 ( .IN1(n28922), .IN2(n25966), .IN3(n28921), .IN4(n25957), .Q(
        n25954) );
  OA22X1 U29733 ( .IN1(n28926), .IN2(n25970), .IN3(n28923), .IN4(n25969), .Q(
        n25953) );
  OA22X1 U29734 ( .IN1(n28920), .IN2(n25950), .IN3(n28919), .IN4(n25963), .Q(
        n25952) );
  OA22X1 U29735 ( .IN1(n28924), .IN2(n25955), .IN3(n28925), .IN4(n25965), .Q(
        n25951) );
  NAND4X0 U29736 ( .IN1(n25954), .IN2(n25953), .IN3(n25952), .IN4(n25951), 
        .QN(s8_addr_o[29]) );
  OA22X1 U29737 ( .IN1(n28932), .IN2(n25956), .IN3(n28935), .IN4(n25955), .Q(
        n25962) );
  OA22X1 U29738 ( .IN1(n28931), .IN2(n25965), .IN3(n28940), .IN4(n25963), .Q(
        n25961) );
  OA22X1 U29739 ( .IN1(n28933), .IN2(n25957), .IN3(n28936), .IN4(n25967), .Q(
        n25960) );
  OA22X1 U29740 ( .IN1(n28937), .IN2(n25958), .IN3(n28939), .IN4(n25969), .Q(
        n25959) );
  NAND4X0 U29741 ( .IN1(n25962), .IN2(n25961), .IN3(n25960), .IN4(n25959), 
        .QN(s8_addr_o[30]) );
  OA22X1 U29742 ( .IN1(n28960), .IN2(n25964), .IN3(n28958), .IN4(n25963), .Q(
        n25974) );
  OA22X1 U29743 ( .IN1(n28956), .IN2(n25966), .IN3(n28950), .IN4(n25965), .Q(
        n25973) );
  OA22X1 U29744 ( .IN1(n28952), .IN2(n25968), .IN3(n28954), .IN4(n25967), .Q(
        n25972) );
  OA22X1 U29745 ( .IN1(n28948), .IN2(n25970), .IN3(n28946), .IN4(n25969), .Q(
        n25971) );
  NAND4X0 U29746 ( .IN1(n25974), .IN2(n25973), .IN3(n25972), .IN4(n25971), 
        .QN(s8_addr_o[31]) );
  OA22X1 U29747 ( .IN1(n29330), .IN2(n25976), .IN3(n29311), .IN4(n25975), .Q(
        n25986) );
  OA22X1 U29748 ( .IN1(n29235), .IN2(n25978), .IN3(n29292), .IN4(n25977), .Q(
        n25985) );
  OA22X1 U29749 ( .IN1(n29349), .IN2(n25980), .IN3(n29254), .IN4(n25979), .Q(
        n25984) );
  OA22X1 U29750 ( .IN1(n29273), .IN2(n25982), .IN3(n29368), .IN4(n25981), .Q(
        n25983) );
  NAND4X0 U29751 ( .IN1(n25986), .IN2(n25985), .IN3(n25984), .IN4(n25983), 
        .QN(s7_stb_o) );
  INVX0 U29752 ( .INP(n29091), .ZN(n26262) );
  INVX0 U29753 ( .INP(n29100), .ZN(n26274) );
  OA22X1 U29754 ( .IN1(n26262), .IN2(n28123), .IN3(n26274), .IN4(n28127), .Q(
        n25990) );
  INVX0 U29755 ( .INP(n29092), .ZN(n26253) );
  INVX0 U29756 ( .INP(n29094), .ZN(n26269) );
  OA22X1 U29757 ( .IN1(n26253), .IN2(n28126), .IN3(n26269), .IN4(n28125), .Q(
        n25989) );
  INVX0 U29758 ( .INP(n29099), .ZN(n26272) );
  INVX0 U29759 ( .INP(n29101), .ZN(n26227) );
  OA22X1 U29760 ( .IN1(n26272), .IN2(n28124), .IN3(n26227), .IN4(n28122), .Q(
        n25988) );
  INVX0 U29761 ( .INP(n29093), .ZN(n26236) );
  INVX0 U29762 ( .INP(n29102), .ZN(n26261) );
  OA22X1 U29763 ( .IN1(n26236), .IN2(n28128), .IN3(n26261), .IN4(n28121), .Q(
        n25987) );
  NAND4X0 U29764 ( .IN1(n25990), .IN2(n25989), .IN3(n25988), .IN4(n25987), 
        .QN(s7_we_o) );
  INVX0 U29765 ( .INP(n29091), .ZN(n26270) );
  OA22X1 U29766 ( .IN1(n26270), .IN2(n28133), .IN3(n26227), .IN4(n28138), .Q(
        n25994) );
  INVX0 U29767 ( .INP(n29093), .ZN(n26268) );
  OA22X1 U29768 ( .IN1(n26268), .IN2(n28140), .IN3(n26269), .IN4(n28136), .Q(
        n25993) );
  OA22X1 U29769 ( .IN1(n26272), .IN2(n28134), .IN3(n26253), .IN4(n28139), .Q(
        n25992) );
  INVX0 U29770 ( .INP(n29100), .ZN(n26260) );
  INVX0 U29771 ( .INP(n29102), .ZN(n26273) );
  OA22X1 U29772 ( .IN1(n26260), .IN2(n28137), .IN3(n26273), .IN4(n28135), .Q(
        n25991) );
  NAND4X0 U29773 ( .IN1(n25994), .IN2(n25993), .IN3(n25992), .IN4(n25991), 
        .QN(s7_data_o[0]) );
  OA22X1 U29774 ( .IN1(n26236), .IN2(n28146), .IN3(n26227), .IN4(n28149), .Q(
        n25998) );
  OA22X1 U29775 ( .IN1(n26270), .IN2(n28148), .IN3(n26273), .IN4(n28147), .Q(
        n25997) );
  INVX0 U29776 ( .INP(n29092), .ZN(n26267) );
  OA22X1 U29777 ( .IN1(n26267), .IN2(n28145), .IN3(n26269), .IN4(n28152), .Q(
        n25996) );
  INVX0 U29778 ( .INP(n29099), .ZN(n26258) );
  OA22X1 U29779 ( .IN1(n26258), .IN2(n28150), .IN3(n26274), .IN4(n28151), .Q(
        n25995) );
  NAND4X0 U29780 ( .IN1(n25998), .IN2(n25997), .IN3(n25996), .IN4(n25995), 
        .QN(s7_data_o[1]) );
  OA22X1 U29781 ( .IN1(n26258), .IN2(n28160), .IN3(n26274), .IN4(n28157), .Q(
        n26002) );
  OA22X1 U29782 ( .IN1(n26253), .IN2(n28159), .IN3(n26269), .IN4(n28162), .Q(
        n26001) );
  OA22X1 U29783 ( .IN1(n26236), .IN2(n28164), .IN3(n26227), .IN4(n28158), .Q(
        n26000) );
  OA22X1 U29784 ( .IN1(n26270), .IN2(n28163), .IN3(n26273), .IN4(n28161), .Q(
        n25999) );
  NAND4X0 U29785 ( .IN1(n26002), .IN2(n26001), .IN3(n26000), .IN4(n25999), 
        .QN(s7_data_o[2]) );
  INVX0 U29786 ( .INP(n29101), .ZN(n26271) );
  OA22X1 U29787 ( .IN1(n26271), .IN2(n28171), .IN3(n26274), .IN4(n28169), .Q(
        n26006) );
  OA22X1 U29788 ( .IN1(n26258), .IN2(n28172), .IN3(n26269), .IN4(n28175), .Q(
        n26005) );
  OA22X1 U29789 ( .IN1(n26236), .IN2(n28174), .IN3(n26273), .IN4(n28173), .Q(
        n26004) );
  OA22X1 U29790 ( .IN1(n26270), .IN2(n28176), .IN3(n26253), .IN4(n28170), .Q(
        n26003) );
  NAND4X0 U29791 ( .IN1(n26006), .IN2(n26005), .IN3(n26004), .IN4(n26003), 
        .QN(s7_data_o[3]) );
  OA22X1 U29792 ( .IN1(n26258), .IN2(n28182), .IN3(n26273), .IN4(n28181), .Q(
        n26010) );
  OA22X1 U29793 ( .IN1(n26236), .IN2(n28184), .IN3(n26253), .IN4(n28188), .Q(
        n26009) );
  OA22X1 U29794 ( .IN1(n26262), .IN2(n28186), .IN3(n26274), .IN4(n28187), .Q(
        n26008) );
  OA22X1 U29795 ( .IN1(n26271), .IN2(n28185), .IN3(n26269), .IN4(n28183), .Q(
        n26007) );
  NAND4X0 U29796 ( .IN1(n26010), .IN2(n26009), .IN3(n26008), .IN4(n26007), 
        .QN(s7_data_o[4]) );
  OA22X1 U29797 ( .IN1(n26267), .IN2(n28193), .IN3(n26227), .IN4(n28198), .Q(
        n26014) );
  OA22X1 U29798 ( .IN1(n26258), .IN2(n28196), .IN3(n26273), .IN4(n28199), .Q(
        n26013) );
  OA22X1 U29799 ( .IN1(n26236), .IN2(n28200), .IN3(n26269), .IN4(n28197), .Q(
        n26012) );
  OA22X1 U29800 ( .IN1(n26262), .IN2(n28194), .IN3(n26274), .IN4(n28195), .Q(
        n26011) );
  NAND4X0 U29801 ( .IN1(n26014), .IN2(n26013), .IN3(n26012), .IN4(n26011), 
        .QN(s7_data_o[5]) );
  OA22X1 U29802 ( .IN1(n26269), .IN2(n28205), .IN3(n26274), .IN4(n28210), .Q(
        n26018) );
  OA22X1 U29803 ( .IN1(n26236), .IN2(n28207), .IN3(n26273), .IN4(n28209), .Q(
        n26017) );
  OA22X1 U29804 ( .IN1(n26253), .IN2(n28212), .IN3(n26227), .IN4(n28211), .Q(
        n26016) );
  OA22X1 U29805 ( .IN1(n26258), .IN2(n28208), .IN3(n26270), .IN4(n28206), .Q(
        n26015) );
  NAND4X0 U29806 ( .IN1(n26018), .IN2(n26017), .IN3(n26016), .IN4(n26015), 
        .QN(s7_data_o[6]) );
  OA22X1 U29807 ( .IN1(n26267), .IN2(n28218), .IN3(n26269), .IN4(n28223), .Q(
        n26022) );
  OA22X1 U29808 ( .IN1(n26262), .IN2(n28224), .IN3(n26227), .IN4(n28217), .Q(
        n26021) );
  OA22X1 U29809 ( .IN1(n26274), .IN2(n28222), .IN3(n26261), .IN4(n28221), .Q(
        n26020) );
  OA22X1 U29810 ( .IN1(n26258), .IN2(n28220), .IN3(n26236), .IN4(n28219), .Q(
        n26019) );
  NAND4X0 U29811 ( .IN1(n26022), .IN2(n26021), .IN3(n26020), .IN4(n26019), 
        .QN(s7_data_o[7]) );
  OA22X1 U29812 ( .IN1(n26253), .IN2(n28234), .IN3(n26269), .IN4(n28229), .Q(
        n26026) );
  OA22X1 U29813 ( .IN1(n26272), .IN2(n28230), .IN3(n26274), .IN4(n28233), .Q(
        n26025) );
  OA22X1 U29814 ( .IN1(n26236), .IN2(n28232), .IN3(n26270), .IN4(n28231), .Q(
        n26024) );
  OA22X1 U29815 ( .IN1(n26227), .IN2(n28236), .IN3(n26261), .IN4(n28235), .Q(
        n26023) );
  NAND4X0 U29816 ( .IN1(n26026), .IN2(n26025), .IN3(n26024), .IN4(n26023), 
        .QN(s7_data_o[8]) );
  OA22X1 U29817 ( .IN1(n26272), .IN2(n28242), .IN3(n26227), .IN4(n28241), .Q(
        n26030) );
  OA22X1 U29818 ( .IN1(n26236), .IN2(n28244), .IN3(n26261), .IN4(n28247), .Q(
        n26029) );
  OA22X1 U29819 ( .IN1(n26267), .IN2(n28248), .IN3(n26269), .IN4(n28245), .Q(
        n26028) );
  OA22X1 U29820 ( .IN1(n26270), .IN2(n28246), .IN3(n26274), .IN4(n28243), .Q(
        n26027) );
  NAND4X0 U29821 ( .IN1(n26030), .IN2(n26029), .IN3(n26028), .IN4(n26027), 
        .QN(s7_data_o[9]) );
  OA22X1 U29822 ( .IN1(n26262), .IN2(n28260), .IN3(n26227), .IN4(n28254), .Q(
        n26034) );
  OA22X1 U29823 ( .IN1(n26272), .IN2(n28258), .IN3(n26236), .IN4(n28257), .Q(
        n26033) );
  OA22X1 U29824 ( .IN1(n26253), .IN2(n28256), .IN3(n26274), .IN4(n28253), .Q(
        n26032) );
  INVX0 U29825 ( .INP(n29094), .ZN(n26259) );
  OA22X1 U29826 ( .IN1(n26259), .IN2(n28255), .IN3(n26261), .IN4(n28259), .Q(
        n26031) );
  NAND4X0 U29827 ( .IN1(n26034), .IN2(n26033), .IN3(n26032), .IN4(n26031), 
        .QN(s7_data_o[10]) );
  OA22X1 U29828 ( .IN1(n26262), .IN2(n28265), .IN3(n26269), .IN4(n28270), .Q(
        n26038) );
  OA22X1 U29829 ( .IN1(n26271), .IN2(n28268), .IN3(n26261), .IN4(n28269), .Q(
        n26037) );
  OA22X1 U29830 ( .IN1(n26272), .IN2(n28266), .IN3(n26260), .IN4(n28267), .Q(
        n26036) );
  OA22X1 U29831 ( .IN1(n26268), .IN2(n28272), .IN3(n26253), .IN4(n28271), .Q(
        n26035) );
  NAND4X0 U29832 ( .IN1(n26038), .IN2(n26037), .IN3(n26036), .IN4(n26035), 
        .QN(s7_data_o[11]) );
  OA22X1 U29833 ( .IN1(n26262), .IN2(n28280), .IN3(n26261), .IN4(n28277), .Q(
        n26042) );
  OA22X1 U29834 ( .IN1(n26236), .IN2(n28278), .IN3(n26260), .IN4(n28279), .Q(
        n26041) );
  OA22X1 U29835 ( .IN1(n26267), .IN2(n28282), .IN3(n26227), .IN4(n28283), .Q(
        n26040) );
  OA22X1 U29836 ( .IN1(n26272), .IN2(n28284), .IN3(n26259), .IN4(n28281), .Q(
        n26039) );
  NAND4X0 U29837 ( .IN1(n26042), .IN2(n26041), .IN3(n26040), .IN4(n26039), 
        .QN(s7_data_o[12]) );
  OA22X1 U29838 ( .IN1(n26272), .IN2(n28290), .IN3(n26253), .IN4(n28292), .Q(
        n26046) );
  OA22X1 U29839 ( .IN1(n26268), .IN2(n28294), .IN3(n26227), .IN4(n28289), .Q(
        n26045) );
  OA22X1 U29840 ( .IN1(n26260), .IN2(n28291), .IN3(n26261), .IN4(n28295), .Q(
        n26044) );
  OA22X1 U29841 ( .IN1(n26270), .IN2(n28296), .IN3(n26259), .IN4(n28293), .Q(
        n26043) );
  NAND4X0 U29842 ( .IN1(n26046), .IN2(n26045), .IN3(n26044), .IN4(n26043), 
        .QN(s7_data_o[13]) );
  OA22X1 U29843 ( .IN1(n26272), .IN2(n28306), .IN3(n26253), .IN4(n28305), .Q(
        n26050) );
  OA22X1 U29844 ( .IN1(n26227), .IN2(n28307), .IN3(n26260), .IN4(n28301), .Q(
        n26049) );
  OA22X1 U29845 ( .IN1(n26236), .IN2(n28304), .IN3(n26261), .IN4(n28303), .Q(
        n26048) );
  OA22X1 U29846 ( .IN1(n26270), .IN2(n28308), .IN3(n26269), .IN4(n28302), .Q(
        n26047) );
  NAND4X0 U29847 ( .IN1(n26050), .IN2(n26049), .IN3(n26048), .IN4(n26047), 
        .QN(s7_data_o[14]) );
  OA22X1 U29848 ( .IN1(n26272), .IN2(n28316), .IN3(n26270), .IN4(n28314), .Q(
        n26054) );
  OA22X1 U29849 ( .IN1(n26269), .IN2(n28318), .IN3(n26261), .IN4(n28319), .Q(
        n26053) );
  OA22X1 U29850 ( .IN1(n26271), .IN2(n28320), .IN3(n26260), .IN4(n28317), .Q(
        n26052) );
  OA22X1 U29851 ( .IN1(n26268), .IN2(n28315), .IN3(n26253), .IN4(n28313), .Q(
        n26051) );
  NAND4X0 U29852 ( .IN1(n26054), .IN2(n26053), .IN3(n26052), .IN4(n26051), 
        .QN(s7_data_o[15]) );
  OA22X1 U29853 ( .IN1(n26272), .IN2(n28330), .IN3(n26259), .IN4(n28325), .Q(
        n26058) );
  OA22X1 U29854 ( .IN1(n26262), .IN2(n28331), .IN3(n26253), .IN4(n28326), .Q(
        n26057) );
  OA22X1 U29855 ( .IN1(n26236), .IN2(n28332), .IN3(n26261), .IN4(n28327), .Q(
        n26056) );
  OA22X1 U29856 ( .IN1(n26227), .IN2(n28329), .IN3(n26260), .IN4(n28328), .Q(
        n26055) );
  NAND4X0 U29857 ( .IN1(n26058), .IN2(n26057), .IN3(n26056), .IN4(n26055), 
        .QN(s7_data_o[16]) );
  OA22X1 U29858 ( .IN1(n26270), .IN2(n28342), .IN3(n26227), .IN4(n28337), .Q(
        n26062) );
  OA22X1 U29859 ( .IN1(n26268), .IN2(n28344), .IN3(n26253), .IN4(n28338), .Q(
        n26061) );
  OA22X1 U29860 ( .IN1(n26274), .IN2(n28343), .IN3(n26261), .IN4(n28341), .Q(
        n26060) );
  OA22X1 U29861 ( .IN1(n26272), .IN2(n28340), .IN3(n26269), .IN4(n28339), .Q(
        n26059) );
  NAND4X0 U29862 ( .IN1(n26062), .IN2(n26061), .IN3(n26060), .IN4(n26059), 
        .QN(s7_data_o[17]) );
  OA22X1 U29863 ( .IN1(n26272), .IN2(n28352), .IN3(n26269), .IN4(n28349), .Q(
        n26066) );
  OA22X1 U29864 ( .IN1(n26270), .IN2(n28350), .IN3(n26227), .IN4(n28354), .Q(
        n26065) );
  OA22X1 U29865 ( .IN1(n26253), .IN2(n28355), .IN3(n26261), .IN4(n28353), .Q(
        n26064) );
  OA22X1 U29866 ( .IN1(n26236), .IN2(n28356), .IN3(n26260), .IN4(n28351), .Q(
        n26063) );
  NAND4X0 U29867 ( .IN1(n26066), .IN2(n26065), .IN3(n26064), .IN4(n26063), 
        .QN(s7_data_o[18]) );
  OA22X1 U29868 ( .IN1(n26267), .IN2(n28363), .IN3(n26227), .IN4(n28365), .Q(
        n26070) );
  OA22X1 U29869 ( .IN1(n26262), .IN2(n28362), .IN3(n26269), .IN4(n28361), .Q(
        n26069) );
  OA22X1 U29870 ( .IN1(n26272), .IN2(n28366), .IN3(n26261), .IN4(n28367), .Q(
        n26068) );
  OA22X1 U29871 ( .IN1(n26268), .IN2(n28364), .IN3(n26260), .IN4(n28368), .Q(
        n26067) );
  NAND4X0 U29872 ( .IN1(n26070), .IN2(n26069), .IN3(n26068), .IN4(n26067), 
        .QN(s7_data_o[19]) );
  OA22X1 U29873 ( .IN1(n26259), .IN2(n28380), .IN3(n26260), .IN4(n28379), .Q(
        n26074) );
  OA22X1 U29874 ( .IN1(n26271), .IN2(n28376), .IN3(n26261), .IN4(n28375), .Q(
        n26073) );
  OA22X1 U29875 ( .IN1(n26272), .IN2(n28378), .IN3(n26236), .IN4(n28377), .Q(
        n26072) );
  OA22X1 U29876 ( .IN1(n26262), .IN2(n28374), .IN3(n26253), .IN4(n28373), .Q(
        n26071) );
  NAND4X0 U29877 ( .IN1(n26074), .IN2(n26073), .IN3(n26072), .IN4(n26071), 
        .QN(s7_data_o[20]) );
  OA22X1 U29878 ( .IN1(n26236), .IN2(n28386), .IN3(n26270), .IN4(n28390), .Q(
        n26078) );
  OA22X1 U29879 ( .IN1(n26267), .IN2(n28388), .IN3(n26227), .IN4(n28387), .Q(
        n26077) );
  OA22X1 U29880 ( .IN1(n26272), .IN2(n28392), .IN3(n26261), .IN4(n28391), .Q(
        n26076) );
  OA22X1 U29881 ( .IN1(n26259), .IN2(n28385), .IN3(n26260), .IN4(n28389), .Q(
        n26075) );
  NAND4X0 U29882 ( .IN1(n26078), .IN2(n26077), .IN3(n26076), .IN4(n26075), 
        .QN(s7_data_o[21]) );
  OA22X1 U29883 ( .IN1(n26268), .IN2(n28402), .IN3(n26270), .IN4(n28404), .Q(
        n26082) );
  OA22X1 U29884 ( .IN1(n26258), .IN2(n28400), .IN3(n26261), .IN4(n28397), .Q(
        n26081) );
  OA22X1 U29885 ( .IN1(n26267), .IN2(n28403), .IN3(n26260), .IN4(n28401), .Q(
        n26080) );
  OA22X1 U29886 ( .IN1(n26271), .IN2(n28398), .IN3(n26259), .IN4(n28399), .Q(
        n26079) );
  NAND4X0 U29887 ( .IN1(n26082), .IN2(n26081), .IN3(n26080), .IN4(n26079), 
        .QN(s7_data_o[22]) );
  OA22X1 U29888 ( .IN1(n26236), .IN2(n28415), .IN3(n26260), .IN4(n28409), .Q(
        n26086) );
  OA22X1 U29889 ( .IN1(n26272), .IN2(n28416), .IN3(n26273), .IN4(n28411), .Q(
        n26085) );
  OA22X1 U29890 ( .IN1(n26270), .IN2(n28414), .IN3(n26227), .IN4(n28410), .Q(
        n26084) );
  OA22X1 U29891 ( .IN1(n26267), .IN2(n28413), .IN3(n26259), .IN4(n28412), .Q(
        n26083) );
  NAND4X0 U29892 ( .IN1(n26086), .IN2(n26085), .IN3(n26084), .IN4(n26083), 
        .QN(s7_data_o[23]) );
  OA22X1 U29893 ( .IN1(n26262), .IN2(n28422), .IN3(n26261), .IN4(n28423), .Q(
        n26090) );
  OA22X1 U29894 ( .IN1(n26272), .IN2(n28426), .IN3(n26253), .IN4(n28421), .Q(
        n26089) );
  OA22X1 U29895 ( .IN1(n26271), .IN2(n28425), .IN3(n26260), .IN4(n28427), .Q(
        n26088) );
  OA22X1 U29896 ( .IN1(n26236), .IN2(n28424), .IN3(n26269), .IN4(n28428), .Q(
        n26087) );
  NAND4X0 U29897 ( .IN1(n26090), .IN2(n26089), .IN3(n26088), .IN4(n26087), 
        .QN(s7_data_o[24]) );
  OA22X1 U29898 ( .IN1(n26236), .IN2(n28440), .IN3(n26253), .IN4(n28439), .Q(
        n26094) );
  OA22X1 U29899 ( .IN1(n26258), .IN2(n28438), .IN3(n26262), .IN4(n28434), .Q(
        n26093) );
  OA22X1 U29900 ( .IN1(n26259), .IN2(n28437), .IN3(n26273), .IN4(n28435), .Q(
        n26092) );
  OA22X1 U29901 ( .IN1(n26227), .IN2(n28433), .IN3(n26260), .IN4(n28436), .Q(
        n26091) );
  NAND4X0 U29902 ( .IN1(n26094), .IN2(n26093), .IN3(n26092), .IN4(n26091), 
        .QN(s7_data_o[25]) );
  OA22X1 U29903 ( .IN1(n26259), .IN2(n28448), .IN3(n26260), .IN4(n28447), .Q(
        n26098) );
  OA22X1 U29904 ( .IN1(n26270), .IN2(n28450), .IN3(n26227), .IN4(n28449), .Q(
        n26097) );
  OA22X1 U29905 ( .IN1(n26258), .IN2(n28452), .IN3(n26267), .IN4(n28446), .Q(
        n26096) );
  OA22X1 U29906 ( .IN1(n26236), .IN2(n28451), .IN3(n26273), .IN4(n28445), .Q(
        n26095) );
  NAND4X0 U29907 ( .IN1(n26098), .IN2(n26097), .IN3(n26096), .IN4(n26095), 
        .QN(s7_data_o[26]) );
  OA22X1 U29908 ( .IN1(n26272), .IN2(n28462), .IN3(n26270), .IN4(n28464), .Q(
        n26102) );
  OA22X1 U29909 ( .IN1(n26236), .IN2(n28461), .IN3(n26227), .IN4(n28457), .Q(
        n26101) );
  OA22X1 U29910 ( .IN1(n26259), .IN2(n28463), .IN3(n26261), .IN4(n28459), .Q(
        n26100) );
  OA22X1 U29911 ( .IN1(n26267), .IN2(n28458), .IN3(n26260), .IN4(n28460), .Q(
        n26099) );
  NAND4X0 U29912 ( .IN1(n26102), .IN2(n26101), .IN3(n26100), .IN4(n26099), 
        .QN(s7_data_o[27]) );
  OA22X1 U29913 ( .IN1(n26258), .IN2(n28474), .IN3(n26227), .IN4(n28471), .Q(
        n26106) );
  OA22X1 U29914 ( .IN1(n26274), .IN2(n28469), .IN3(n26261), .IN4(n28473), .Q(
        n26105) );
  OA22X1 U29915 ( .IN1(n26253), .IN2(n28470), .IN3(n26269), .IN4(n28475), .Q(
        n26104) );
  OA22X1 U29916 ( .IN1(n26268), .IN2(n28476), .IN3(n26270), .IN4(n28472), .Q(
        n26103) );
  NAND4X0 U29917 ( .IN1(n26106), .IN2(n26105), .IN3(n26104), .IN4(n26103), 
        .QN(s7_data_o[28]) );
  OA22X1 U29918 ( .IN1(n26268), .IN2(n28482), .IN3(n26260), .IN4(n28485), .Q(
        n26110) );
  OA22X1 U29919 ( .IN1(n26272), .IN2(n28484), .IN3(n26262), .IN4(n28488), .Q(
        n26109) );
  OA22X1 U29920 ( .IN1(n26271), .IN2(n28487), .IN3(n26259), .IN4(n28483), .Q(
        n26108) );
  OA22X1 U29921 ( .IN1(n26253), .IN2(n28486), .IN3(n26273), .IN4(n28481), .Q(
        n26107) );
  NAND4X0 U29922 ( .IN1(n26110), .IN2(n26109), .IN3(n26108), .IN4(n26107), 
        .QN(s7_data_o[29]) );
  OA22X1 U29923 ( .IN1(n26270), .IN2(n28497), .IN3(n26260), .IN4(n28500), .Q(
        n26114) );
  OA22X1 U29924 ( .IN1(n26272), .IN2(n28494), .IN3(n26269), .IN4(n28495), .Q(
        n26113) );
  OA22X1 U29925 ( .IN1(n26267), .IN2(n28496), .IN3(n26261), .IN4(n28499), .Q(
        n26112) );
  OA22X1 U29926 ( .IN1(n26268), .IN2(n28498), .IN3(n26271), .IN4(n28493), .Q(
        n26111) );
  NAND4X0 U29927 ( .IN1(n26114), .IN2(n26113), .IN3(n26112), .IN4(n26111), 
        .QN(s7_data_o[30]) );
  OA22X1 U29928 ( .IN1(n26262), .IN2(n28506), .IN3(n26260), .IN4(n28511), .Q(
        n26118) );
  OA22X1 U29929 ( .IN1(n26253), .IN2(n28505), .IN3(n26227), .IN4(n28512), .Q(
        n26117) );
  OA22X1 U29930 ( .IN1(n26259), .IN2(n28508), .IN3(n26273), .IN4(n28507), .Q(
        n26116) );
  OA22X1 U29931 ( .IN1(n26258), .IN2(n28510), .IN3(n26236), .IN4(n28509), .Q(
        n26115) );
  NAND4X0 U29932 ( .IN1(n26118), .IN2(n26117), .IN3(n26116), .IN4(n26115), 
        .QN(s7_data_o[31]) );
  OA22X1 U29933 ( .IN1(n26258), .IN2(n28518), .IN3(n26259), .IN4(n28520), .Q(
        n26122) );
  OA22X1 U29934 ( .IN1(n26253), .IN2(n28524), .IN3(n26274), .IN4(n28521), .Q(
        n26121) );
  OA22X1 U29935 ( .IN1(n26236), .IN2(n28517), .IN3(n26273), .IN4(n28519), .Q(
        n26120) );
  OA22X1 U29936 ( .IN1(n26262), .IN2(n28522), .IN3(n26227), .IN4(n28523), .Q(
        n26119) );
  NAND4X0 U29937 ( .IN1(n26122), .IN2(n26121), .IN3(n26120), .IN4(n26119), 
        .QN(s7_sel_o[0]) );
  OA22X1 U29938 ( .IN1(n26262), .IN2(n28530), .IN3(n26267), .IN4(n28536), .Q(
        n26126) );
  OA22X1 U29939 ( .IN1(n26227), .IN2(n28535), .IN3(n26269), .IN4(n28533), .Q(
        n26125) );
  OA22X1 U29940 ( .IN1(n26272), .IN2(n28534), .IN3(n26261), .IN4(n28529), .Q(
        n26124) );
  OA22X1 U29941 ( .IN1(n26268), .IN2(n28532), .IN3(n26274), .IN4(n28531), .Q(
        n26123) );
  NAND4X0 U29942 ( .IN1(n26126), .IN2(n26125), .IN3(n26124), .IN4(n26123), 
        .QN(s7_sel_o[1]) );
  OA22X1 U29943 ( .IN1(n26259), .IN2(n28542), .IN3(n26261), .IN4(n28541), .Q(
        n26130) );
  OA22X1 U29944 ( .IN1(n26258), .IN2(n28544), .IN3(n26253), .IN4(n28548), .Q(
        n26129) );
  OA22X1 U29945 ( .IN1(n26262), .IN2(n28543), .IN3(n26260), .IN4(n28545), .Q(
        n26128) );
  OA22X1 U29946 ( .IN1(n26236), .IN2(n28546), .IN3(n26271), .IN4(n28547), .Q(
        n26127) );
  NAND4X0 U29947 ( .IN1(n26130), .IN2(n26129), .IN3(n26128), .IN4(n26127), 
        .QN(s7_sel_o[2]) );
  OA22X1 U29948 ( .IN1(n26262), .IN2(n28553), .IN3(n26271), .IN4(n28556), .Q(
        n26134) );
  OA22X1 U29949 ( .IN1(n26253), .IN2(n28557), .IN3(n26274), .IN4(n28559), .Q(
        n26133) );
  OA22X1 U29950 ( .IN1(n26258), .IN2(n28558), .IN3(n26259), .IN4(n28560), .Q(
        n26132) );
  OA22X1 U29951 ( .IN1(n26268), .IN2(n28554), .IN3(n26273), .IN4(n28555), .Q(
        n26131) );
  NAND4X0 U29952 ( .IN1(n26134), .IN2(n26133), .IN3(n26132), .IN4(n26131), 
        .QN(s7_sel_o[3]) );
  OA22X1 U29953 ( .IN1(n26259), .IN2(n28567), .IN3(n26260), .IN4(n28565), .Q(
        n26138) );
  OA22X1 U29954 ( .IN1(n26272), .IN2(n28572), .IN3(n26267), .IN4(n28566), .Q(
        n26137) );
  OA22X1 U29955 ( .IN1(n26271), .IN2(n28568), .IN3(n26261), .IN4(n28569), .Q(
        n26136) );
  OA22X1 U29956 ( .IN1(n26236), .IN2(n28570), .IN3(n26270), .IN4(n28571), .Q(
        n26135) );
  NAND4X0 U29957 ( .IN1(n26138), .IN2(n26137), .IN3(n26136), .IN4(n26135), 
        .QN(s7_addr_o[0]) );
  OA22X1 U29958 ( .IN1(n26268), .IN2(n28578), .IN3(n26270), .IN4(n28582), .Q(
        n26142) );
  OA22X1 U29959 ( .IN1(n26272), .IN2(n28580), .IN3(n26271), .IN4(n28579), .Q(
        n26141) );
  OA22X1 U29960 ( .IN1(n26274), .IN2(n28577), .IN3(n26273), .IN4(n28583), .Q(
        n26140) );
  OA22X1 U29961 ( .IN1(n26253), .IN2(n28581), .IN3(n26259), .IN4(n28584), .Q(
        n26139) );
  NAND4X0 U29962 ( .IN1(n26142), .IN2(n26141), .IN3(n26140), .IN4(n26139), 
        .QN(s7_addr_o[1]) );
  OA22X1 U29963 ( .IN1(n28596), .IN2(n26261), .IN3(n28593), .IN4(n26269), .Q(
        n26146) );
  OA22X1 U29964 ( .IN1(n28592), .IN2(n26253), .IN3(n28590), .IN4(n26227), .Q(
        n26145) );
  OA22X1 U29965 ( .IN1(n28594), .IN2(n26270), .IN3(n28589), .IN4(n26236), .Q(
        n26144) );
  OA22X1 U29966 ( .IN1(n28591), .IN2(n26272), .IN3(n28595), .IN4(n26274), .Q(
        n26143) );
  NAND4X0 U29967 ( .IN1(n26146), .IN2(n26145), .IN3(n26144), .IN4(n26143), 
        .QN(s7_addr_o[2]) );
  OA22X1 U29968 ( .IN1(n28606), .IN2(n26227), .IN3(n28603), .IN4(n26274), .Q(
        n26150) );
  OA22X1 U29969 ( .IN1(n28604), .IN2(n26262), .IN3(n28607), .IN4(n26267), .Q(
        n26149) );
  OA22X1 U29970 ( .IN1(n28605), .IN2(n26268), .IN3(n28608), .IN4(n26273), .Q(
        n26148) );
  OA22X1 U29971 ( .IN1(n28602), .IN2(n26269), .IN3(n28601), .IN4(n26258), .Q(
        n26147) );
  NAND4X0 U29972 ( .IN1(n26150), .IN2(n26149), .IN3(n26148), .IN4(n26147), 
        .QN(s7_addr_o[3]) );
  OA22X1 U29973 ( .IN1(n28618), .IN2(n26267), .IN3(n28617), .IN4(n26258), .Q(
        n26154) );
  OA22X1 U29974 ( .IN1(n28619), .IN2(n26273), .IN3(n28615), .IN4(n26271), .Q(
        n26153) );
  OA22X1 U29975 ( .IN1(n28616), .IN2(n26268), .IN3(n28620), .IN4(n26274), .Q(
        n26152) );
  OA22X1 U29976 ( .IN1(n28614), .IN2(n26259), .IN3(n28613), .IN4(n26262), .Q(
        n26151) );
  NAND4X0 U29977 ( .IN1(n26154), .IN2(n26153), .IN3(n26152), .IN4(n26151), 
        .QN(s7_addr_o[4]) );
  OA22X1 U29978 ( .IN1(n28628), .IN2(n26260), .IN3(n28626), .IN4(n26267), .Q(
        n26158) );
  OA22X1 U29979 ( .IN1(n28632), .IN2(n26270), .IN3(n28625), .IN4(n26261), .Q(
        n26157) );
  OA22X1 U29980 ( .IN1(n28627), .IN2(n26269), .IN3(n28631), .IN4(n26271), .Q(
        n26156) );
  OA22X1 U29981 ( .IN1(n28630), .IN2(n26268), .IN3(n28629), .IN4(n26258), .Q(
        n26155) );
  NAND4X0 U29982 ( .IN1(n26158), .IN2(n26157), .IN3(n26156), .IN4(n26155), 
        .QN(s7_addr_o[5]) );
  OA22X1 U29983 ( .IN1(n26267), .IN2(n28643), .IN3(n26227), .IN4(n28638), .Q(
        n26162) );
  OA22X1 U29984 ( .IN1(n26259), .IN2(n28637), .IN3(n26273), .IN4(n28639), .Q(
        n26161) );
  OA22X1 U29985 ( .IN1(n26268), .IN2(n28640), .IN3(n26270), .IN4(n28644), .Q(
        n26160) );
  OA22X1 U29986 ( .IN1(n26258), .IN2(n28642), .IN3(n26260), .IN4(n28641), .Q(
        n26159) );
  NAND4X0 U29987 ( .IN1(n26162), .IN2(n26161), .IN3(n26160), .IN4(n26159), 
        .QN(s7_addr_o[6]) );
  OA22X1 U29988 ( .IN1(n26272), .IN2(n28654), .IN3(n26273), .IN4(n28655), .Q(
        n26166) );
  OA22X1 U29989 ( .IN1(n26268), .IN2(n28652), .IN3(n26269), .IN4(n28649), .Q(
        n26165) );
  OA22X1 U29990 ( .IN1(n26253), .IN2(n28653), .IN3(n26274), .IN4(n28651), .Q(
        n26164) );
  OA22X1 U29991 ( .IN1(n26262), .IN2(n28656), .IN3(n26271), .IN4(n28650), .Q(
        n26163) );
  NAND4X0 U29992 ( .IN1(n26166), .IN2(n26165), .IN3(n26164), .IN4(n26163), 
        .QN(s7_addr_o[7]) );
  OA22X1 U29993 ( .IN1(n26259), .IN2(n28662), .IN3(n26274), .IN4(n28661), .Q(
        n26170) );
  OA22X1 U29994 ( .IN1(n26262), .IN2(n28666), .IN3(n26273), .IN4(n28667), .Q(
        n26169) );
  OA22X1 U29995 ( .IN1(n26272), .IN2(n28664), .IN3(n26253), .IN4(n28665), .Q(
        n26168) );
  OA22X1 U29996 ( .IN1(n26236), .IN2(n28663), .IN3(n26271), .IN4(n28668), .Q(
        n26167) );
  NAND4X0 U29997 ( .IN1(n26170), .IN2(n26169), .IN3(n26168), .IN4(n26167), 
        .QN(s7_addr_o[8]) );
  OA22X1 U29998 ( .IN1(n26271), .IN2(n28673), .IN3(n26269), .IN4(n28678), .Q(
        n26174) );
  OA22X1 U29999 ( .IN1(n26258), .IN2(n28680), .IN3(n26253), .IN4(n28676), .Q(
        n26173) );
  OA22X1 U30000 ( .IN1(n26262), .IN2(n28674), .IN3(n26260), .IN4(n28675), .Q(
        n26172) );
  OA22X1 U30001 ( .IN1(n26268), .IN2(n28679), .IN3(n26273), .IN4(n28677), .Q(
        n26171) );
  NAND4X0 U30002 ( .IN1(n26174), .IN2(n26173), .IN3(n26172), .IN4(n26171), 
        .QN(s7_addr_o[9]) );
  OA22X1 U30003 ( .IN1(n26258), .IN2(n28692), .IN3(n26267), .IN4(n28687), .Q(
        n26178) );
  OA22X1 U30004 ( .IN1(n26262), .IN2(n28688), .IN3(n26274), .IN4(n28690), .Q(
        n26177) );
  OA22X1 U30005 ( .IN1(n26236), .IN2(n28686), .IN3(n26227), .IN4(n28685), .Q(
        n26176) );
  OA22X1 U30006 ( .IN1(n26259), .IN2(n28691), .IN3(n26273), .IN4(n28689), .Q(
        n26175) );
  NAND4X0 U30007 ( .IN1(n26178), .IN2(n26177), .IN3(n26176), .IN4(n26175), 
        .QN(s7_addr_o[10]) );
  OA22X1 U30008 ( .IN1(n26262), .IN2(n28697), .IN3(n26271), .IN4(n28701), .Q(
        n26182) );
  OA22X1 U30009 ( .IN1(n26267), .IN2(n28704), .IN3(n26274), .IN4(n28700), .Q(
        n26181) );
  OA22X1 U30010 ( .IN1(n26258), .IN2(n28702), .IN3(n26259), .IN4(n28703), .Q(
        n26180) );
  OA22X1 U30011 ( .IN1(n26236), .IN2(n28698), .IN3(n26273), .IN4(n28699), .Q(
        n26179) );
  NAND4X0 U30012 ( .IN1(n26182), .IN2(n26181), .IN3(n26180), .IN4(n26179), 
        .QN(s7_addr_o[11]) );
  OA22X1 U30013 ( .IN1(n26268), .IN2(n28710), .IN3(n26260), .IN4(n28711), .Q(
        n26186) );
  OA22X1 U30014 ( .IN1(n26267), .IN2(n28716), .IN3(n26259), .IN4(n28715), .Q(
        n26185) );
  OA22X1 U30015 ( .IN1(n26271), .IN2(n28709), .IN3(n26273), .IN4(n28713), .Q(
        n26184) );
  OA22X1 U30016 ( .IN1(n26272), .IN2(n28714), .IN3(n26270), .IN4(n28712), .Q(
        n26183) );
  NAND4X0 U30017 ( .IN1(n26186), .IN2(n26185), .IN3(n26184), .IN4(n26183), 
        .QN(s7_addr_o[12]) );
  OA22X1 U30018 ( .IN1(n26268), .IN2(n28728), .IN3(n26270), .IN4(n28726), .Q(
        n26190) );
  OA22X1 U30019 ( .IN1(n26272), .IN2(n28722), .IN3(n26227), .IN4(n28723), .Q(
        n26189) );
  OA22X1 U30020 ( .IN1(n26269), .IN2(n28721), .IN3(n26273), .IN4(n28727), .Q(
        n26188) );
  OA22X1 U30021 ( .IN1(n26267), .IN2(n28724), .IN3(n26274), .IN4(n28725), .Q(
        n26187) );
  NAND4X0 U30022 ( .IN1(n26190), .IN2(n26189), .IN3(n26188), .IN4(n26187), 
        .QN(s7_addr_o[13]) );
  OA22X1 U30023 ( .IN1(n26258), .IN2(n28734), .IN3(n26269), .IN4(n28737), .Q(
        n26194) );
  OA22X1 U30024 ( .IN1(n26271), .IN2(n28740), .IN3(n26273), .IN4(n28739), .Q(
        n26193) );
  OA22X1 U30025 ( .IN1(n26267), .IN2(n28735), .IN3(n26260), .IN4(n28733), .Q(
        n26192) );
  OA22X1 U30026 ( .IN1(n26236), .IN2(n28738), .IN3(n26270), .IN4(n28736), .Q(
        n26191) );
  NAND4X0 U30027 ( .IN1(n26194), .IN2(n26193), .IN3(n26192), .IN4(n26191), 
        .QN(s7_addr_o[14]) );
  OA22X1 U30028 ( .IN1(n26262), .IN2(n28750), .IN3(n26227), .IN4(n28747), .Q(
        n26198) );
  OA22X1 U30029 ( .IN1(n26259), .IN2(n28751), .IN3(n26273), .IN4(n28745), .Q(
        n26197) );
  OA22X1 U30030 ( .IN1(n26258), .IN2(n28746), .IN3(n26267), .IN4(n28752), .Q(
        n26196) );
  OA22X1 U30031 ( .IN1(n26236), .IN2(n28748), .IN3(n26260), .IN4(n28749), .Q(
        n26195) );
  NAND4X0 U30032 ( .IN1(n26198), .IN2(n26197), .IN3(n26196), .IN4(n26195), 
        .QN(s7_addr_o[15]) );
  OA22X1 U30033 ( .IN1(n26269), .IN2(n28757), .IN3(n26274), .IN4(n28764), .Q(
        n26202) );
  OA22X1 U30034 ( .IN1(n26262), .IN2(n28760), .IN3(n26271), .IN4(n28759), .Q(
        n26201) );
  OA22X1 U30035 ( .IN1(n26258), .IN2(n28758), .IN3(n26236), .IN4(n28762), .Q(
        n26200) );
  OA22X1 U30036 ( .IN1(n26267), .IN2(n28761), .IN3(n26261), .IN4(n28763), .Q(
        n26199) );
  NAND4X0 U30037 ( .IN1(n26202), .IN2(n26201), .IN3(n26200), .IN4(n26199), 
        .QN(s7_addr_o[16]) );
  OA22X1 U30038 ( .IN1(n26262), .IN2(n28774), .IN3(n26273), .IN4(n28769), .Q(
        n26206) );
  OA22X1 U30039 ( .IN1(n26268), .IN2(n28776), .IN3(n26260), .IN4(n28770), .Q(
        n26205) );
  OA22X1 U30040 ( .IN1(n26267), .IN2(n28773), .IN3(n26259), .IN4(n28771), .Q(
        n26204) );
  OA22X1 U30041 ( .IN1(n26258), .IN2(n28772), .IN3(n26271), .IN4(n28775), .Q(
        n26203) );
  NAND4X0 U30042 ( .IN1(n26206), .IN2(n26205), .IN3(n26204), .IN4(n26203), 
        .QN(s7_addr_o[17]) );
  OA22X1 U30043 ( .IN1(n26272), .IN2(n28786), .IN3(n26270), .IN4(n28787), .Q(
        n26210) );
  OA22X1 U30044 ( .IN1(n26271), .IN2(n28784), .IN3(n26274), .IN4(n28785), .Q(
        n26209) );
  OA22X1 U30045 ( .IN1(n26236), .IN2(n28788), .IN3(n26261), .IN4(n28781), .Q(
        n26208) );
  OA22X1 U30046 ( .IN1(n26267), .IN2(n28782), .IN3(n26269), .IN4(n28783), .Q(
        n26207) );
  NAND4X0 U30047 ( .IN1(n26210), .IN2(n26209), .IN3(n26208), .IN4(n26207), 
        .QN(s7_addr_o[18]) );
  OA22X1 U30048 ( .IN1(n26258), .IN2(n28796), .IN3(n26253), .IN4(n28794), .Q(
        n26214) );
  OA22X1 U30049 ( .IN1(n26268), .IN2(n28800), .IN3(n26269), .IN4(n28795), .Q(
        n26213) );
  OA22X1 U30050 ( .IN1(n26262), .IN2(n28798), .IN3(n26274), .IN4(n28793), .Q(
        n26212) );
  OA22X1 U30051 ( .IN1(n26271), .IN2(n28797), .IN3(n26273), .IN4(n28799), .Q(
        n26211) );
  NAND4X0 U30052 ( .IN1(n26214), .IN2(n26213), .IN3(n26212), .IN4(n26211), 
        .QN(s7_addr_o[19]) );
  OA22X1 U30053 ( .IN1(n26272), .IN2(n28812), .IN3(n26261), .IN4(n28805), .Q(
        n26218) );
  OA22X1 U30054 ( .IN1(n26236), .IN2(n28808), .IN3(n26259), .IN4(n28811), .Q(
        n26217) );
  OA22X1 U30055 ( .IN1(n26262), .IN2(n28807), .IN3(n26227), .IN4(n28806), .Q(
        n26216) );
  OA22X1 U30056 ( .IN1(n26267), .IN2(n28810), .IN3(n26260), .IN4(n28809), .Q(
        n26215) );
  NAND4X0 U30057 ( .IN1(n26218), .IN2(n26217), .IN3(n26216), .IN4(n26215), 
        .QN(s7_addr_o[20]) );
  OA22X1 U30058 ( .IN1(n26258), .IN2(n28822), .IN3(n26260), .IN4(n28818), .Q(
        n26222) );
  OA22X1 U30059 ( .IN1(n26227), .IN2(n28821), .IN3(n26273), .IN4(n28817), .Q(
        n26221) );
  OA22X1 U30060 ( .IN1(n26268), .IN2(n28824), .IN3(n26267), .IN4(n28819), .Q(
        n26220) );
  OA22X1 U30061 ( .IN1(n26270), .IN2(n28820), .IN3(n26259), .IN4(n28823), .Q(
        n26219) );
  NAND4X0 U30062 ( .IN1(n26222), .IN2(n26221), .IN3(n26220), .IN4(n26219), 
        .QN(s7_addr_o[21]) );
  OA22X1 U30063 ( .IN1(n26272), .IN2(n28833), .IN3(n26270), .IN4(n28831), .Q(
        n26226) );
  OA22X1 U30064 ( .IN1(n26259), .IN2(n28834), .IN3(n26261), .IN4(n28829), .Q(
        n26225) );
  OA22X1 U30065 ( .IN1(n26268), .IN2(n28832), .IN3(n26274), .IN4(n28837), .Q(
        n26224) );
  OA22X1 U30066 ( .IN1(n26267), .IN2(n28838), .IN3(n26271), .IN4(n28836), .Q(
        n26223) );
  NAND4X0 U30067 ( .IN1(n26226), .IN2(n26225), .IN3(n26224), .IN4(n26223), 
        .QN(s7_addr_o[22]) );
  OA22X1 U30068 ( .IN1(n26267), .IN2(n28850), .IN3(n26227), .IN4(n28852), .Q(
        n26231) );
  OA22X1 U30069 ( .IN1(n26268), .IN2(n28845), .IN3(n26270), .IN4(n28843), .Q(
        n26230) );
  OA22X1 U30070 ( .IN1(n26260), .IN2(n28846), .IN3(n26273), .IN4(n28851), .Q(
        n26229) );
  OA22X1 U30071 ( .IN1(n26258), .IN2(n28848), .IN3(n26269), .IN4(n28849), .Q(
        n26228) );
  NAND4X0 U30072 ( .IN1(n26231), .IN2(n26230), .IN3(n26229), .IN4(n26228), 
        .QN(s7_addr_o[23]) );
  OA22X1 U30073 ( .IN1(n28858), .IN2(n26262), .IN3(n28860), .IN4(n26273), .Q(
        n26235) );
  OA22X1 U30074 ( .IN1(n28859), .IN2(n26259), .IN3(n28861), .IN4(n26271), .Q(
        n26234) );
  OA22X1 U30075 ( .IN1(n28864), .IN2(n26268), .IN3(n28857), .IN4(n26253), .Q(
        n26233) );
  OA22X1 U30076 ( .IN1(n28865), .IN2(n26274), .IN3(n28863), .IN4(n26258), .Q(
        n26232) );
  NAND4X0 U30077 ( .IN1(n26235), .IN2(n26234), .IN3(n26233), .IN4(n26232), 
        .QN(s7_addr_o[24]) );
  OA22X1 U30078 ( .IN1(n28873), .IN2(n26270), .IN3(n28877), .IN4(n26236), .Q(
        n26240) );
  OA22X1 U30079 ( .IN1(n28870), .IN2(n26258), .IN3(n28874), .IN4(n26253), .Q(
        n26239) );
  OA22X1 U30080 ( .IN1(n28871), .IN2(n26260), .IN3(n28872), .IN4(n26271), .Q(
        n26238) );
  OA22X1 U30081 ( .IN1(n28875), .IN2(n26261), .IN3(n28876), .IN4(n26259), .Q(
        n26237) );
  NAND4X0 U30082 ( .IN1(n26240), .IN2(n26239), .IN3(n26238), .IN4(n26237), 
        .QN(s7_addr_o[25]) );
  OA22X1 U30083 ( .IN1(n28887), .IN2(n26268), .IN3(n28886), .IN4(n26271), .Q(
        n26244) );
  OA22X1 U30084 ( .IN1(n28889), .IN2(n26273), .IN3(n28888), .IN4(n26269), .Q(
        n26243) );
  OA22X1 U30085 ( .IN1(n28885), .IN2(n26262), .IN3(n28883), .IN4(n26274), .Q(
        n26242) );
  OA22X1 U30086 ( .IN1(n28884), .IN2(n26272), .IN3(n28882), .IN4(n26267), .Q(
        n26241) );
  NAND4X0 U30087 ( .IN1(n26244), .IN2(n26243), .IN3(n26242), .IN4(n26241), 
        .QN(s7_addr_o[26]) );
  OA22X1 U30088 ( .IN1(n28897), .IN2(n26274), .IN3(n28900), .IN4(n26271), .Q(
        n26248) );
  OA22X1 U30089 ( .IN1(n28895), .IN2(n26268), .IN3(n28901), .IN4(n26253), .Q(
        n26247) );
  OA22X1 U30090 ( .IN1(n28899), .IN2(n26270), .IN3(n28898), .IN4(n26261), .Q(
        n26246) );
  OA22X1 U30091 ( .IN1(n28896), .IN2(n26269), .IN3(n28894), .IN4(n26258), .Q(
        n26245) );
  NAND4X0 U30092 ( .IN1(n26248), .IN2(n26247), .IN3(n26246), .IN4(n26245), 
        .QN(s7_addr_o[27]) );
  OA22X1 U30093 ( .IN1(n28907), .IN2(n26260), .IN3(n28913), .IN4(n26273), .Q(
        n26252) );
  OA22X1 U30094 ( .IN1(n28912), .IN2(n26258), .IN3(n28908), .IN4(n26253), .Q(
        n26251) );
  OA22X1 U30095 ( .IN1(n28911), .IN2(n26268), .IN3(n28906), .IN4(n26271), .Q(
        n26250) );
  OA22X1 U30096 ( .IN1(n28909), .IN2(n26262), .IN3(n28910), .IN4(n26259), .Q(
        n26249) );
  NAND4X0 U30097 ( .IN1(n26252), .IN2(n26251), .IN3(n26250), .IN4(n26249), 
        .QN(s7_addr_o[28]) );
  OA22X1 U30098 ( .IN1(n28926), .IN2(n26270), .IN3(n28920), .IN4(n26259), .Q(
        n26257) );
  OA22X1 U30099 ( .IN1(n28921), .IN2(n26261), .IN3(n28923), .IN4(n26271), .Q(
        n26256) );
  OA22X1 U30100 ( .IN1(n28924), .IN2(n26268), .IN3(n28925), .IN4(n26258), .Q(
        n26255) );
  OA22X1 U30101 ( .IN1(n28922), .IN2(n26274), .IN3(n28919), .IN4(n26253), .Q(
        n26254) );
  NAND4X0 U30102 ( .IN1(n26257), .IN2(n26256), .IN3(n26255), .IN4(n26254), 
        .QN(s7_addr_o[29]) );
  OA22X1 U30103 ( .IN1(n28936), .IN2(n26259), .IN3(n28931), .IN4(n26258), .Q(
        n26266) );
  OA22X1 U30104 ( .IN1(n28937), .IN2(n26260), .IN3(n28940), .IN4(n26267), .Q(
        n26265) );
  OA22X1 U30105 ( .IN1(n28935), .IN2(n26268), .IN3(n28933), .IN4(n26261), .Q(
        n26264) );
  OA22X1 U30106 ( .IN1(n28932), .IN2(n26262), .IN3(n28939), .IN4(n26271), .Q(
        n26263) );
  NAND4X0 U30107 ( .IN1(n26266), .IN2(n26265), .IN3(n26264), .IN4(n26263), 
        .QN(s7_addr_o[30]) );
  OA22X1 U30108 ( .IN1(n28952), .IN2(n26268), .IN3(n28958), .IN4(n26267), .Q(
        n26278) );
  OA22X1 U30109 ( .IN1(n28948), .IN2(n26270), .IN3(n28954), .IN4(n26269), .Q(
        n26277) );
  OA22X1 U30110 ( .IN1(n28950), .IN2(n26272), .IN3(n28946), .IN4(n26271), .Q(
        n26276) );
  OA22X1 U30111 ( .IN1(n28956), .IN2(n26274), .IN3(n28960), .IN4(n26273), .Q(
        n26275) );
  NAND4X0 U30112 ( .IN1(n26278), .IN2(n26277), .IN3(n26276), .IN4(n26275), 
        .QN(s7_addr_o[31]) );
  OA22X1 U30113 ( .IN1(n29254), .IN2(n26280), .IN3(n29292), .IN4(n26279), .Q(
        n26290) );
  OA22X1 U30114 ( .IN1(n29273), .IN2(n26282), .IN3(n29235), .IN4(n26281), .Q(
        n26289) );
  OA22X1 U30115 ( .IN1(n29349), .IN2(n26284), .IN3(n29311), .IN4(n26283), .Q(
        n26288) );
  OA22X1 U30116 ( .IN1(n29368), .IN2(n26286), .IN3(n29330), .IN4(n26285), .Q(
        n26287) );
  NAND4X0 U30117 ( .IN1(n26290), .IN2(n26289), .IN3(n26288), .IN4(n26287), 
        .QN(s6_stb_o) );
  INVX0 U30118 ( .INP(n29082), .ZN(n26576) );
  INVX0 U30119 ( .INP(n26527), .ZN(n29075) );
  INVX0 U30120 ( .INP(n29075), .ZN(n26577) );
  OA22X1 U30121 ( .IN1(n26576), .IN2(n28123), .IN3(n26577), .IN4(n28121), .Q(
        n26294) );
  INVX0 U30122 ( .INP(n29084), .ZN(n26558) );
  OA22X1 U30123 ( .IN1(n26558), .IN2(n28125), .IN3(n26541), .IN4(n28127), .Q(
        n26293) );
  INVX0 U30124 ( .INP(n29081), .ZN(n26575) );
  INVX0 U30125 ( .INP(n29073), .ZN(n26565) );
  OA22X1 U30126 ( .IN1(n26575), .IN2(n28124), .IN3(n26565), .IN4(n28126), .Q(
        n26292) );
  INVX0 U30127 ( .INP(n29083), .ZN(n26573) );
  OA22X1 U30128 ( .IN1(n26560), .IN2(n28128), .IN3(n26573), .IN4(n28122), .Q(
        n26291) );
  NAND4X0 U30129 ( .IN1(n26294), .IN2(n26293), .IN3(n26292), .IN4(n26291), 
        .QN(s6_we_o) );
  INVX0 U30130 ( .INP(n29084), .ZN(n26571) );
  OA22X1 U30131 ( .IN1(n26560), .IN2(n28140), .IN3(n26571), .IN4(n28136), .Q(
        n26298) );
  OA22X1 U30132 ( .IN1(n26541), .IN2(n28137), .IN3(n26527), .IN4(n28135), .Q(
        n26297) );
  INVX0 U30133 ( .INP(n29082), .ZN(n26532) );
  OA22X1 U30134 ( .IN1(n26575), .IN2(n28134), .IN3(n26532), .IN4(n28133), .Q(
        n26296) );
  OA22X1 U30135 ( .IN1(n26565), .IN2(n28139), .IN3(n26573), .IN4(n28138), .Q(
        n26295) );
  NAND4X0 U30136 ( .IN1(n26298), .IN2(n26297), .IN3(n26296), .IN4(n26295), 
        .QN(s6_data_o[0]) );
  INVX0 U30137 ( .INP(n29083), .ZN(n26566) );
  OA22X1 U30138 ( .IN1(n26566), .IN2(n28149), .IN3(n26571), .IN4(n28152), .Q(
        n26302) );
  OA22X1 U30139 ( .IN1(n26575), .IN2(n28150), .IN3(n26560), .IN4(n28146), .Q(
        n26301) );
  INVX0 U30140 ( .INP(n29073), .ZN(n26574) );
  OA22X1 U30141 ( .IN1(n26574), .IN2(n28145), .IN3(n26527), .IN4(n28147), .Q(
        n26300) );
  OA22X1 U30142 ( .IN1(n26532), .IN2(n28148), .IN3(n26541), .IN4(n28151), .Q(
        n26299) );
  NAND4X0 U30143 ( .IN1(n26302), .IN2(n26301), .IN3(n26300), .IN4(n26299), 
        .QN(s6_data_o[1]) );
  OA22X1 U30144 ( .IN1(n26575), .IN2(n28160), .IN3(n26571), .IN4(n28162), .Q(
        n26306) );
  OA22X1 U30145 ( .IN1(n26576), .IN2(n28163), .IN3(n26541), .IN4(n28157), .Q(
        n26305) );
  INVX0 U30146 ( .INP(n29076), .ZN(n26572) );
  OA22X1 U30147 ( .IN1(n26572), .IN2(n28164), .IN3(n26527), .IN4(n28161), .Q(
        n26304) );
  OA22X1 U30148 ( .IN1(n26565), .IN2(n28159), .IN3(n26573), .IN4(n28158), .Q(
        n26303) );
  NAND4X0 U30149 ( .IN1(n26306), .IN2(n26305), .IN3(n26304), .IN4(n26303), 
        .QN(s6_data_o[2]) );
  OA22X1 U30150 ( .IN1(n26576), .IN2(n28176), .IN3(n26573), .IN4(n28171), .Q(
        n26310) );
  OA22X1 U30151 ( .IN1(n26559), .IN2(n28172), .IN3(n26541), .IN4(n28169), .Q(
        n26309) );
  OA22X1 U30152 ( .IN1(n26560), .IN2(n28174), .IN3(n26571), .IN4(n28175), .Q(
        n26308) );
  OA22X1 U30153 ( .IN1(n26574), .IN2(n28170), .IN3(n26527), .IN4(n28173), .Q(
        n26307) );
  NAND4X0 U30154 ( .IN1(n26310), .IN2(n26309), .IN3(n26308), .IN4(n26307), 
        .QN(s6_data_o[3]) );
  OA22X1 U30155 ( .IN1(n26576), .IN2(n28186), .IN3(n26571), .IN4(n28183), .Q(
        n26314) );
  OA22X1 U30156 ( .IN1(n26575), .IN2(n28182), .IN3(n26574), .IN4(n28188), .Q(
        n26313) );
  OA22X1 U30157 ( .IN1(n26560), .IN2(n28184), .IN3(n26527), .IN4(n28181), .Q(
        n26312) );
  OA22X1 U30158 ( .IN1(n26573), .IN2(n28185), .IN3(n26541), .IN4(n28187), .Q(
        n26311) );
  NAND4X0 U30159 ( .IN1(n26314), .IN2(n26313), .IN3(n26312), .IN4(n26311), 
        .QN(s6_data_o[4]) );
  OA22X1 U30160 ( .IN1(n26576), .IN2(n28194), .IN3(n26571), .IN4(n28197), .Q(
        n26318) );
  OA22X1 U30161 ( .IN1(n26559), .IN2(n28196), .IN3(n26560), .IN4(n28200), .Q(
        n26317) );
  OA22X1 U30162 ( .IN1(n26565), .IN2(n28193), .IN3(n26573), .IN4(n28198), .Q(
        n26316) );
  OA22X1 U30163 ( .IN1(n26541), .IN2(n28195), .IN3(n26527), .IN4(n28199), .Q(
        n26315) );
  NAND4X0 U30164 ( .IN1(n26318), .IN2(n26317), .IN3(n26316), .IN4(n26315), 
        .QN(s6_data_o[5]) );
  OA22X1 U30165 ( .IN1(n26532), .IN2(n28206), .IN3(n26571), .IN4(n28205), .Q(
        n26322) );
  OA22X1 U30166 ( .IN1(n26572), .IN2(n28207), .IN3(n26541), .IN4(n28210), .Q(
        n26321) );
  OA22X1 U30167 ( .IN1(n26565), .IN2(n28212), .IN3(n26573), .IN4(n28211), .Q(
        n26320) );
  OA22X1 U30168 ( .IN1(n26575), .IN2(n28208), .IN3(n26527), .IN4(n28209), .Q(
        n26319) );
  NAND4X0 U30169 ( .IN1(n26322), .IN2(n26321), .IN3(n26320), .IN4(n26319), 
        .QN(s6_data_o[6]) );
  OA22X1 U30170 ( .IN1(n26566), .IN2(n28217), .IN3(n26571), .IN4(n28223), .Q(
        n26326) );
  OA22X1 U30171 ( .IN1(n26559), .IN2(n28220), .IN3(n26574), .IN4(n28218), .Q(
        n26325) );
  OA22X1 U30172 ( .IN1(n26576), .IN2(n28224), .IN3(n26577), .IN4(n28221), .Q(
        n26324) );
  OA22X1 U30173 ( .IN1(n26560), .IN2(n28219), .IN3(n26541), .IN4(n28222), .Q(
        n26323) );
  NAND4X0 U30174 ( .IN1(n26326), .IN2(n26325), .IN3(n26324), .IN4(n26323), 
        .QN(s6_data_o[7]) );
  OA22X1 U30175 ( .IN1(n26532), .IN2(n28231), .IN3(n26577), .IN4(n28235), .Q(
        n26330) );
  OA22X1 U30176 ( .IN1(n26574), .IN2(n28234), .IN3(n26573), .IN4(n28236), .Q(
        n26329) );
  INVX0 U30177 ( .INP(n26541), .ZN(n29074) );
  INVX0 U30178 ( .INP(n29074), .ZN(n26578) );
  OA22X1 U30179 ( .IN1(n26571), .IN2(n28229), .IN3(n26578), .IN4(n28233), .Q(
        n26328) );
  OA22X1 U30180 ( .IN1(n26575), .IN2(n28230), .IN3(n26560), .IN4(n28232), .Q(
        n26327) );
  NAND4X0 U30181 ( .IN1(n26330), .IN2(n26329), .IN3(n26328), .IN4(n26327), 
        .QN(s6_data_o[8]) );
  OA22X1 U30182 ( .IN1(n26559), .IN2(n28242), .IN3(n26571), .IN4(n28245), .Q(
        n26334) );
  OA22X1 U30183 ( .IN1(n26576), .IN2(n28246), .IN3(n26577), .IN4(n28247), .Q(
        n26333) );
  OA22X1 U30184 ( .IN1(n26572), .IN2(n28244), .IN3(n26573), .IN4(n28241), .Q(
        n26332) );
  OA22X1 U30185 ( .IN1(n26565), .IN2(n28248), .IN3(n26578), .IN4(n28243), .Q(
        n26331) );
  NAND4X0 U30186 ( .IN1(n26334), .IN2(n26333), .IN3(n26332), .IN4(n26331), 
        .QN(s6_data_o[9]) );
  OA22X1 U30187 ( .IN1(n26560), .IN2(n28257), .IN3(n26574), .IN4(n28256), .Q(
        n26338) );
  OA22X1 U30188 ( .IN1(n26575), .IN2(n28258), .IN3(n26577), .IN4(n28259), .Q(
        n26337) );
  OA22X1 U30189 ( .IN1(n26573), .IN2(n28254), .IN3(n26541), .IN4(n28253), .Q(
        n26336) );
  OA22X1 U30190 ( .IN1(n26532), .IN2(n28260), .IN3(n26571), .IN4(n28255), .Q(
        n26335) );
  NAND4X0 U30191 ( .IN1(n26338), .IN2(n26337), .IN3(n26336), .IN4(n26335), 
        .QN(s6_data_o[10]) );
  OA22X1 U30192 ( .IN1(n26559), .IN2(n28266), .IN3(n26573), .IN4(n28268), .Q(
        n26342) );
  OA22X1 U30193 ( .IN1(n26576), .IN2(n28265), .IN3(n26571), .IN4(n28270), .Q(
        n26341) );
  OA22X1 U30194 ( .IN1(n26574), .IN2(n28271), .IN3(n26577), .IN4(n28269), .Q(
        n26340) );
  OA22X1 U30195 ( .IN1(n26572), .IN2(n28272), .IN3(n26541), .IN4(n28267), .Q(
        n26339) );
  NAND4X0 U30196 ( .IN1(n26342), .IN2(n26341), .IN3(n26340), .IN4(n26339), 
        .QN(s6_data_o[11]) );
  OA22X1 U30197 ( .IN1(n26532), .IN2(n28280), .IN3(n26571), .IN4(n28281), .Q(
        n26346) );
  OA22X1 U30198 ( .IN1(n26560), .IN2(n28278), .IN3(n26541), .IN4(n28279), .Q(
        n26345) );
  OA22X1 U30199 ( .IN1(n26565), .IN2(n28282), .IN3(n26577), .IN4(n28277), .Q(
        n26344) );
  OA22X1 U30200 ( .IN1(n26575), .IN2(n28284), .IN3(n26566), .IN4(n28283), .Q(
        n26343) );
  NAND4X0 U30201 ( .IN1(n26346), .IN2(n26345), .IN3(n26344), .IN4(n26343), 
        .QN(s6_data_o[12]) );
  OA22X1 U30202 ( .IN1(n26572), .IN2(n28294), .IN3(n26532), .IN4(n28296), .Q(
        n26350) );
  OA22X1 U30203 ( .IN1(n26566), .IN2(n28289), .IN3(n26541), .IN4(n28291), .Q(
        n26349) );
  OA22X1 U30204 ( .IN1(n26565), .IN2(n28292), .IN3(n26571), .IN4(n28293), .Q(
        n26348) );
  OA22X1 U30205 ( .IN1(n26559), .IN2(n28290), .IN3(n26577), .IN4(n28295), .Q(
        n26347) );
  NAND4X0 U30206 ( .IN1(n26350), .IN2(n26349), .IN3(n26348), .IN4(n26347), 
        .QN(s6_data_o[13]) );
  OA22X1 U30207 ( .IN1(n26576), .IN2(n28308), .IN3(n26574), .IN4(n28305), .Q(
        n26354) );
  OA22X1 U30208 ( .IN1(n26560), .IN2(n28304), .IN3(n26541), .IN4(n28301), .Q(
        n26353) );
  OA22X1 U30209 ( .IN1(n26573), .IN2(n28307), .IN3(n26577), .IN4(n28303), .Q(
        n26352) );
  OA22X1 U30210 ( .IN1(n26575), .IN2(n28306), .IN3(n26571), .IN4(n28302), .Q(
        n26351) );
  NAND4X0 U30211 ( .IN1(n26354), .IN2(n26353), .IN3(n26352), .IN4(n26351), 
        .QN(s6_data_o[14]) );
  OA22X1 U30212 ( .IN1(n26559), .IN2(n28316), .IN3(n26558), .IN4(n28318), .Q(
        n26358) );
  OA22X1 U30213 ( .IN1(n26572), .IN2(n28315), .IN3(n26541), .IN4(n28317), .Q(
        n26357) );
  OA22X1 U30214 ( .IN1(n26532), .IN2(n28314), .IN3(n26573), .IN4(n28320), .Q(
        n26356) );
  OA22X1 U30215 ( .IN1(n26565), .IN2(n28313), .IN3(n26577), .IN4(n28319), .Q(
        n26355) );
  NAND4X0 U30216 ( .IN1(n26358), .IN2(n26357), .IN3(n26356), .IN4(n26355), 
        .QN(s6_data_o[15]) );
  OA22X1 U30217 ( .IN1(n26558), .IN2(n28325), .IN3(n26541), .IN4(n28328), .Q(
        n26362) );
  OA22X1 U30218 ( .IN1(n26565), .IN2(n28326), .IN3(n26566), .IN4(n28329), .Q(
        n26361) );
  OA22X1 U30219 ( .IN1(n26560), .IN2(n28332), .IN3(n26532), .IN4(n28331), .Q(
        n26360) );
  OA22X1 U30220 ( .IN1(n26559), .IN2(n28330), .IN3(n26577), .IN4(n28327), .Q(
        n26359) );
  NAND4X0 U30221 ( .IN1(n26362), .IN2(n26361), .IN3(n26360), .IN4(n26359), 
        .QN(s6_data_o[16]) );
  OA22X1 U30222 ( .IN1(n26575), .IN2(n28340), .IN3(n26571), .IN4(n28339), .Q(
        n26366) );
  OA22X1 U30223 ( .IN1(n26541), .IN2(n28343), .IN3(n26577), .IN4(n28341), .Q(
        n26365) );
  OA22X1 U30224 ( .IN1(n26572), .IN2(n28344), .IN3(n26574), .IN4(n28338), .Q(
        n26364) );
  OA22X1 U30225 ( .IN1(n26532), .IN2(n28342), .IN3(n26566), .IN4(n28337), .Q(
        n26363) );
  NAND4X0 U30226 ( .IN1(n26366), .IN2(n26365), .IN3(n26364), .IN4(n26363), 
        .QN(s6_data_o[17]) );
  OA22X1 U30227 ( .IN1(n26576), .IN2(n28350), .IN3(n26574), .IN4(n28355), .Q(
        n26370) );
  OA22X1 U30228 ( .IN1(n26566), .IN2(n28354), .IN3(n26571), .IN4(n28349), .Q(
        n26369) );
  OA22X1 U30229 ( .IN1(n26560), .IN2(n28356), .IN3(n26577), .IN4(n28353), .Q(
        n26368) );
  OA22X1 U30230 ( .IN1(n26559), .IN2(n28352), .IN3(n26541), .IN4(n28351), .Q(
        n26367) );
  NAND4X0 U30231 ( .IN1(n26370), .IN2(n26369), .IN3(n26368), .IN4(n26367), 
        .QN(s6_data_o[18]) );
  OA22X1 U30232 ( .IN1(n26532), .IN2(n28362), .IN3(n26573), .IN4(n28365), .Q(
        n26374) );
  OA22X1 U30233 ( .IN1(n26565), .IN2(n28363), .IN3(n26571), .IN4(n28361), .Q(
        n26373) );
  OA22X1 U30234 ( .IN1(n26559), .IN2(n28366), .IN3(n26560), .IN4(n28364), .Q(
        n26372) );
  OA22X1 U30235 ( .IN1(n26541), .IN2(n28368), .IN3(n26577), .IN4(n28367), .Q(
        n26371) );
  NAND4X0 U30236 ( .IN1(n26374), .IN2(n26373), .IN3(n26372), .IN4(n26371), 
        .QN(s6_data_o[19]) );
  OA22X1 U30237 ( .IN1(n26572), .IN2(n28377), .IN3(n26532), .IN4(n28374), .Q(
        n26378) );
  OA22X1 U30238 ( .IN1(n26541), .IN2(n28379), .IN3(n26577), .IN4(n28375), .Q(
        n26377) );
  OA22X1 U30239 ( .IN1(n26559), .IN2(n28378), .IN3(n26573), .IN4(n28376), .Q(
        n26376) );
  OA22X1 U30240 ( .IN1(n26565), .IN2(n28373), .IN3(n26558), .IN4(n28380), .Q(
        n26375) );
  NAND4X0 U30241 ( .IN1(n26378), .IN2(n26377), .IN3(n26376), .IN4(n26375), 
        .QN(s6_data_o[20]) );
  OA22X1 U30242 ( .IN1(n26571), .IN2(n28385), .IN3(n26577), .IN4(n28391), .Q(
        n26382) );
  OA22X1 U30243 ( .IN1(n26566), .IN2(n28387), .IN3(n26541), .IN4(n28389), .Q(
        n26381) );
  OA22X1 U30244 ( .IN1(n26559), .IN2(n28392), .IN3(n26574), .IN4(n28388), .Q(
        n26380) );
  OA22X1 U30245 ( .IN1(n26572), .IN2(n28386), .IN3(n26532), .IN4(n28390), .Q(
        n26379) );
  NAND4X0 U30246 ( .IN1(n26382), .IN2(n26381), .IN3(n26380), .IN4(n26379), 
        .QN(s6_data_o[21]) );
  OA22X1 U30247 ( .IN1(n26572), .IN2(n28402), .IN3(n26574), .IN4(n28403), .Q(
        n26386) );
  OA22X1 U30248 ( .IN1(n26558), .IN2(n28399), .IN3(n26577), .IN4(n28397), .Q(
        n26385) );
  OA22X1 U30249 ( .IN1(n26559), .IN2(n28400), .IN3(n26541), .IN4(n28401), .Q(
        n26384) );
  OA22X1 U30250 ( .IN1(n26532), .IN2(n28404), .IN3(n26566), .IN4(n28398), .Q(
        n26383) );
  NAND4X0 U30251 ( .IN1(n26386), .IN2(n26385), .IN3(n26384), .IN4(n26383), 
        .QN(s6_data_o[22]) );
  OA22X1 U30252 ( .IN1(n26572), .IN2(n28415), .IN3(n26532), .IN4(n28414), .Q(
        n26390) );
  OA22X1 U30253 ( .IN1(n26565), .IN2(n28413), .IN3(n26541), .IN4(n28409), .Q(
        n26389) );
  OA22X1 U30254 ( .IN1(n26559), .IN2(n28416), .IN3(n26558), .IN4(n28412), .Q(
        n26388) );
  OA22X1 U30255 ( .IN1(n26566), .IN2(n28410), .IN3(n26527), .IN4(n28411), .Q(
        n26387) );
  NAND4X0 U30256 ( .IN1(n26390), .IN2(n26389), .IN3(n26388), .IN4(n26387), 
        .QN(s6_data_o[23]) );
  OA22X1 U30257 ( .IN1(n26576), .IN2(n28422), .IN3(n26541), .IN4(n28427), .Q(
        n26394) );
  OA22X1 U30258 ( .IN1(n26572), .IN2(n28424), .IN3(n26574), .IN4(n28421), .Q(
        n26393) );
  OA22X1 U30259 ( .IN1(n26566), .IN2(n28425), .IN3(n26571), .IN4(n28428), .Q(
        n26392) );
  OA22X1 U30260 ( .IN1(n26559), .IN2(n28426), .IN3(n26527), .IN4(n28423), .Q(
        n26391) );
  NAND4X0 U30261 ( .IN1(n26394), .IN2(n26393), .IN3(n26392), .IN4(n26391), 
        .QN(s6_data_o[24]) );
  OA22X1 U30262 ( .IN1(n26565), .IN2(n28439), .IN3(n26573), .IN4(n28433), .Q(
        n26398) );
  OA22X1 U30263 ( .IN1(n26572), .IN2(n28440), .IN3(n26532), .IN4(n28434), .Q(
        n26397) );
  OA22X1 U30264 ( .IN1(n26541), .IN2(n28436), .IN3(n26527), .IN4(n28435), .Q(
        n26396) );
  OA22X1 U30265 ( .IN1(n26559), .IN2(n28438), .IN3(n26558), .IN4(n28437), .Q(
        n26395) );
  NAND4X0 U30266 ( .IN1(n26398), .IN2(n26397), .IN3(n26396), .IN4(n26395), 
        .QN(s6_data_o[25]) );
  OA22X1 U30267 ( .IN1(n26565), .IN2(n28446), .IN3(n26527), .IN4(n28445), .Q(
        n26402) );
  OA22X1 U30268 ( .IN1(n26576), .IN2(n28450), .IN3(n26566), .IN4(n28449), .Q(
        n26401) );
  OA22X1 U30269 ( .IN1(n26558), .IN2(n28448), .IN3(n26541), .IN4(n28447), .Q(
        n26400) );
  OA22X1 U30270 ( .IN1(n26559), .IN2(n28452), .IN3(n26560), .IN4(n28451), .Q(
        n26399) );
  NAND4X0 U30271 ( .IN1(n26402), .IN2(n26401), .IN3(n26400), .IN4(n26399), 
        .QN(s6_data_o[26]) );
  OA22X1 U30272 ( .IN1(n26572), .IN2(n28461), .IN3(n26532), .IN4(n28464), .Q(
        n26406) );
  OA22X1 U30273 ( .IN1(n26559), .IN2(n28462), .IN3(n26574), .IN4(n28458), .Q(
        n26405) );
  OA22X1 U30274 ( .IN1(n26578), .IN2(n28460), .IN3(n26527), .IN4(n28459), .Q(
        n26404) );
  OA22X1 U30275 ( .IN1(n26566), .IN2(n28457), .IN3(n26571), .IN4(n28463), .Q(
        n26403) );
  NAND4X0 U30276 ( .IN1(n26406), .IN2(n26405), .IN3(n26404), .IN4(n26403), 
        .QN(s6_data_o[27]) );
  OA22X1 U30277 ( .IN1(n26572), .IN2(n28476), .IN3(n26574), .IN4(n28470), .Q(
        n26410) );
  OA22X1 U30278 ( .IN1(n26566), .IN2(n28471), .IN3(n26527), .IN4(n28473), .Q(
        n26409) );
  OA22X1 U30279 ( .IN1(n26559), .IN2(n28474), .IN3(n26558), .IN4(n28475), .Q(
        n26408) );
  OA22X1 U30280 ( .IN1(n26532), .IN2(n28472), .IN3(n26541), .IN4(n28469), .Q(
        n26407) );
  NAND4X0 U30281 ( .IN1(n26410), .IN2(n26409), .IN3(n26408), .IN4(n26407), 
        .QN(s6_data_o[28]) );
  OA22X1 U30282 ( .IN1(n26559), .IN2(n28484), .IN3(n26573), .IN4(n28487), .Q(
        n26414) );
  OA22X1 U30283 ( .IN1(n26565), .IN2(n28486), .IN3(n26571), .IN4(n28483), .Q(
        n26413) );
  OA22X1 U30284 ( .IN1(n26576), .IN2(n28488), .IN3(n26527), .IN4(n28481), .Q(
        n26412) );
  OA22X1 U30285 ( .IN1(n26572), .IN2(n28482), .IN3(n26541), .IN4(n28485), .Q(
        n26411) );
  NAND4X0 U30286 ( .IN1(n26414), .IN2(n26413), .IN3(n26412), .IN4(n26411), 
        .QN(s6_data_o[29]) );
  OA22X1 U30287 ( .IN1(n26572), .IN2(n28498), .IN3(n26532), .IN4(n28497), .Q(
        n26418) );
  OA22X1 U30288 ( .IN1(n26574), .IN2(n28496), .IN3(n26527), .IN4(n28499), .Q(
        n26417) );
  OA22X1 U30289 ( .IN1(n26559), .IN2(n28494), .IN3(n26573), .IN4(n28493), .Q(
        n26416) );
  OA22X1 U30290 ( .IN1(n26558), .IN2(n28495), .IN3(n26541), .IN4(n28500), .Q(
        n26415) );
  NAND4X0 U30291 ( .IN1(n26418), .IN2(n26417), .IN3(n26416), .IN4(n26415), 
        .QN(s6_data_o[30]) );
  OA22X1 U30292 ( .IN1(n26566), .IN2(n28512), .IN3(n26541), .IN4(n28511), .Q(
        n26422) );
  OA22X1 U30293 ( .IN1(n26572), .IN2(n28509), .IN3(n26527), .IN4(n28507), .Q(
        n26421) );
  OA22X1 U30294 ( .IN1(n26576), .IN2(n28506), .IN3(n26571), .IN4(n28508), .Q(
        n26420) );
  OA22X1 U30295 ( .IN1(n26575), .IN2(n28510), .IN3(n26574), .IN4(n28505), .Q(
        n26419) );
  NAND4X0 U30296 ( .IN1(n26422), .IN2(n26421), .IN3(n26420), .IN4(n26419), 
        .QN(s6_data_o[31]) );
  OA22X1 U30297 ( .IN1(n26574), .IN2(n28524), .IN3(n26541), .IN4(n28521), .Q(
        n26426) );
  OA22X1 U30298 ( .IN1(n26558), .IN2(n28520), .IN3(n26527), .IN4(n28519), .Q(
        n26425) );
  OA22X1 U30299 ( .IN1(n26575), .IN2(n28518), .IN3(n26573), .IN4(n28523), .Q(
        n26424) );
  OA22X1 U30300 ( .IN1(n26572), .IN2(n28517), .IN3(n26532), .IN4(n28522), .Q(
        n26423) );
  NAND4X0 U30301 ( .IN1(n26426), .IN2(n26425), .IN3(n26424), .IN4(n26423), 
        .QN(s6_sel_o[0]) );
  OA22X1 U30302 ( .IN1(n26574), .IN2(n28536), .IN3(n26527), .IN4(n28529), .Q(
        n26430) );
  OA22X1 U30303 ( .IN1(n26572), .IN2(n28532), .IN3(n26558), .IN4(n28533), .Q(
        n26429) );
  OA22X1 U30304 ( .IN1(n26575), .IN2(n28534), .IN3(n26532), .IN4(n28530), .Q(
        n26428) );
  OA22X1 U30305 ( .IN1(n26566), .IN2(n28535), .IN3(n26541), .IN4(n28531), .Q(
        n26427) );
  NAND4X0 U30306 ( .IN1(n26430), .IN2(n26429), .IN3(n26428), .IN4(n26427), 
        .QN(s6_sel_o[1]) );
  OA22X1 U30307 ( .IN1(n26574), .IN2(n28548), .IN3(n26541), .IN4(n28545), .Q(
        n26434) );
  OA22X1 U30308 ( .IN1(n26572), .IN2(n28546), .IN3(n26532), .IN4(n28543), .Q(
        n26433) );
  OA22X1 U30309 ( .IN1(n26558), .IN2(n28542), .IN3(n26527), .IN4(n28541), .Q(
        n26432) );
  OA22X1 U30310 ( .IN1(n26575), .IN2(n28544), .IN3(n26566), .IN4(n28547), .Q(
        n26431) );
  NAND4X0 U30311 ( .IN1(n26434), .IN2(n26433), .IN3(n26432), .IN4(n26431), 
        .QN(s6_sel_o[2]) );
  OA22X1 U30312 ( .IN1(n26560), .IN2(n28554), .IN3(n26566), .IN4(n28556), .Q(
        n26438) );
  OA22X1 U30313 ( .IN1(n26532), .IN2(n28553), .IN3(n26574), .IN4(n28557), .Q(
        n26437) );
  OA22X1 U30314 ( .IN1(n26575), .IN2(n28558), .IN3(n26541), .IN4(n28559), .Q(
        n26436) );
  OA22X1 U30315 ( .IN1(n26558), .IN2(n28560), .IN3(n26527), .IN4(n28555), .Q(
        n26435) );
  NAND4X0 U30316 ( .IN1(n26438), .IN2(n26437), .IN3(n26436), .IN4(n26435), 
        .QN(s6_sel_o[3]) );
  OA22X1 U30317 ( .IN1(n26560), .IN2(n28570), .IN3(n26573), .IN4(n28568), .Q(
        n26442) );
  OA22X1 U30318 ( .IN1(n26559), .IN2(n28572), .IN3(n26565), .IN4(n28566), .Q(
        n26441) );
  OA22X1 U30319 ( .IN1(n26532), .IN2(n28571), .IN3(n26558), .IN4(n28567), .Q(
        n26440) );
  OA22X1 U30320 ( .IN1(n26578), .IN2(n28565), .IN3(n26527), .IN4(n28569), .Q(
        n26439) );
  NAND4X0 U30321 ( .IN1(n26442), .IN2(n26441), .IN3(n26440), .IN4(n26439), 
        .QN(s6_addr_o[0]) );
  OA22X1 U30322 ( .IN1(n26575), .IN2(n28580), .IN3(n26571), .IN4(n28584), .Q(
        n26446) );
  OA22X1 U30323 ( .IN1(n26576), .IN2(n28582), .IN3(n26573), .IN4(n28579), .Q(
        n26445) );
  OA22X1 U30324 ( .IN1(n26560), .IN2(n28578), .IN3(n26541), .IN4(n28577), .Q(
        n26444) );
  OA22X1 U30325 ( .IN1(n26565), .IN2(n28581), .IN3(n26527), .IN4(n28583), .Q(
        n26443) );
  NAND4X0 U30326 ( .IN1(n26446), .IN2(n26445), .IN3(n26444), .IN4(n26443), 
        .QN(s6_addr_o[1]) );
  OA22X1 U30327 ( .IN1(n28596), .IN2(n26577), .IN3(n28595), .IN4(n26541), .Q(
        n26450) );
  OA22X1 U30328 ( .IN1(n28590), .IN2(n26573), .IN3(n28589), .IN4(n26560), .Q(
        n26449) );
  OA22X1 U30329 ( .IN1(n28592), .IN2(n26574), .IN3(n28591), .IN4(n26575), .Q(
        n26448) );
  OA22X1 U30330 ( .IN1(n28594), .IN2(n26576), .IN3(n28593), .IN4(n26571), .Q(
        n26447) );
  NAND4X0 U30331 ( .IN1(n26450), .IN2(n26449), .IN3(n26448), .IN4(n26447), 
        .QN(s6_addr_o[2]) );
  OA22X1 U30332 ( .IN1(n28604), .IN2(n26576), .IN3(n28606), .IN4(n26573), .Q(
        n26454) );
  OA22X1 U30333 ( .IN1(n28602), .IN2(n26571), .IN3(n28603), .IN4(n26541), .Q(
        n26453) );
  OA22X1 U30334 ( .IN1(n28608), .IN2(n26577), .IN3(n28607), .IN4(n26565), .Q(
        n26452) );
  OA22X1 U30335 ( .IN1(n28605), .IN2(n26560), .IN3(n28601), .IN4(n26575), .Q(
        n26451) );
  NAND4X0 U30336 ( .IN1(n26454), .IN2(n26453), .IN3(n26452), .IN4(n26451), 
        .QN(s6_addr_o[3]) );
  OA22X1 U30337 ( .IN1(n28620), .IN2(n26578), .IN3(n28614), .IN4(n26558), .Q(
        n26458) );
  OA22X1 U30338 ( .IN1(n28617), .IN2(n26575), .IN3(n28613), .IN4(n26532), .Q(
        n26457) );
  OA22X1 U30339 ( .IN1(n28618), .IN2(n26565), .IN3(n28615), .IN4(n26573), .Q(
        n26456) );
  OA22X1 U30340 ( .IN1(n28616), .IN2(n26572), .IN3(n28619), .IN4(n26577), .Q(
        n26455) );
  NAND4X0 U30341 ( .IN1(n26458), .IN2(n26457), .IN3(n26456), .IN4(n26455), 
        .QN(s6_addr_o[4]) );
  OA22X1 U30342 ( .IN1(n28632), .IN2(n26576), .IN3(n28631), .IN4(n26573), .Q(
        n26462) );
  OA22X1 U30343 ( .IN1(n28630), .IN2(n26572), .IN3(n28629), .IN4(n26575), .Q(
        n26461) );
  OA22X1 U30344 ( .IN1(n28628), .IN2(n26578), .IN3(n28627), .IN4(n26558), .Q(
        n26460) );
  OA22X1 U30345 ( .IN1(n28626), .IN2(n26574), .IN3(n28625), .IN4(n26577), .Q(
        n26459) );
  NAND4X0 U30346 ( .IN1(n26462), .IN2(n26461), .IN3(n26460), .IN4(n26459), 
        .QN(s6_addr_o[5]) );
  OA22X1 U30347 ( .IN1(n26560), .IN2(n28640), .IN3(n26527), .IN4(n28639), .Q(
        n26466) );
  OA22X1 U30348 ( .IN1(n26532), .IN2(n28644), .IN3(n26565), .IN4(n28643), .Q(
        n26465) );
  OA22X1 U30349 ( .IN1(n26559), .IN2(n28642), .IN3(n26566), .IN4(n28638), .Q(
        n26464) );
  OA22X1 U30350 ( .IN1(n26558), .IN2(n28637), .IN3(n26578), .IN4(n28641), .Q(
        n26463) );
  NAND4X0 U30351 ( .IN1(n26466), .IN2(n26465), .IN3(n26464), .IN4(n26463), 
        .QN(s6_addr_o[6]) );
  OA22X1 U30352 ( .IN1(n26575), .IN2(n28654), .IN3(n26578), .IN4(n28651), .Q(
        n26470) );
  OA22X1 U30353 ( .IN1(n26558), .IN2(n28649), .IN3(n26527), .IN4(n28655), .Q(
        n26469) );
  OA22X1 U30354 ( .IN1(n26560), .IN2(n28652), .IN3(n26532), .IN4(n28656), .Q(
        n26468) );
  OA22X1 U30355 ( .IN1(n26565), .IN2(n28653), .IN3(n26566), .IN4(n28650), .Q(
        n26467) );
  NAND4X0 U30356 ( .IN1(n26470), .IN2(n26469), .IN3(n26468), .IN4(n26467), 
        .QN(s6_addr_o[7]) );
  OA22X1 U30357 ( .IN1(n26574), .IN2(n28665), .IN3(n26527), .IN4(n28667), .Q(
        n26474) );
  OA22X1 U30358 ( .IN1(n26575), .IN2(n28664), .IN3(n26532), .IN4(n28666), .Q(
        n26473) );
  OA22X1 U30359 ( .IN1(n26560), .IN2(n28663), .IN3(n26566), .IN4(n28668), .Q(
        n26472) );
  OA22X1 U30360 ( .IN1(n26558), .IN2(n28662), .IN3(n26578), .IN4(n28661), .Q(
        n26471) );
  NAND4X0 U30361 ( .IN1(n26474), .IN2(n26473), .IN3(n26472), .IN4(n26471), 
        .QN(s6_addr_o[8]) );
  OA22X1 U30362 ( .IN1(n26574), .IN2(n28676), .IN3(n26573), .IN4(n28673), .Q(
        n26478) );
  OA22X1 U30363 ( .IN1(n26572), .IN2(n28679), .IN3(n26576), .IN4(n28674), .Q(
        n26477) );
  OA22X1 U30364 ( .IN1(n26558), .IN2(n28678), .IN3(n26527), .IN4(n28677), .Q(
        n26476) );
  OA22X1 U30365 ( .IN1(n26575), .IN2(n28680), .IN3(n26578), .IN4(n28675), .Q(
        n26475) );
  NAND4X0 U30366 ( .IN1(n26478), .IN2(n26477), .IN3(n26476), .IN4(n26475), 
        .QN(s6_addr_o[9]) );
  OA22X1 U30367 ( .IN1(n26560), .IN2(n28686), .IN3(n26578), .IN4(n28690), .Q(
        n26482) );
  OA22X1 U30368 ( .IN1(n26559), .IN2(n28692), .IN3(n26573), .IN4(n28685), .Q(
        n26481) );
  OA22X1 U30369 ( .IN1(n26532), .IN2(n28688), .IN3(n26574), .IN4(n28687), .Q(
        n26480) );
  OA22X1 U30370 ( .IN1(n26571), .IN2(n28691), .IN3(n26527), .IN4(n28689), .Q(
        n26479) );
  NAND4X0 U30371 ( .IN1(n26482), .IN2(n26481), .IN3(n26480), .IN4(n26479), 
        .QN(s6_addr_o[10]) );
  OA22X1 U30372 ( .IN1(n26566), .IN2(n28701), .IN3(n26527), .IN4(n28699), .Q(
        n26486) );
  OA22X1 U30373 ( .IN1(n26558), .IN2(n28703), .IN3(n26578), .IN4(n28700), .Q(
        n26485) );
  OA22X1 U30374 ( .IN1(n26560), .IN2(n28698), .IN3(n26574), .IN4(n28704), .Q(
        n26484) );
  OA22X1 U30375 ( .IN1(n26559), .IN2(n28702), .IN3(n26532), .IN4(n28697), .Q(
        n26483) );
  NAND4X0 U30376 ( .IN1(n26486), .IN2(n26485), .IN3(n26484), .IN4(n26483), 
        .QN(s6_addr_o[11]) );
  OA22X1 U30377 ( .IN1(n26558), .IN2(n28715), .IN3(n26527), .IN4(n28713), .Q(
        n26490) );
  OA22X1 U30378 ( .IN1(n26574), .IN2(n28716), .IN3(n26566), .IN4(n28709), .Q(
        n26489) );
  OA22X1 U30379 ( .IN1(n26559), .IN2(n28714), .IN3(n26578), .IN4(n28711), .Q(
        n26488) );
  OA22X1 U30380 ( .IN1(n26560), .IN2(n28710), .IN3(n26576), .IN4(n28712), .Q(
        n26487) );
  NAND4X0 U30381 ( .IN1(n26490), .IN2(n26489), .IN3(n26488), .IN4(n26487), 
        .QN(s6_addr_o[12]) );
  OA22X1 U30382 ( .IN1(n26575), .IN2(n28722), .IN3(n26558), .IN4(n28721), .Q(
        n26494) );
  OA22X1 U30383 ( .IN1(n26566), .IN2(n28723), .IN3(n26527), .IN4(n28727), .Q(
        n26493) );
  OA22X1 U30384 ( .IN1(n26572), .IN2(n28728), .IN3(n26532), .IN4(n28726), .Q(
        n26492) );
  OA22X1 U30385 ( .IN1(n26565), .IN2(n28724), .IN3(n26578), .IN4(n28725), .Q(
        n26491) );
  NAND4X0 U30386 ( .IN1(n26494), .IN2(n26493), .IN3(n26492), .IN4(n26491), 
        .QN(s6_addr_o[13]) );
  OA22X1 U30387 ( .IN1(n26565), .IN2(n28735), .IN3(n26578), .IN4(n28733), .Q(
        n26498) );
  OA22X1 U30388 ( .IN1(n26575), .IN2(n28734), .IN3(n26560), .IN4(n28738), .Q(
        n26497) );
  OA22X1 U30389 ( .IN1(n26566), .IN2(n28740), .IN3(n26527), .IN4(n28739), .Q(
        n26496) );
  OA22X1 U30390 ( .IN1(n26576), .IN2(n28736), .IN3(n26558), .IN4(n28737), .Q(
        n26495) );
  NAND4X0 U30391 ( .IN1(n26498), .IN2(n26497), .IN3(n26496), .IN4(n26495), 
        .QN(s6_addr_o[14]) );
  OA22X1 U30392 ( .IN1(n26573), .IN2(n28747), .IN3(n26578), .IN4(n28749), .Q(
        n26502) );
  OA22X1 U30393 ( .IN1(n26558), .IN2(n28751), .IN3(n26527), .IN4(n28745), .Q(
        n26501) );
  OA22X1 U30394 ( .IN1(n26559), .IN2(n28746), .IN3(n26565), .IN4(n28752), .Q(
        n26500) );
  OA22X1 U30395 ( .IN1(n26572), .IN2(n28748), .IN3(n26576), .IN4(n28750), .Q(
        n26499) );
  NAND4X0 U30396 ( .IN1(n26502), .IN2(n26501), .IN3(n26500), .IN4(n26499), 
        .QN(s6_addr_o[15]) );
  OA22X1 U30397 ( .IN1(n26572), .IN2(n28762), .IN3(n26573), .IN4(n28759), .Q(
        n26506) );
  OA22X1 U30398 ( .IN1(n26532), .IN2(n28760), .IN3(n26527), .IN4(n28763), .Q(
        n26505) );
  OA22X1 U30399 ( .IN1(n26565), .IN2(n28761), .IN3(n26571), .IN4(n28757), .Q(
        n26504) );
  OA22X1 U30400 ( .IN1(n26559), .IN2(n28758), .IN3(n26578), .IN4(n28764), .Q(
        n26503) );
  NAND4X0 U30401 ( .IN1(n26506), .IN2(n26505), .IN3(n26504), .IN4(n26503), 
        .QN(s6_addr_o[16]) );
  OA22X1 U30402 ( .IN1(n26559), .IN2(n28772), .IN3(n26566), .IN4(n28775), .Q(
        n26510) );
  OA22X1 U30403 ( .IN1(n26558), .IN2(n28771), .IN3(n26578), .IN4(n28770), .Q(
        n26509) );
  OA22X1 U30404 ( .IN1(n26572), .IN2(n28776), .IN3(n26532), .IN4(n28774), .Q(
        n26508) );
  OA22X1 U30405 ( .IN1(n26574), .IN2(n28773), .IN3(n26527), .IN4(n28769), .Q(
        n26507) );
  NAND4X0 U30406 ( .IN1(n26510), .IN2(n26509), .IN3(n26508), .IN4(n26507), 
        .QN(s6_addr_o[17]) );
  OA22X1 U30407 ( .IN1(n26532), .IN2(n28787), .IN3(n26578), .IN4(n28785), .Q(
        n26514) );
  OA22X1 U30408 ( .IN1(n26560), .IN2(n28788), .IN3(n26574), .IN4(n28782), .Q(
        n26513) );
  OA22X1 U30409 ( .IN1(n26575), .IN2(n28786), .IN3(n26527), .IN4(n28781), .Q(
        n26512) );
  OA22X1 U30410 ( .IN1(n26566), .IN2(n28784), .IN3(n26571), .IN4(n28783), .Q(
        n26511) );
  NAND4X0 U30411 ( .IN1(n26514), .IN2(n26513), .IN3(n26512), .IN4(n26511), 
        .QN(s6_addr_o[18]) );
  OA22X1 U30412 ( .IN1(n26574), .IN2(n28794), .IN3(n26527), .IN4(n28799), .Q(
        n26518) );
  OA22X1 U30413 ( .IN1(n26573), .IN2(n28797), .IN3(n26558), .IN4(n28795), .Q(
        n26517) );
  OA22X1 U30414 ( .IN1(n26559), .IN2(n28796), .IN3(n26560), .IN4(n28800), .Q(
        n26516) );
  OA22X1 U30415 ( .IN1(n26576), .IN2(n28798), .IN3(n26578), .IN4(n28793), .Q(
        n26515) );
  NAND4X0 U30416 ( .IN1(n26518), .IN2(n26517), .IN3(n26516), .IN4(n26515), 
        .QN(s6_addr_o[19]) );
  OA22X1 U30417 ( .IN1(n26575), .IN2(n28812), .IN3(n26527), .IN4(n28805), .Q(
        n26522) );
  OA22X1 U30418 ( .IN1(n26566), .IN2(n28806), .IN3(n26541), .IN4(n28809), .Q(
        n26521) );
  OA22X1 U30419 ( .IN1(n26565), .IN2(n28810), .IN3(n26571), .IN4(n28811), .Q(
        n26520) );
  OA22X1 U30420 ( .IN1(n26560), .IN2(n28808), .IN3(n26532), .IN4(n28807), .Q(
        n26519) );
  NAND4X0 U30421 ( .IN1(n26522), .IN2(n26521), .IN3(n26520), .IN4(n26519), 
        .QN(s6_addr_o[20]) );
  OA22X1 U30422 ( .IN1(n26575), .IN2(n28822), .IN3(n26565), .IN4(n28819), .Q(
        n26526) );
  OA22X1 U30423 ( .IN1(n26572), .IN2(n28824), .IN3(n26576), .IN4(n28820), .Q(
        n26525) );
  OA22X1 U30424 ( .IN1(n26573), .IN2(n28821), .IN3(n26558), .IN4(n28823), .Q(
        n26524) );
  OA22X1 U30425 ( .IN1(n26578), .IN2(n28818), .IN3(n26527), .IN4(n28817), .Q(
        n26523) );
  NAND4X0 U30426 ( .IN1(n26526), .IN2(n26525), .IN3(n26524), .IN4(n26523), 
        .QN(s6_addr_o[21]) );
  OA22X1 U30427 ( .IN1(n26572), .IN2(n28832), .IN3(n26576), .IN4(n28831), .Q(
        n26531) );
  OA22X1 U30428 ( .IN1(n26559), .IN2(n28833), .IN3(n26566), .IN4(n28836), .Q(
        n26530) );
  OA22X1 U30429 ( .IN1(n26565), .IN2(n28838), .IN3(n26541), .IN4(n28837), .Q(
        n26529) );
  OA22X1 U30430 ( .IN1(n26571), .IN2(n28834), .IN3(n26527), .IN4(n28829), .Q(
        n26528) );
  NAND4X0 U30431 ( .IN1(n26531), .IN2(n26530), .IN3(n26529), .IN4(n26528), 
        .QN(s6_addr_o[22]) );
  OA22X1 U30432 ( .IN1(n26578), .IN2(n28846), .IN3(n26577), .IN4(n28851), .Q(
        n26536) );
  OA22X1 U30433 ( .IN1(n26566), .IN2(n28852), .IN3(n26558), .IN4(n28849), .Q(
        n26535) );
  OA22X1 U30434 ( .IN1(n26572), .IN2(n28845), .IN3(n26532), .IN4(n28843), .Q(
        n26534) );
  OA22X1 U30435 ( .IN1(n26559), .IN2(n28848), .IN3(n26565), .IN4(n28850), .Q(
        n26533) );
  NAND4X0 U30436 ( .IN1(n26536), .IN2(n26535), .IN3(n26534), .IN4(n26533), 
        .QN(s6_addr_o[23]) );
  OA22X1 U30437 ( .IN1(n28858), .IN2(n26576), .IN3(n28859), .IN4(n26571), .Q(
        n26540) );
  OA22X1 U30438 ( .IN1(n28857), .IN2(n26565), .IN3(n28861), .IN4(n26573), .Q(
        n26539) );
  OA22X1 U30439 ( .IN1(n28860), .IN2(n26577), .IN3(n28863), .IN4(n26575), .Q(
        n26538) );
  OA22X1 U30440 ( .IN1(n28865), .IN2(n26578), .IN3(n28864), .IN4(n26560), .Q(
        n26537) );
  NAND4X0 U30441 ( .IN1(n26540), .IN2(n26539), .IN3(n26538), .IN4(n26537), 
        .QN(s6_addr_o[24]) );
  OA22X1 U30442 ( .IN1(n28875), .IN2(n26577), .IN3(n28872), .IN4(n26573), .Q(
        n26545) );
  OA22X1 U30443 ( .IN1(n28873), .IN2(n26576), .IN3(n28871), .IN4(n26541), .Q(
        n26544) );
  OA22X1 U30444 ( .IN1(n28877), .IN2(n26560), .IN3(n28870), .IN4(n26575), .Q(
        n26543) );
  OA22X1 U30445 ( .IN1(n28876), .IN2(n26558), .IN3(n28874), .IN4(n26574), .Q(
        n26542) );
  NAND4X0 U30446 ( .IN1(n26545), .IN2(n26544), .IN3(n26543), .IN4(n26542), 
        .QN(s6_addr_o[25]) );
  OA22X1 U30447 ( .IN1(n28887), .IN2(n26572), .IN3(n28889), .IN4(n26577), .Q(
        n26549) );
  OA22X1 U30448 ( .IN1(n28885), .IN2(n26576), .IN3(n28888), .IN4(n26558), .Q(
        n26548) );
  OA22X1 U30449 ( .IN1(n28884), .IN2(n26575), .IN3(n28882), .IN4(n26565), .Q(
        n26547) );
  OA22X1 U30450 ( .IN1(n28883), .IN2(n26578), .IN3(n28886), .IN4(n26566), .Q(
        n26546) );
  NAND4X0 U30451 ( .IN1(n26549), .IN2(n26548), .IN3(n26547), .IN4(n26546), 
        .QN(s6_addr_o[26]) );
  OA22X1 U30452 ( .IN1(n28896), .IN2(n26571), .IN3(n28901), .IN4(n26565), .Q(
        n26553) );
  OA22X1 U30453 ( .IN1(n28897), .IN2(n26578), .IN3(n28894), .IN4(n26575), .Q(
        n26552) );
  OA22X1 U30454 ( .IN1(n28895), .IN2(n26560), .IN3(n28898), .IN4(n26577), .Q(
        n26551) );
  OA22X1 U30455 ( .IN1(n28899), .IN2(n26576), .IN3(n28900), .IN4(n26566), .Q(
        n26550) );
  NAND4X0 U30456 ( .IN1(n26553), .IN2(n26552), .IN3(n26551), .IN4(n26550), 
        .QN(s6_addr_o[27]) );
  OA22X1 U30457 ( .IN1(n28907), .IN2(n26578), .IN3(n28913), .IN4(n26577), .Q(
        n26557) );
  OA22X1 U30458 ( .IN1(n28911), .IN2(n26560), .IN3(n28912), .IN4(n26575), .Q(
        n26556) );
  OA22X1 U30459 ( .IN1(n28909), .IN2(n26576), .IN3(n28908), .IN4(n26574), .Q(
        n26555) );
  OA22X1 U30460 ( .IN1(n28910), .IN2(n26558), .IN3(n28906), .IN4(n26573), .Q(
        n26554) );
  NAND4X0 U30461 ( .IN1(n26557), .IN2(n26556), .IN3(n26555), .IN4(n26554), 
        .QN(s6_addr_o[28]) );
  OA22X1 U30462 ( .IN1(n28926), .IN2(n26576), .IN3(n28920), .IN4(n26558), .Q(
        n26564) );
  OA22X1 U30463 ( .IN1(n28925), .IN2(n26559), .IN3(n28923), .IN4(n26566), .Q(
        n26563) );
  OA22X1 U30464 ( .IN1(n28922), .IN2(n26578), .IN3(n28924), .IN4(n26560), .Q(
        n26562) );
  OA22X1 U30465 ( .IN1(n28921), .IN2(n26577), .IN3(n28919), .IN4(n26574), .Q(
        n26561) );
  NAND4X0 U30466 ( .IN1(n26564), .IN2(n26563), .IN3(n26562), .IN4(n26561), 
        .QN(s6_addr_o[29]) );
  OA22X1 U30467 ( .IN1(n28932), .IN2(n26576), .IN3(n28931), .IN4(n26575), .Q(
        n26570) );
  OA22X1 U30468 ( .IN1(n28935), .IN2(n26572), .IN3(n28940), .IN4(n26565), .Q(
        n26569) );
  OA22X1 U30469 ( .IN1(n28937), .IN2(n26578), .IN3(n28933), .IN4(n26577), .Q(
        n26568) );
  OA22X1 U30470 ( .IN1(n28936), .IN2(n26571), .IN3(n28939), .IN4(n26566), .Q(
        n26567) );
  NAND4X0 U30471 ( .IN1(n26570), .IN2(n26569), .IN3(n26568), .IN4(n26567), 
        .QN(s6_addr_o[30]) );
  OA22X1 U30472 ( .IN1(n28952), .IN2(n26572), .IN3(n28954), .IN4(n26571), .Q(
        n26582) );
  OA22X1 U30473 ( .IN1(n28958), .IN2(n26574), .IN3(n28946), .IN4(n26573), .Q(
        n26581) );
  OA22X1 U30474 ( .IN1(n28948), .IN2(n26576), .IN3(n28950), .IN4(n26575), .Q(
        n26580) );
  OA22X1 U30475 ( .IN1(n28956), .IN2(n26578), .IN3(n28960), .IN4(n26577), .Q(
        n26579) );
  NAND4X0 U30476 ( .IN1(n26582), .IN2(n26581), .IN3(n26580), .IN4(n26579), 
        .QN(s6_addr_o[31]) );
  INVX0 U30477 ( .INP(n26583), .ZN(n26585) );
  OA22X1 U30478 ( .IN1(n29254), .IN2(n26585), .IN3(n29311), .IN4(n26584), .Q(
        n26596) );
  OA22X1 U30479 ( .IN1(n29368), .IN2(n26587), .IN3(n29330), .IN4(n26586), .Q(
        n26595) );
  INVX0 U30480 ( .INP(n26588), .ZN(n26590) );
  OA22X1 U30481 ( .IN1(n29235), .IN2(n26590), .IN3(n29292), .IN4(n26589), .Q(
        n26594) );
  OA22X1 U30482 ( .IN1(n29273), .IN2(n26592), .IN3(n29349), .IN4(n26591), .Q(
        n26593) );
  NAND4X0 U30483 ( .IN1(n26596), .IN2(n26595), .IN3(n26594), .IN4(n26593), 
        .QN(s5_stb_o) );
  INVX0 U30484 ( .INP(n29055), .ZN(n26882) );
  INVX0 U30485 ( .INP(n29063), .ZN(n26881) );
  OA22X1 U30486 ( .IN1(n26882), .IN2(n28123), .IN3(n26881), .IN4(n28122), .Q(
        n26600) );
  INVX0 U30487 ( .INP(n29064), .ZN(n26883) );
  INVX0 U30488 ( .INP(n29057), .ZN(n26880) );
  OA22X1 U30489 ( .IN1(n26883), .IN2(n28126), .IN3(n26880), .IN4(n28127), .Q(
        n26599) );
  INVX0 U30490 ( .INP(n29066), .ZN(n26842) );
  INVX0 U30491 ( .INP(n29058), .ZN(n26872) );
  OA22X1 U30492 ( .IN1(n26842), .IN2(n28124), .IN3(n26872), .IN4(n28128), .Q(
        n26598) );
  INVX0 U30493 ( .INP(n29056), .ZN(n26868) );
  INVX0 U30494 ( .INP(n26833), .ZN(n29065) );
  INVX0 U30495 ( .INP(n29065), .ZN(n26877) );
  OA22X1 U30496 ( .IN1(n26868), .IN2(n28125), .IN3(n26877), .IN4(n28121), .Q(
        n26597) );
  NAND4X0 U30497 ( .IN1(n26600), .IN2(n26599), .IN3(n26598), .IN4(n26597), 
        .QN(s5_we_o) );
  INVX0 U30498 ( .INP(n29064), .ZN(n26870) );
  OA22X1 U30499 ( .IN1(n26870), .IN2(n28139), .IN3(n26833), .IN4(n28135), .Q(
        n26604) );
  OA22X1 U30500 ( .IN1(n26879), .IN2(n28134), .IN3(n26872), .IN4(n28140), .Q(
        n26603) );
  INVX0 U30501 ( .INP(n29057), .ZN(n26871) );
  OA22X1 U30502 ( .IN1(n26882), .IN2(n28133), .IN3(n26871), .IN4(n28137), .Q(
        n26602) );
  OA22X1 U30503 ( .IN1(n26881), .IN2(n28138), .IN3(n26868), .IN4(n28136), .Q(
        n26601) );
  NAND4X0 U30504 ( .IN1(n26604), .IN2(n26603), .IN3(n26602), .IN4(n26601), 
        .QN(s5_data_o[0]) );
  INVX0 U30505 ( .INP(n29056), .ZN(n26884) );
  OA22X1 U30506 ( .IN1(n26870), .IN2(n28145), .IN3(n26884), .IN4(n28152), .Q(
        n26608) );
  OA22X1 U30507 ( .IN1(n26842), .IN2(n28150), .IN3(n26833), .IN4(n28147), .Q(
        n26607) );
  OA22X1 U30508 ( .IN1(n26878), .IN2(n28146), .IN3(n26881), .IN4(n28149), .Q(
        n26606) );
  INVX0 U30509 ( .INP(n29055), .ZN(n26869) );
  OA22X1 U30510 ( .IN1(n26869), .IN2(n28148), .IN3(n26871), .IN4(n28151), .Q(
        n26605) );
  NAND4X0 U30511 ( .IN1(n26608), .IN2(n26607), .IN3(n26606), .IN4(n26605), 
        .QN(s5_data_o[1]) );
  OA22X1 U30512 ( .IN1(n26879), .IN2(n28160), .IN3(n26884), .IN4(n28162), .Q(
        n26612) );
  OA22X1 U30513 ( .IN1(n26882), .IN2(n28163), .IN3(n26870), .IN4(n28159), .Q(
        n26611) );
  INVX0 U30514 ( .INP(n29063), .ZN(n26863) );
  OA22X1 U30515 ( .IN1(n26863), .IN2(n28158), .IN3(n26871), .IN4(n28157), .Q(
        n26610) );
  OA22X1 U30516 ( .IN1(n26872), .IN2(n28164), .IN3(n26833), .IN4(n28161), .Q(
        n26609) );
  NAND4X0 U30517 ( .IN1(n26612), .IN2(n26611), .IN3(n26610), .IN4(n26609), 
        .QN(s5_data_o[2]) );
  OA22X1 U30518 ( .IN1(n26882), .IN2(n28176), .IN3(n26870), .IN4(n28170), .Q(
        n26616) );
  OA22X1 U30519 ( .IN1(n26842), .IN2(n28172), .IN3(n26872), .IN4(n28174), .Q(
        n26615) );
  OA22X1 U30520 ( .IN1(n26880), .IN2(n28169), .IN3(n26833), .IN4(n28173), .Q(
        n26614) );
  OA22X1 U30521 ( .IN1(n26881), .IN2(n28171), .IN3(n26884), .IN4(n28175), .Q(
        n26613) );
  NAND4X0 U30522 ( .IN1(n26616), .IN2(n26615), .IN3(n26614), .IN4(n26613), 
        .QN(s5_data_o[3]) );
  OA22X1 U30523 ( .IN1(n26869), .IN2(n28186), .IN3(n26884), .IN4(n28183), .Q(
        n26620) );
  OA22X1 U30524 ( .IN1(n26883), .IN2(n28188), .IN3(n26881), .IN4(n28185), .Q(
        n26619) );
  OA22X1 U30525 ( .IN1(n26879), .IN2(n28182), .IN3(n26833), .IN4(n28181), .Q(
        n26618) );
  OA22X1 U30526 ( .IN1(n26878), .IN2(n28184), .IN3(n26871), .IN4(n28187), .Q(
        n26617) );
  NAND4X0 U30527 ( .IN1(n26620), .IN2(n26619), .IN3(n26618), .IN4(n26617), 
        .QN(s5_data_o[4]) );
  OA22X1 U30528 ( .IN1(n26842), .IN2(n28196), .IN3(n26884), .IN4(n28197), .Q(
        n26624) );
  OA22X1 U30529 ( .IN1(n26869), .IN2(n28194), .IN3(n26833), .IN4(n28199), .Q(
        n26623) );
  OA22X1 U30530 ( .IN1(n26872), .IN2(n28200), .IN3(n26881), .IN4(n28198), .Q(
        n26622) );
  OA22X1 U30531 ( .IN1(n26870), .IN2(n28193), .IN3(n26871), .IN4(n28195), .Q(
        n26621) );
  NAND4X0 U30532 ( .IN1(n26624), .IN2(n26623), .IN3(n26622), .IN4(n26621), 
        .QN(s5_data_o[5]) );
  OA22X1 U30533 ( .IN1(n26882), .IN2(n28206), .IN3(n26871), .IN4(n28210), .Q(
        n26628) );
  OA22X1 U30534 ( .IN1(n26879), .IN2(n28208), .IN3(n26872), .IN4(n28207), .Q(
        n26627) );
  OA22X1 U30535 ( .IN1(n26863), .IN2(n28211), .IN3(n26833), .IN4(n28209), .Q(
        n26626) );
  OA22X1 U30536 ( .IN1(n26870), .IN2(n28212), .IN3(n26884), .IN4(n28205), .Q(
        n26625) );
  NAND4X0 U30537 ( .IN1(n26628), .IN2(n26627), .IN3(n26626), .IN4(n26625), 
        .QN(s5_data_o[6]) );
  OA22X1 U30538 ( .IN1(n26881), .IN2(n28217), .IN3(n26884), .IN4(n28223), .Q(
        n26632) );
  OA22X1 U30539 ( .IN1(n26869), .IN2(n28224), .IN3(n26877), .IN4(n28221), .Q(
        n26631) );
  OA22X1 U30540 ( .IN1(n26842), .IN2(n28220), .IN3(n26872), .IN4(n28219), .Q(
        n26630) );
  OA22X1 U30541 ( .IN1(n26870), .IN2(n28218), .IN3(n26871), .IN4(n28222), .Q(
        n26629) );
  NAND4X0 U30542 ( .IN1(n26632), .IN2(n26631), .IN3(n26630), .IN4(n26629), 
        .QN(s5_data_o[7]) );
  OA22X1 U30543 ( .IN1(n26871), .IN2(n28233), .IN3(n26877), .IN4(n28235), .Q(
        n26636) );
  OA22X1 U30544 ( .IN1(n26863), .IN2(n28236), .IN3(n26884), .IN4(n28229), .Q(
        n26635) );
  OA22X1 U30545 ( .IN1(n26842), .IN2(n28230), .IN3(n26872), .IN4(n28232), .Q(
        n26634) );
  OA22X1 U30546 ( .IN1(n26869), .IN2(n28231), .IN3(n26870), .IN4(n28234), .Q(
        n26633) );
  NAND4X0 U30547 ( .IN1(n26636), .IN2(n26635), .IN3(n26634), .IN4(n26633), 
        .QN(s5_data_o[8]) );
  OA22X1 U30548 ( .IN1(n26878), .IN2(n28244), .IN3(n26877), .IN4(n28247), .Q(
        n26640) );
  OA22X1 U30549 ( .IN1(n26881), .IN2(n28241), .IN3(n26871), .IN4(n28243), .Q(
        n26639) );
  OA22X1 U30550 ( .IN1(n26879), .IN2(n28242), .IN3(n26869), .IN4(n28246), .Q(
        n26638) );
  OA22X1 U30551 ( .IN1(n26870), .IN2(n28248), .IN3(n26868), .IN4(n28245), .Q(
        n26637) );
  NAND4X0 U30552 ( .IN1(n26640), .IN2(n26639), .IN3(n26638), .IN4(n26637), 
        .QN(s5_data_o[9]) );
  OA22X1 U30553 ( .IN1(n26872), .IN2(n28257), .IN3(n26868), .IN4(n28255), .Q(
        n26644) );
  OA22X1 U30554 ( .IN1(n26882), .IN2(n28260), .IN3(n26870), .IN4(n28256), .Q(
        n26643) );
  OA22X1 U30555 ( .IN1(n26842), .IN2(n28258), .IN3(n26871), .IN4(n28253), .Q(
        n26642) );
  OA22X1 U30556 ( .IN1(n26863), .IN2(n28254), .IN3(n26877), .IN4(n28259), .Q(
        n26641) );
  NAND4X0 U30557 ( .IN1(n26644), .IN2(n26643), .IN3(n26642), .IN4(n26641), 
        .QN(s5_data_o[10]) );
  OA22X1 U30558 ( .IN1(n26879), .IN2(n28266), .IN3(n26884), .IN4(n28270), .Q(
        n26648) );
  OA22X1 U30559 ( .IN1(n26878), .IN2(n28272), .IN3(n26869), .IN4(n28265), .Q(
        n26647) );
  OA22X1 U30560 ( .IN1(n26881), .IN2(n28268), .IN3(n26880), .IN4(n28267), .Q(
        n26646) );
  OA22X1 U30561 ( .IN1(n26883), .IN2(n28271), .IN3(n26877), .IN4(n28269), .Q(
        n26645) );
  NAND4X0 U30562 ( .IN1(n26648), .IN2(n26647), .IN3(n26646), .IN4(n26645), 
        .QN(s5_data_o[11]) );
  OA22X1 U30563 ( .IN1(n26863), .IN2(n28283), .IN3(n26880), .IN4(n28279), .Q(
        n26652) );
  OA22X1 U30564 ( .IN1(n26842), .IN2(n28284), .IN3(n26869), .IN4(n28280), .Q(
        n26651) );
  OA22X1 U30565 ( .IN1(n26870), .IN2(n28282), .IN3(n26877), .IN4(n28277), .Q(
        n26650) );
  OA22X1 U30566 ( .IN1(n26872), .IN2(n28278), .IN3(n26868), .IN4(n28281), .Q(
        n26649) );
  NAND4X0 U30567 ( .IN1(n26652), .IN2(n26651), .IN3(n26650), .IN4(n26649), 
        .QN(s5_data_o[12]) );
  OA22X1 U30568 ( .IN1(n26878), .IN2(n28294), .IN3(n26877), .IN4(n28295), .Q(
        n26656) );
  OA22X1 U30569 ( .IN1(n26882), .IN2(n28296), .IN3(n26870), .IN4(n28292), .Q(
        n26655) );
  OA22X1 U30570 ( .IN1(n26881), .IN2(n28289), .IN3(n26884), .IN4(n28293), .Q(
        n26654) );
  OA22X1 U30571 ( .IN1(n26879), .IN2(n28290), .IN3(n26880), .IN4(n28291), .Q(
        n26653) );
  NAND4X0 U30572 ( .IN1(n26656), .IN2(n26655), .IN3(n26654), .IN4(n26653), 
        .QN(s5_data_o[13]) );
  OA22X1 U30573 ( .IN1(n26878), .IN2(n28304), .IN3(n26880), .IN4(n28301), .Q(
        n26660) );
  OA22X1 U30574 ( .IN1(n26869), .IN2(n28308), .IN3(n26877), .IN4(n28303), .Q(
        n26659) );
  OA22X1 U30575 ( .IN1(n26842), .IN2(n28306), .IN3(n26863), .IN4(n28307), .Q(
        n26658) );
  OA22X1 U30576 ( .IN1(n26870), .IN2(n28305), .IN3(n26884), .IN4(n28302), .Q(
        n26657) );
  NAND4X0 U30577 ( .IN1(n26660), .IN2(n26659), .IN3(n26658), .IN4(n26657), 
        .QN(s5_data_o[14]) );
  OA22X1 U30578 ( .IN1(n26872), .IN2(n28315), .IN3(n26869), .IN4(n28314), .Q(
        n26664) );
  OA22X1 U30579 ( .IN1(n26842), .IN2(n28316), .IN3(n26880), .IN4(n28317), .Q(
        n26663) );
  OA22X1 U30580 ( .IN1(n26863), .IN2(n28320), .IN3(n26877), .IN4(n28319), .Q(
        n26662) );
  OA22X1 U30581 ( .IN1(n26870), .IN2(n28313), .IN3(n26868), .IN4(n28318), .Q(
        n26661) );
  NAND4X0 U30582 ( .IN1(n26664), .IN2(n26663), .IN3(n26662), .IN4(n26661), 
        .QN(s5_data_o[15]) );
  OA22X1 U30583 ( .IN1(n26878), .IN2(n28332), .IN3(n26869), .IN4(n28331), .Q(
        n26668) );
  OA22X1 U30584 ( .IN1(n26868), .IN2(n28325), .IN3(n26880), .IN4(n28328), .Q(
        n26667) );
  OA22X1 U30585 ( .IN1(n26883), .IN2(n28326), .IN3(n26863), .IN4(n28329), .Q(
        n26666) );
  OA22X1 U30586 ( .IN1(n26842), .IN2(n28330), .IN3(n26877), .IN4(n28327), .Q(
        n26665) );
  NAND4X0 U30587 ( .IN1(n26668), .IN2(n26667), .IN3(n26666), .IN4(n26665), 
        .QN(s5_data_o[16]) );
  OA22X1 U30588 ( .IN1(n26884), .IN2(n28339), .IN3(n26877), .IN4(n28341), .Q(
        n26672) );
  OA22X1 U30589 ( .IN1(n26842), .IN2(n28340), .IN3(n26880), .IN4(n28343), .Q(
        n26671) );
  OA22X1 U30590 ( .IN1(n26878), .IN2(n28344), .IN3(n26869), .IN4(n28342), .Q(
        n26670) );
  OA22X1 U30591 ( .IN1(n26883), .IN2(n28338), .IN3(n26881), .IN4(n28337), .Q(
        n26669) );
  NAND4X0 U30592 ( .IN1(n26672), .IN2(n26671), .IN3(n26670), .IN4(n26669), 
        .QN(s5_data_o[17]) );
  OA22X1 U30593 ( .IN1(n26863), .IN2(n28354), .IN3(n26877), .IN4(n28353), .Q(
        n26676) );
  OA22X1 U30594 ( .IN1(n26842), .IN2(n28352), .IN3(n26872), .IN4(n28356), .Q(
        n26675) );
  OA22X1 U30595 ( .IN1(n26869), .IN2(n28350), .IN3(n26880), .IN4(n28351), .Q(
        n26674) );
  OA22X1 U30596 ( .IN1(n26883), .IN2(n28355), .IN3(n26868), .IN4(n28349), .Q(
        n26673) );
  NAND4X0 U30597 ( .IN1(n26676), .IN2(n26675), .IN3(n26674), .IN4(n26673), 
        .QN(s5_data_o[18]) );
  OA22X1 U30598 ( .IN1(n26842), .IN2(n28366), .IN3(n26884), .IN4(n28361), .Q(
        n26680) );
  OA22X1 U30599 ( .IN1(n26870), .IN2(n28363), .IN3(n26863), .IN4(n28365), .Q(
        n26679) );
  OA22X1 U30600 ( .IN1(n26880), .IN2(n28368), .IN3(n26877), .IN4(n28367), .Q(
        n26678) );
  OA22X1 U30601 ( .IN1(n26878), .IN2(n28364), .IN3(n26869), .IN4(n28362), .Q(
        n26677) );
  NAND4X0 U30602 ( .IN1(n26680), .IN2(n26679), .IN3(n26678), .IN4(n26677), 
        .QN(s5_data_o[19]) );
  OA22X1 U30603 ( .IN1(n26842), .IN2(n28378), .IN3(n26863), .IN4(n28376), .Q(
        n26684) );
  OA22X1 U30604 ( .IN1(n26878), .IN2(n28377), .IN3(n26877), .IN4(n28375), .Q(
        n26683) );
  OA22X1 U30605 ( .IN1(n26882), .IN2(n28374), .IN3(n26870), .IN4(n28373), .Q(
        n26682) );
  OA22X1 U30606 ( .IN1(n26868), .IN2(n28380), .IN3(n26880), .IN4(n28379), .Q(
        n26681) );
  NAND4X0 U30607 ( .IN1(n26684), .IN2(n26683), .IN3(n26682), .IN4(n26681), 
        .QN(s5_data_o[20]) );
  OA22X1 U30608 ( .IN1(n26878), .IN2(n28386), .IN3(n26881), .IN4(n28387), .Q(
        n26688) );
  OA22X1 U30609 ( .IN1(n26842), .IN2(n28392), .IN3(n26880), .IN4(n28389), .Q(
        n26687) );
  OA22X1 U30610 ( .IN1(n26869), .IN2(n28390), .IN3(n26877), .IN4(n28391), .Q(
        n26686) );
  OA22X1 U30611 ( .IN1(n26883), .IN2(n28388), .IN3(n26868), .IN4(n28385), .Q(
        n26685) );
  NAND4X0 U30612 ( .IN1(n26688), .IN2(n26687), .IN3(n26686), .IN4(n26685), 
        .QN(s5_data_o[21]) );
  OA22X1 U30613 ( .IN1(n26882), .IN2(n28404), .IN3(n26880), .IN4(n28401), .Q(
        n26692) );
  OA22X1 U30614 ( .IN1(n26842), .IN2(n28400), .IN3(n26870), .IN4(n28403), .Q(
        n26691) );
  OA22X1 U30615 ( .IN1(n26863), .IN2(n28398), .IN3(n26877), .IN4(n28397), .Q(
        n26690) );
  OA22X1 U30616 ( .IN1(n26878), .IN2(n28402), .IN3(n26884), .IN4(n28399), .Q(
        n26689) );
  NAND4X0 U30617 ( .IN1(n26692), .IN2(n26691), .IN3(n26690), .IN4(n26689), 
        .QN(s5_data_o[22]) );
  OA22X1 U30618 ( .IN1(n26870), .IN2(n28413), .IN3(n26881), .IN4(n28410), .Q(
        n26696) );
  OA22X1 U30619 ( .IN1(n26871), .IN2(n28409), .IN3(n26833), .IN4(n28411), .Q(
        n26695) );
  OA22X1 U30620 ( .IN1(n26878), .IN2(n28415), .IN3(n26884), .IN4(n28412), .Q(
        n26694) );
  OA22X1 U30621 ( .IN1(n26842), .IN2(n28416), .IN3(n26869), .IN4(n28414), .Q(
        n26693) );
  NAND4X0 U30622 ( .IN1(n26696), .IN2(n26695), .IN3(n26694), .IN4(n26693), 
        .QN(s5_data_o[23]) );
  OA22X1 U30623 ( .IN1(n26842), .IN2(n28426), .IN3(n26863), .IN4(n28425), .Q(
        n26700) );
  OA22X1 U30624 ( .IN1(n26882), .IN2(n28422), .IN3(n26880), .IN4(n28427), .Q(
        n26699) );
  OA22X1 U30625 ( .IN1(n26878), .IN2(n28424), .IN3(n26833), .IN4(n28423), .Q(
        n26698) );
  OA22X1 U30626 ( .IN1(n26883), .IN2(n28421), .IN3(n26868), .IN4(n28428), .Q(
        n26697) );
  NAND4X0 U30627 ( .IN1(n26700), .IN2(n26699), .IN3(n26698), .IN4(n26697), 
        .QN(s5_data_o[24]) );
  OA22X1 U30628 ( .IN1(n26871), .IN2(n28436), .IN3(n26833), .IN4(n28435), .Q(
        n26704) );
  OA22X1 U30629 ( .IN1(n26842), .IN2(n28438), .IN3(n26869), .IN4(n28434), .Q(
        n26703) );
  OA22X1 U30630 ( .IN1(n26878), .IN2(n28440), .IN3(n26863), .IN4(n28433), .Q(
        n26702) );
  OA22X1 U30631 ( .IN1(n26870), .IN2(n28439), .IN3(n26868), .IN4(n28437), .Q(
        n26701) );
  NAND4X0 U30632 ( .IN1(n26704), .IN2(n26703), .IN3(n26702), .IN4(n26701), 
        .QN(s5_data_o[25]) );
  OA22X1 U30633 ( .IN1(n26878), .IN2(n28451), .IN3(n26880), .IN4(n28447), .Q(
        n26708) );
  OA22X1 U30634 ( .IN1(n26842), .IN2(n28452), .IN3(n26833), .IN4(n28445), .Q(
        n26707) );
  OA22X1 U30635 ( .IN1(n26863), .IN2(n28449), .IN3(n26884), .IN4(n28448), .Q(
        n26706) );
  OA22X1 U30636 ( .IN1(n26869), .IN2(n28450), .IN3(n26870), .IN4(n28446), .Q(
        n26705) );
  NAND4X0 U30637 ( .IN1(n26708), .IN2(n26707), .IN3(n26706), .IN4(n26705), 
        .QN(s5_data_o[26]) );
  OA22X1 U30638 ( .IN1(n26842), .IN2(n28462), .IN3(n26872), .IN4(n28461), .Q(
        n26712) );
  OA22X1 U30639 ( .IN1(n26869), .IN2(n28464), .IN3(n26833), .IN4(n28459), .Q(
        n26711) );
  OA22X1 U30640 ( .IN1(n26883), .IN2(n28458), .IN3(n26863), .IN4(n28457), .Q(
        n26710) );
  OA22X1 U30641 ( .IN1(n26884), .IN2(n28463), .IN3(n26880), .IN4(n28460), .Q(
        n26709) );
  NAND4X0 U30642 ( .IN1(n26712), .IN2(n26711), .IN3(n26710), .IN4(n26709), 
        .QN(s5_data_o[27]) );
  OA22X1 U30643 ( .IN1(n26869), .IN2(n28472), .IN3(n26880), .IN4(n28469), .Q(
        n26716) );
  OA22X1 U30644 ( .IN1(n26879), .IN2(n28474), .IN3(n26868), .IN4(n28475), .Q(
        n26715) );
  OA22X1 U30645 ( .IN1(n26878), .IN2(n28476), .IN3(n26881), .IN4(n28471), .Q(
        n26714) );
  OA22X1 U30646 ( .IN1(n26870), .IN2(n28470), .IN3(n26833), .IN4(n28473), .Q(
        n26713) );
  NAND4X0 U30647 ( .IN1(n26716), .IN2(n26715), .IN3(n26714), .IN4(n26713), 
        .QN(s5_data_o[28]) );
  OA22X1 U30648 ( .IN1(n26879), .IN2(n28484), .IN3(n26878), .IN4(n28482), .Q(
        n26720) );
  OA22X1 U30649 ( .IN1(n26883), .IN2(n28486), .IN3(n26833), .IN4(n28481), .Q(
        n26719) );
  OA22X1 U30650 ( .IN1(n26863), .IN2(n28487), .IN3(n26884), .IN4(n28483), .Q(
        n26718) );
  OA22X1 U30651 ( .IN1(n26882), .IN2(n28488), .IN3(n26880), .IN4(n28485), .Q(
        n26717) );
  NAND4X0 U30652 ( .IN1(n26720), .IN2(n26719), .IN3(n26718), .IN4(n26717), 
        .QN(s5_data_o[29]) );
  OA22X1 U30653 ( .IN1(n26880), .IN2(n28500), .IN3(n26833), .IN4(n28499), .Q(
        n26724) );
  OA22X1 U30654 ( .IN1(n26879), .IN2(n28494), .IN3(n26884), .IN4(n28495), .Q(
        n26723) );
  OA22X1 U30655 ( .IN1(n26869), .IN2(n28497), .IN3(n26881), .IN4(n28493), .Q(
        n26722) );
  OA22X1 U30656 ( .IN1(n26878), .IN2(n28498), .IN3(n26883), .IN4(n28496), .Q(
        n26721) );
  NAND4X0 U30657 ( .IN1(n26724), .IN2(n26723), .IN3(n26722), .IN4(n26721), 
        .QN(s5_data_o[30]) );
  OA22X1 U30658 ( .IN1(n26870), .IN2(n28505), .IN3(n26884), .IN4(n28508), .Q(
        n26728) );
  OA22X1 U30659 ( .IN1(n26869), .IN2(n28506), .IN3(n26863), .IN4(n28512), .Q(
        n26727) );
  OA22X1 U30660 ( .IN1(n26879), .IN2(n28510), .IN3(n26872), .IN4(n28509), .Q(
        n26726) );
  OA22X1 U30661 ( .IN1(n26880), .IN2(n28511), .IN3(n26833), .IN4(n28507), .Q(
        n26725) );
  NAND4X0 U30662 ( .IN1(n26728), .IN2(n26727), .IN3(n26726), .IN4(n26725), 
        .QN(s5_data_o[31]) );
  OA22X1 U30663 ( .IN1(n26879), .IN2(n28518), .IN3(n26883), .IN4(n28524), .Q(
        n26732) );
  OA22X1 U30664 ( .IN1(n26878), .IN2(n28517), .IN3(n26871), .IN4(n28521), .Q(
        n26731) );
  OA22X1 U30665 ( .IN1(n26863), .IN2(n28523), .IN3(n26884), .IN4(n28520), .Q(
        n26730) );
  OA22X1 U30666 ( .IN1(n26882), .IN2(n28522), .IN3(n26833), .IN4(n28519), .Q(
        n26729) );
  NAND4X0 U30667 ( .IN1(n26732), .IN2(n26731), .IN3(n26730), .IN4(n26729), 
        .QN(s5_sel_o[0]) );
  OA22X1 U30668 ( .IN1(n26883), .IN2(n28536), .IN3(n26884), .IN4(n28533), .Q(
        n26736) );
  OA22X1 U30669 ( .IN1(n26882), .IN2(n28530), .IN3(n26833), .IN4(n28529), .Q(
        n26735) );
  OA22X1 U30670 ( .IN1(n26879), .IN2(n28534), .IN3(n26871), .IN4(n28531), .Q(
        n26734) );
  OA22X1 U30671 ( .IN1(n26872), .IN2(n28532), .IN3(n26863), .IN4(n28535), .Q(
        n26733) );
  NAND4X0 U30672 ( .IN1(n26736), .IN2(n26735), .IN3(n26734), .IN4(n26733), 
        .QN(s5_sel_o[1]) );
  OA22X1 U30673 ( .IN1(n26879), .IN2(n28544), .IN3(n26869), .IN4(n28543), .Q(
        n26740) );
  OA22X1 U30674 ( .IN1(n26872), .IN2(n28546), .IN3(n26884), .IN4(n28542), .Q(
        n26739) );
  OA22X1 U30675 ( .IN1(n26870), .IN2(n28548), .IN3(n26871), .IN4(n28545), .Q(
        n26738) );
  OA22X1 U30676 ( .IN1(n26863), .IN2(n28547), .IN3(n26833), .IN4(n28541), .Q(
        n26737) );
  NAND4X0 U30677 ( .IN1(n26740), .IN2(n26739), .IN3(n26738), .IN4(n26737), 
        .QN(s5_sel_o[2]) );
  OA22X1 U30678 ( .IN1(n26883), .IN2(n28557), .IN3(n26833), .IN4(n28555), .Q(
        n26744) );
  OA22X1 U30679 ( .IN1(n26869), .IN2(n28553), .IN3(n26884), .IN4(n28560), .Q(
        n26743) );
  OA22X1 U30680 ( .IN1(n26863), .IN2(n28556), .IN3(n26871), .IN4(n28559), .Q(
        n26742) );
  OA22X1 U30681 ( .IN1(n26842), .IN2(n28558), .IN3(n26872), .IN4(n28554), .Q(
        n26741) );
  NAND4X0 U30682 ( .IN1(n26744), .IN2(n26743), .IN3(n26742), .IN4(n26741), 
        .QN(s5_sel_o[3]) );
  OA22X1 U30683 ( .IN1(n26842), .IN2(n28572), .IN3(n26872), .IN4(n28570), .Q(
        n26748) );
  OA22X1 U30684 ( .IN1(n26870), .IN2(n28566), .IN3(n26884), .IN4(n28567), .Q(
        n26747) );
  OA22X1 U30685 ( .IN1(n26882), .IN2(n28571), .IN3(n26881), .IN4(n28568), .Q(
        n26746) );
  OA22X1 U30686 ( .IN1(n26871), .IN2(n28565), .IN3(n26833), .IN4(n28569), .Q(
        n26745) );
  NAND4X0 U30687 ( .IN1(n26748), .IN2(n26747), .IN3(n26746), .IN4(n26745), 
        .QN(s5_addr_o[0]) );
  OA22X1 U30688 ( .IN1(n26882), .IN2(n28582), .IN3(n26833), .IN4(n28583), .Q(
        n26752) );
  OA22X1 U30689 ( .IN1(n26868), .IN2(n28584), .IN3(n26871), .IN4(n28577), .Q(
        n26751) );
  OA22X1 U30690 ( .IN1(n26879), .IN2(n28580), .IN3(n26870), .IN4(n28581), .Q(
        n26750) );
  OA22X1 U30691 ( .IN1(n26872), .IN2(n28578), .IN3(n26863), .IN4(n28579), .Q(
        n26749) );
  NAND4X0 U30692 ( .IN1(n26752), .IN2(n26751), .IN3(n26750), .IN4(n26749), 
        .QN(s5_addr_o[1]) );
  OA22X1 U30693 ( .IN1(n28596), .IN2(n26877), .IN3(n28590), .IN4(n26881), .Q(
        n26756) );
  OA22X1 U30694 ( .IN1(n28594), .IN2(n26882), .IN3(n28593), .IN4(n26868), .Q(
        n26755) );
  OA22X1 U30695 ( .IN1(n28589), .IN2(n26872), .IN3(n28595), .IN4(n26871), .Q(
        n26754) );
  OA22X1 U30696 ( .IN1(n28592), .IN2(n26883), .IN3(n28591), .IN4(n26879), .Q(
        n26753) );
  NAND4X0 U30697 ( .IN1(n26756), .IN2(n26755), .IN3(n26754), .IN4(n26753), 
        .QN(s5_addr_o[2]) );
  OA22X1 U30698 ( .IN1(n28604), .IN2(n26869), .IN3(n28606), .IN4(n26863), .Q(
        n26760) );
  OA22X1 U30699 ( .IN1(n28608), .IN2(n26877), .IN3(n28607), .IN4(n26883), .Q(
        n26759) );
  OA22X1 U30700 ( .IN1(n28602), .IN2(n26884), .IN3(n28601), .IN4(n26879), .Q(
        n26758) );
  OA22X1 U30701 ( .IN1(n28605), .IN2(n26872), .IN3(n28603), .IN4(n26880), .Q(
        n26757) );
  NAND4X0 U30702 ( .IN1(n26760), .IN2(n26759), .IN3(n26758), .IN4(n26757), 
        .QN(s5_addr_o[3]) );
  OA22X1 U30703 ( .IN1(n28620), .IN2(n26871), .IN3(n28614), .IN4(n26868), .Q(
        n26764) );
  OA22X1 U30704 ( .IN1(n28618), .IN2(n26883), .IN3(n28615), .IN4(n26881), .Q(
        n26763) );
  OA22X1 U30705 ( .IN1(n28619), .IN2(n26877), .IN3(n28617), .IN4(n26879), .Q(
        n26762) );
  OA22X1 U30706 ( .IN1(n28616), .IN2(n26878), .IN3(n28613), .IN4(n26869), .Q(
        n26761) );
  NAND4X0 U30707 ( .IN1(n26764), .IN2(n26763), .IN3(n26762), .IN4(n26761), 
        .QN(s5_addr_o[4]) );
  OA22X1 U30708 ( .IN1(n28627), .IN2(n26868), .IN3(n28629), .IN4(n26879), .Q(
        n26768) );
  OA22X1 U30709 ( .IN1(n28628), .IN2(n26880), .IN3(n28626), .IN4(n26883), .Q(
        n26767) );
  OA22X1 U30710 ( .IN1(n28631), .IN2(n26863), .IN3(n28625), .IN4(n26877), .Q(
        n26766) );
  OA22X1 U30711 ( .IN1(n28632), .IN2(n26882), .IN3(n28630), .IN4(n26878), .Q(
        n26765) );
  NAND4X0 U30712 ( .IN1(n26768), .IN2(n26767), .IN3(n26766), .IN4(n26765), 
        .QN(s5_addr_o[5]) );
  OA22X1 U30713 ( .IN1(n26879), .IN2(n28642), .IN3(n26870), .IN4(n28643), .Q(
        n26772) );
  OA22X1 U30714 ( .IN1(n26872), .IN2(n28640), .IN3(n26884), .IN4(n28637), .Q(
        n26771) );
  OA22X1 U30715 ( .IN1(n26882), .IN2(n28644), .IN3(n26871), .IN4(n28641), .Q(
        n26770) );
  OA22X1 U30716 ( .IN1(n26863), .IN2(n28638), .IN3(n26833), .IN4(n28639), .Q(
        n26769) );
  NAND4X0 U30717 ( .IN1(n26772), .IN2(n26771), .IN3(n26770), .IN4(n26769), 
        .QN(s5_addr_o[6]) );
  OA22X1 U30718 ( .IN1(n26883), .IN2(n28653), .IN3(n26884), .IN4(n28649), .Q(
        n26776) );
  OA22X1 U30719 ( .IN1(n26879), .IN2(n28654), .IN3(n26871), .IN4(n28651), .Q(
        n26775) );
  OA22X1 U30720 ( .IN1(n26882), .IN2(n28656), .IN3(n26881), .IN4(n28650), .Q(
        n26774) );
  OA22X1 U30721 ( .IN1(n26872), .IN2(n28652), .IN3(n26833), .IN4(n28655), .Q(
        n26773) );
  NAND4X0 U30722 ( .IN1(n26776), .IN2(n26775), .IN3(n26774), .IN4(n26773), 
        .QN(s5_addr_o[7]) );
  OA22X1 U30723 ( .IN1(n26872), .IN2(n28663), .IN3(n26869), .IN4(n28666), .Q(
        n26780) );
  OA22X1 U30724 ( .IN1(n26880), .IN2(n28661), .IN3(n26833), .IN4(n28667), .Q(
        n26779) );
  OA22X1 U30725 ( .IN1(n26870), .IN2(n28665), .IN3(n26868), .IN4(n28662), .Q(
        n26778) );
  OA22X1 U30726 ( .IN1(n26842), .IN2(n28664), .IN3(n26881), .IN4(n28668), .Q(
        n26777) );
  NAND4X0 U30727 ( .IN1(n26780), .IN2(n26779), .IN3(n26778), .IN4(n26777), 
        .QN(s5_addr_o[8]) );
  OA22X1 U30728 ( .IN1(n26883), .IN2(n28676), .IN3(n26833), .IN4(n28677), .Q(
        n26784) );
  OA22X1 U30729 ( .IN1(n26872), .IN2(n28679), .IN3(n26881), .IN4(n28673), .Q(
        n26783) );
  OA22X1 U30730 ( .IN1(n26882), .IN2(n28674), .IN3(n26868), .IN4(n28678), .Q(
        n26782) );
  OA22X1 U30731 ( .IN1(n26842), .IN2(n28680), .IN3(n26871), .IN4(n28675), .Q(
        n26781) );
  NAND4X0 U30732 ( .IN1(n26784), .IN2(n26783), .IN3(n26782), .IN4(n26781), 
        .QN(s5_addr_o[9]) );
  OA22X1 U30733 ( .IN1(n26878), .IN2(n28686), .IN3(n26880), .IN4(n28690), .Q(
        n26788) );
  OA22X1 U30734 ( .IN1(n26882), .IN2(n28688), .IN3(n26884), .IN4(n28691), .Q(
        n26787) );
  OA22X1 U30735 ( .IN1(n26879), .IN2(n28692), .IN3(n26863), .IN4(n28685), .Q(
        n26786) );
  OA22X1 U30736 ( .IN1(n26883), .IN2(n28687), .IN3(n26833), .IN4(n28689), .Q(
        n26785) );
  NAND4X0 U30737 ( .IN1(n26788), .IN2(n26787), .IN3(n26786), .IN4(n26785), 
        .QN(s5_addr_o[10]) );
  OA22X1 U30738 ( .IN1(n26878), .IN2(n28698), .IN3(n26884), .IN4(n28703), .Q(
        n26792) );
  OA22X1 U30739 ( .IN1(n26870), .IN2(n28704), .IN3(n26871), .IN4(n28700), .Q(
        n26791) );
  OA22X1 U30740 ( .IN1(n26879), .IN2(n28702), .IN3(n26881), .IN4(n28701), .Q(
        n26790) );
  OA22X1 U30741 ( .IN1(n26882), .IN2(n28697), .IN3(n26833), .IN4(n28699), .Q(
        n26789) );
  NAND4X0 U30742 ( .IN1(n26792), .IN2(n26791), .IN3(n26790), .IN4(n26789), 
        .QN(s5_addr_o[11]) );
  OA22X1 U30743 ( .IN1(n26872), .IN2(n28710), .IN3(n26868), .IN4(n28715), .Q(
        n26796) );
  OA22X1 U30744 ( .IN1(n26863), .IN2(n28709), .IN3(n26880), .IN4(n28711), .Q(
        n26795) );
  OA22X1 U30745 ( .IN1(n26879), .IN2(n28714), .IN3(n26833), .IN4(n28713), .Q(
        n26794) );
  OA22X1 U30746 ( .IN1(n26882), .IN2(n28712), .IN3(n26870), .IN4(n28716), .Q(
        n26793) );
  NAND4X0 U30747 ( .IN1(n26796), .IN2(n26795), .IN3(n26794), .IN4(n26793), 
        .QN(s5_addr_o[12]) );
  OA22X1 U30748 ( .IN1(n26882), .IN2(n28726), .IN3(n26870), .IN4(n28724), .Q(
        n26800) );
  OA22X1 U30749 ( .IN1(n26842), .IN2(n28722), .IN3(n26868), .IN4(n28721), .Q(
        n26799) );
  OA22X1 U30750 ( .IN1(n26872), .IN2(n28728), .IN3(n26833), .IN4(n28727), .Q(
        n26798) );
  OA22X1 U30751 ( .IN1(n26863), .IN2(n28723), .IN3(n26871), .IN4(n28725), .Q(
        n26797) );
  NAND4X0 U30752 ( .IN1(n26800), .IN2(n26799), .IN3(n26798), .IN4(n26797), 
        .QN(s5_addr_o[13]) );
  OA22X1 U30753 ( .IN1(n26879), .IN2(n28734), .IN3(n26872), .IN4(n28738), .Q(
        n26804) );
  OA22X1 U30754 ( .IN1(n26880), .IN2(n28733), .IN3(n26833), .IN4(n28739), .Q(
        n26803) );
  OA22X1 U30755 ( .IN1(n26882), .IN2(n28736), .IN3(n26868), .IN4(n28737), .Q(
        n26802) );
  OA22X1 U30756 ( .IN1(n26883), .IN2(n28735), .IN3(n26863), .IN4(n28740), .Q(
        n26801) );
  NAND4X0 U30757 ( .IN1(n26804), .IN2(n26803), .IN3(n26802), .IN4(n26801), 
        .QN(s5_addr_o[14]) );
  OA22X1 U30758 ( .IN1(n26842), .IN2(n28746), .IN3(n26870), .IN4(n28752), .Q(
        n26808) );
  OA22X1 U30759 ( .IN1(n26878), .IN2(n28748), .IN3(n26884), .IN4(n28751), .Q(
        n26807) );
  OA22X1 U30760 ( .IN1(n26869), .IN2(n28750), .IN3(n26833), .IN4(n28745), .Q(
        n26806) );
  OA22X1 U30761 ( .IN1(n26881), .IN2(n28747), .IN3(n26880), .IN4(n28749), .Q(
        n26805) );
  NAND4X0 U30762 ( .IN1(n26808), .IN2(n26807), .IN3(n26806), .IN4(n26805), 
        .QN(s5_addr_o[15]) );
  OA22X1 U30763 ( .IN1(n26878), .IN2(n28762), .IN3(n26881), .IN4(n28759), .Q(
        n26812) );
  OA22X1 U30764 ( .IN1(n26842), .IN2(n28758), .IN3(n26868), .IN4(n28757), .Q(
        n26811) );
  OA22X1 U30765 ( .IN1(n26882), .IN2(n28760), .IN3(n26880), .IN4(n28764), .Q(
        n26810) );
  OA22X1 U30766 ( .IN1(n26883), .IN2(n28761), .IN3(n26833), .IN4(n28763), .Q(
        n26809) );
  NAND4X0 U30767 ( .IN1(n26812), .IN2(n26811), .IN3(n26810), .IN4(n26809), 
        .QN(s5_addr_o[16]) );
  OA22X1 U30768 ( .IN1(n26882), .IN2(n28774), .IN3(n26881), .IN4(n28775), .Q(
        n26816) );
  OA22X1 U30769 ( .IN1(n26878), .IN2(n28776), .IN3(n26868), .IN4(n28771), .Q(
        n26815) );
  OA22X1 U30770 ( .IN1(n26883), .IN2(n28773), .IN3(n26833), .IN4(n28769), .Q(
        n26814) );
  OA22X1 U30771 ( .IN1(n26842), .IN2(n28772), .IN3(n26871), .IN4(n28770), .Q(
        n26813) );
  NAND4X0 U30772 ( .IN1(n26816), .IN2(n26815), .IN3(n26814), .IN4(n26813), 
        .QN(s5_addr_o[17]) );
  OA22X1 U30773 ( .IN1(n26883), .IN2(n28782), .IN3(n26833), .IN4(n28781), .Q(
        n26820) );
  OA22X1 U30774 ( .IN1(n26879), .IN2(n28786), .IN3(n26871), .IN4(n28785), .Q(
        n26819) );
  OA22X1 U30775 ( .IN1(n26863), .IN2(n28784), .IN3(n26868), .IN4(n28783), .Q(
        n26818) );
  OA22X1 U30776 ( .IN1(n26878), .IN2(n28788), .IN3(n26869), .IN4(n28787), .Q(
        n26817) );
  NAND4X0 U30777 ( .IN1(n26820), .IN2(n26819), .IN3(n26818), .IN4(n26817), 
        .QN(s5_addr_o[18]) );
  OA22X1 U30778 ( .IN1(n26882), .IN2(n28798), .IN3(n26870), .IN4(n28794), .Q(
        n26824) );
  OA22X1 U30779 ( .IN1(n26872), .IN2(n28800), .IN3(n26868), .IN4(n28795), .Q(
        n26823) );
  OA22X1 U30780 ( .IN1(n26879), .IN2(n28796), .IN3(n26881), .IN4(n28797), .Q(
        n26822) );
  OA22X1 U30781 ( .IN1(n26871), .IN2(n28793), .IN3(n26833), .IN4(n28799), .Q(
        n26821) );
  NAND4X0 U30782 ( .IN1(n26824), .IN2(n26823), .IN3(n26822), .IN4(n26821), 
        .QN(s5_addr_o[19]) );
  OA22X1 U30783 ( .IN1(n26842), .IN2(n28812), .IN3(n26833), .IN4(n28805), .Q(
        n26828) );
  OA22X1 U30784 ( .IN1(n26872), .IN2(n28808), .IN3(n26869), .IN4(n28807), .Q(
        n26827) );
  OA22X1 U30785 ( .IN1(n26883), .IN2(n28810), .IN3(n26881), .IN4(n28806), .Q(
        n26826) );
  OA22X1 U30786 ( .IN1(n26884), .IN2(n28811), .IN3(n26871), .IN4(n28809), .Q(
        n26825) );
  NAND4X0 U30787 ( .IN1(n26828), .IN2(n26827), .IN3(n26826), .IN4(n26825), 
        .QN(s5_addr_o[20]) );
  OA22X1 U30788 ( .IN1(n26872), .IN2(n28824), .IN3(n26869), .IN4(n28820), .Q(
        n26832) );
  OA22X1 U30789 ( .IN1(n26863), .IN2(n28821), .IN3(n26868), .IN4(n28823), .Q(
        n26831) );
  OA22X1 U30790 ( .IN1(n26879), .IN2(n28822), .IN3(n26880), .IN4(n28818), .Q(
        n26830) );
  OA22X1 U30791 ( .IN1(n26883), .IN2(n28819), .IN3(n26833), .IN4(n28817), .Q(
        n26829) );
  NAND4X0 U30792 ( .IN1(n26832), .IN2(n26831), .IN3(n26830), .IN4(n26829), 
        .QN(s5_addr_o[21]) );
  OA22X1 U30793 ( .IN1(n26869), .IN2(n28831), .IN3(n26833), .IN4(n28829), .Q(
        n26837) );
  OA22X1 U30794 ( .IN1(n26883), .IN2(n28838), .IN3(n26871), .IN4(n28837), .Q(
        n26836) );
  OA22X1 U30795 ( .IN1(n26872), .IN2(n28832), .IN3(n26881), .IN4(n28836), .Q(
        n26835) );
  OA22X1 U30796 ( .IN1(n26842), .IN2(n28833), .IN3(n26868), .IN4(n28834), .Q(
        n26834) );
  NAND4X0 U30797 ( .IN1(n26837), .IN2(n26836), .IN3(n26835), .IN4(n26834), 
        .QN(s5_addr_o[22]) );
  OA22X1 U30798 ( .IN1(n26842), .IN2(n28848), .IN3(n26877), .IN4(n28851), .Q(
        n26841) );
  OA22X1 U30799 ( .IN1(n26882), .IN2(n28843), .IN3(n26870), .IN4(n28850), .Q(
        n26840) );
  OA22X1 U30800 ( .IN1(n26878), .IN2(n28845), .IN3(n26868), .IN4(n28849), .Q(
        n26839) );
  OA22X1 U30801 ( .IN1(n26863), .IN2(n28852), .IN3(n26871), .IN4(n28846), .Q(
        n26838) );
  NAND4X0 U30802 ( .IN1(n26841), .IN2(n26840), .IN3(n26839), .IN4(n26838), 
        .QN(s5_addr_o[23]) );
  OA22X1 U30803 ( .IN1(n28865), .IN2(n26871), .IN3(n28857), .IN4(n26870), .Q(
        n26846) );
  OA22X1 U30804 ( .IN1(n28863), .IN2(n26842), .IN3(n28861), .IN4(n26881), .Q(
        n26845) );
  OA22X1 U30805 ( .IN1(n28858), .IN2(n26869), .IN3(n28860), .IN4(n26877), .Q(
        n26844) );
  OA22X1 U30806 ( .IN1(n28864), .IN2(n26878), .IN3(n28859), .IN4(n26868), .Q(
        n26843) );
  NAND4X0 U30807 ( .IN1(n26846), .IN2(n26845), .IN3(n26844), .IN4(n26843), 
        .QN(s5_addr_o[24]) );
  OA22X1 U30808 ( .IN1(n28871), .IN2(n26880), .IN3(n28874), .IN4(n26883), .Q(
        n26850) );
  OA22X1 U30809 ( .IN1(n28877), .IN2(n26872), .IN3(n28875), .IN4(n26877), .Q(
        n26849) );
  OA22X1 U30810 ( .IN1(n28873), .IN2(n26882), .IN3(n28870), .IN4(n26879), .Q(
        n26848) );
  OA22X1 U30811 ( .IN1(n28876), .IN2(n26884), .IN3(n28872), .IN4(n26881), .Q(
        n26847) );
  NAND4X0 U30812 ( .IN1(n26850), .IN2(n26849), .IN3(n26848), .IN4(n26847), 
        .QN(s5_addr_o[25]) );
  OA22X1 U30813 ( .IN1(n28888), .IN2(n26868), .IN3(n28884), .IN4(n26879), .Q(
        n26854) );
  OA22X1 U30814 ( .IN1(n28882), .IN2(n26883), .IN3(n28886), .IN4(n26881), .Q(
        n26853) );
  OA22X1 U30815 ( .IN1(n28885), .IN2(n26869), .IN3(n28887), .IN4(n26872), .Q(
        n26852) );
  OA22X1 U30816 ( .IN1(n28883), .IN2(n26871), .IN3(n28889), .IN4(n26877), .Q(
        n26851) );
  NAND4X0 U30817 ( .IN1(n26854), .IN2(n26853), .IN3(n26852), .IN4(n26851), 
        .QN(s5_addr_o[26]) );
  OA22X1 U30818 ( .IN1(n28895), .IN2(n26878), .IN3(n28896), .IN4(n26868), .Q(
        n26858) );
  OA22X1 U30819 ( .IN1(n28897), .IN2(n26880), .IN3(n28901), .IN4(n26883), .Q(
        n26857) );
  OA22X1 U30820 ( .IN1(n28899), .IN2(n26882), .IN3(n28894), .IN4(n26879), .Q(
        n26856) );
  OA22X1 U30821 ( .IN1(n28898), .IN2(n26877), .IN3(n28900), .IN4(n26881), .Q(
        n26855) );
  NAND4X0 U30822 ( .IN1(n26858), .IN2(n26857), .IN3(n26856), .IN4(n26855), 
        .QN(s5_addr_o[27]) );
  OA22X1 U30823 ( .IN1(n28908), .IN2(n26883), .IN3(n28906), .IN4(n26881), .Q(
        n26862) );
  OA22X1 U30824 ( .IN1(n28909), .IN2(n26869), .IN3(n28911), .IN4(n26878), .Q(
        n26861) );
  OA22X1 U30825 ( .IN1(n28907), .IN2(n26871), .IN3(n28910), .IN4(n26868), .Q(
        n26860) );
  OA22X1 U30826 ( .IN1(n28913), .IN2(n26877), .IN3(n28912), .IN4(n26879), .Q(
        n26859) );
  NAND4X0 U30827 ( .IN1(n26862), .IN2(n26861), .IN3(n26860), .IN4(n26859), 
        .QN(s5_addr_o[28]) );
  OA22X1 U30828 ( .IN1(n28924), .IN2(n26872), .IN3(n28925), .IN4(n26879), .Q(
        n26867) );
  OA22X1 U30829 ( .IN1(n28926), .IN2(n26882), .IN3(n28921), .IN4(n26877), .Q(
        n26866) );
  OA22X1 U30830 ( .IN1(n28922), .IN2(n26880), .IN3(n28920), .IN4(n26868), .Q(
        n26865) );
  OA22X1 U30831 ( .IN1(n28919), .IN2(n26883), .IN3(n28923), .IN4(n26863), .Q(
        n26864) );
  NAND4X0 U30832 ( .IN1(n26867), .IN2(n26866), .IN3(n26865), .IN4(n26864), 
        .QN(s5_addr_o[29]) );
  OA22X1 U30833 ( .IN1(n28933), .IN2(n26877), .IN3(n28936), .IN4(n26868), .Q(
        n26876) );
  OA22X1 U30834 ( .IN1(n28932), .IN2(n26869), .IN3(n28931), .IN4(n26879), .Q(
        n26875) );
  OA22X1 U30835 ( .IN1(n28937), .IN2(n26871), .IN3(n28940), .IN4(n26870), .Q(
        n26874) );
  OA22X1 U30836 ( .IN1(n28935), .IN2(n26872), .IN3(n28939), .IN4(n26881), .Q(
        n26873) );
  NAND4X0 U30837 ( .IN1(n26876), .IN2(n26875), .IN3(n26874), .IN4(n26873), 
        .QN(s5_addr_o[30]) );
  OA22X1 U30838 ( .IN1(n28952), .IN2(n26878), .IN3(n28960), .IN4(n26877), .Q(
        n26888) );
  OA22X1 U30839 ( .IN1(n28956), .IN2(n26880), .IN3(n28950), .IN4(n26879), .Q(
        n26887) );
  OA22X1 U30840 ( .IN1(n28948), .IN2(n26882), .IN3(n28946), .IN4(n26881), .Q(
        n26886) );
  OA22X1 U30841 ( .IN1(n28954), .IN2(n26884), .IN3(n28958), .IN4(n26883), .Q(
        n26885) );
  NAND4X0 U30842 ( .IN1(n26888), .IN2(n26887), .IN3(n26886), .IN4(n26885), 
        .QN(s5_addr_o[31]) );
  OA22X1 U30843 ( .IN1(n29368), .IN2(n26890), .IN3(n29330), .IN4(n26889), .Q(
        n26900) );
  OA22X1 U30844 ( .IN1(n29235), .IN2(n26892), .IN3(n29311), .IN4(n26891), .Q(
        n26899) );
  OA22X1 U30845 ( .IN1(n29273), .IN2(n26894), .IN3(n29292), .IN4(n26893), .Q(
        n26898) );
  OA22X1 U30846 ( .IN1(n29349), .IN2(n26896), .IN3(n29254), .IN4(n26895), .Q(
        n26897) );
  NAND4X0 U30847 ( .IN1(n26900), .IN2(n26899), .IN3(n26898), .IN4(n26897), 
        .QN(s4_stb_o) );
  INVX0 U30848 ( .INP(n29048), .ZN(n27168) );
  INVX0 U30849 ( .INP(n27137), .ZN(n29047) );
  INVX0 U30850 ( .INP(n29047), .ZN(n27188) );
  OA22X1 U30851 ( .IN1(n27168), .IN2(n28122), .IN3(n27188), .IN4(n28121), .Q(
        n26904) );
  INVX0 U30852 ( .INP(n29040), .ZN(n27186) );
  INVX0 U30853 ( .INP(n29045), .ZN(n27167) );
  OA22X1 U30854 ( .IN1(n27186), .IN2(n28128), .IN3(n27167), .IN4(n28125), .Q(
        n26903) );
  INVX0 U30855 ( .INP(n29038), .ZN(n27185) );
  INVX0 U30856 ( .INP(n29046), .ZN(n27175) );
  OA22X1 U30857 ( .IN1(n27185), .IN2(n28124), .IN3(n27175), .IN4(n28126), .Q(
        n26902) );
  INVX0 U30858 ( .INP(n29037), .ZN(n27184) );
  OA22X1 U30859 ( .IN1(n27184), .IN2(n28123), .IN3(n27183), .IN4(n28127), .Q(
        n26901) );
  NAND4X0 U30860 ( .IN1(n26904), .IN2(n26903), .IN3(n26902), .IN4(n26901), 
        .QN(s4_we_o) );
  INVX0 U30861 ( .INP(n29048), .ZN(n27181) );
  OA22X1 U30862 ( .IN1(n27175), .IN2(n28139), .IN3(n27181), .IN4(n28138), .Q(
        n26908) );
  OA22X1 U30863 ( .IN1(n27167), .IN2(n28136), .IN3(n27137), .IN4(n28135), .Q(
        n26907) );
  INVX0 U30864 ( .INP(n29040), .ZN(n27174) );
  OA22X1 U30865 ( .IN1(n27174), .IN2(n28140), .IN3(n27184), .IN4(n28133), .Q(
        n26906) );
  INVX0 U30866 ( .INP(n29038), .ZN(n27150) );
  OA22X1 U30867 ( .IN1(n27150), .IN2(n28134), .IN3(n27183), .IN4(n28137), .Q(
        n26905) );
  NAND4X0 U30868 ( .IN1(n26908), .IN2(n26907), .IN3(n26906), .IN4(n26905), 
        .QN(s4_data_o[0]) );
  OA22X1 U30869 ( .IN1(n27185), .IN2(n28150), .IN3(n27137), .IN4(n28147), .Q(
        n26912) );
  OA22X1 U30870 ( .IN1(n27174), .IN2(n28146), .IN3(n27167), .IN4(n28152), .Q(
        n26911) );
  INVX0 U30871 ( .INP(n29037), .ZN(n27173) );
  OA22X1 U30872 ( .IN1(n27173), .IN2(n28148), .IN3(n27175), .IN4(n28145), .Q(
        n26910) );
  OA22X1 U30873 ( .IN1(n27181), .IN2(n28149), .IN3(n27183), .IN4(n28151), .Q(
        n26909) );
  NAND4X0 U30874 ( .IN1(n26912), .IN2(n26911), .IN3(n26910), .IN4(n26909), 
        .QN(s4_data_o[1]) );
  OA22X1 U30875 ( .IN1(n27174), .IN2(n28164), .IN3(n27137), .IN4(n28161), .Q(
        n26916) );
  OA22X1 U30876 ( .IN1(n27185), .IN2(n28160), .IN3(n27167), .IN4(n28162), .Q(
        n26915) );
  INVX0 U30877 ( .INP(n29046), .ZN(n27187) );
  OA22X1 U30878 ( .IN1(n27187), .IN2(n28159), .IN3(n27181), .IN4(n28158), .Q(
        n26914) );
  OA22X1 U30879 ( .IN1(n27184), .IN2(n28163), .IN3(n27183), .IN4(n28157), .Q(
        n26913) );
  NAND4X0 U30880 ( .IN1(n26916), .IN2(n26915), .IN3(n26914), .IN4(n26913), 
        .QN(s4_data_o[2]) );
  INVX0 U30881 ( .INP(n27183), .ZN(n29039) );
  INVX0 U30882 ( .INP(n29039), .ZN(n27176) );
  OA22X1 U30883 ( .IN1(n27176), .IN2(n28169), .IN3(n27137), .IN4(n28173), .Q(
        n26920) );
  OA22X1 U30884 ( .IN1(n27185), .IN2(n28172), .IN3(n27167), .IN4(n28175), .Q(
        n26919) );
  OA22X1 U30885 ( .IN1(n27174), .IN2(n28174), .IN3(n27184), .IN4(n28176), .Q(
        n26918) );
  OA22X1 U30886 ( .IN1(n27175), .IN2(n28170), .IN3(n27181), .IN4(n28171), .Q(
        n26917) );
  NAND4X0 U30887 ( .IN1(n26920), .IN2(n26919), .IN3(n26918), .IN4(n26917), 
        .QN(s4_data_o[3]) );
  OA22X1 U30888 ( .IN1(n27185), .IN2(n28182), .IN3(n27167), .IN4(n28183), .Q(
        n26924) );
  OA22X1 U30889 ( .IN1(n27187), .IN2(n28188), .IN3(n27137), .IN4(n28181), .Q(
        n26923) );
  OA22X1 U30890 ( .IN1(n27173), .IN2(n28186), .IN3(n27183), .IN4(n28187), .Q(
        n26922) );
  OA22X1 U30891 ( .IN1(n27174), .IN2(n28184), .IN3(n27181), .IN4(n28185), .Q(
        n26921) );
  NAND4X0 U30892 ( .IN1(n26924), .IN2(n26923), .IN3(n26922), .IN4(n26921), 
        .QN(s4_data_o[4]) );
  OA22X1 U30893 ( .IN1(n27174), .IN2(n28200), .IN3(n27167), .IN4(n28197), .Q(
        n26928) );
  OA22X1 U30894 ( .IN1(n27185), .IN2(n28196), .IN3(n27184), .IN4(n28194), .Q(
        n26927) );
  OA22X1 U30895 ( .IN1(n27176), .IN2(n28195), .IN3(n27137), .IN4(n28199), .Q(
        n26926) );
  OA22X1 U30896 ( .IN1(n27175), .IN2(n28193), .IN3(n27181), .IN4(n28198), .Q(
        n26925) );
  NAND4X0 U30897 ( .IN1(n26928), .IN2(n26927), .IN3(n26926), .IN4(n26925), 
        .QN(s4_data_o[5]) );
  OA22X1 U30898 ( .IN1(n27173), .IN2(n28206), .IN3(n27175), .IN4(n28212), .Q(
        n26932) );
  OA22X1 U30899 ( .IN1(n27168), .IN2(n28211), .IN3(n27137), .IN4(n28209), .Q(
        n26931) );
  OA22X1 U30900 ( .IN1(n27174), .IN2(n28207), .IN3(n27167), .IN4(n28205), .Q(
        n26930) );
  OA22X1 U30901 ( .IN1(n27185), .IN2(n28208), .IN3(n27183), .IN4(n28210), .Q(
        n26929) );
  NAND4X0 U30902 ( .IN1(n26932), .IN2(n26931), .IN3(n26930), .IN4(n26929), 
        .QN(s4_data_o[6]) );
  OA22X1 U30903 ( .IN1(n27186), .IN2(n28219), .IN3(n27175), .IN4(n28218), .Q(
        n26936) );
  INVX0 U30904 ( .INP(n29045), .ZN(n27182) );
  OA22X1 U30905 ( .IN1(n27182), .IN2(n28223), .IN3(n27183), .IN4(n28222), .Q(
        n26935) );
  OA22X1 U30906 ( .IN1(n27185), .IN2(n28220), .IN3(n27188), .IN4(n28221), .Q(
        n26934) );
  OA22X1 U30907 ( .IN1(n27184), .IN2(n28224), .IN3(n27181), .IN4(n28217), .Q(
        n26933) );
  NAND4X0 U30908 ( .IN1(n26936), .IN2(n26935), .IN3(n26934), .IN4(n26933), 
        .QN(s4_data_o[7]) );
  OA22X1 U30909 ( .IN1(n27186), .IN2(n28232), .IN3(n27183), .IN4(n28233), .Q(
        n26940) );
  OA22X1 U30910 ( .IN1(n27185), .IN2(n28230), .IN3(n27184), .IN4(n28231), .Q(
        n26939) );
  OA22X1 U30911 ( .IN1(n27187), .IN2(n28234), .IN3(n27188), .IN4(n28235), .Q(
        n26938) );
  OA22X1 U30912 ( .IN1(n27181), .IN2(n28236), .IN3(n27182), .IN4(n28229), .Q(
        n26937) );
  NAND4X0 U30913 ( .IN1(n26940), .IN2(n26939), .IN3(n26938), .IN4(n26937), 
        .QN(s4_data_o[8]) );
  OA22X1 U30914 ( .IN1(n27167), .IN2(n28245), .IN3(n27188), .IN4(n28247), .Q(
        n26944) );
  OA22X1 U30915 ( .IN1(n27184), .IN2(n28246), .IN3(n27175), .IN4(n28248), .Q(
        n26943) );
  OA22X1 U30916 ( .IN1(n27174), .IN2(n28244), .IN3(n27181), .IN4(n28241), .Q(
        n26942) );
  OA22X1 U30917 ( .IN1(n27150), .IN2(n28242), .IN3(n27183), .IN4(n28243), .Q(
        n26941) );
  NAND4X0 U30918 ( .IN1(n26944), .IN2(n26943), .IN3(n26942), .IN4(n26941), 
        .QN(s4_data_o[9]) );
  OA22X1 U30919 ( .IN1(n27185), .IN2(n28258), .IN3(n27184), .IN4(n28260), .Q(
        n26948) );
  OA22X1 U30920 ( .IN1(n27182), .IN2(n28255), .IN3(n27183), .IN4(n28253), .Q(
        n26947) );
  OA22X1 U30921 ( .IN1(n27175), .IN2(n28256), .IN3(n27181), .IN4(n28254), .Q(
        n26946) );
  OA22X1 U30922 ( .IN1(n27174), .IN2(n28257), .IN3(n27188), .IN4(n28259), .Q(
        n26945) );
  NAND4X0 U30923 ( .IN1(n26948), .IN2(n26947), .IN3(n26946), .IN4(n26945), 
        .QN(s4_data_o[10]) );
  OA22X1 U30924 ( .IN1(n27167), .IN2(n28270), .IN3(n27188), .IN4(n28269), .Q(
        n26952) );
  OA22X1 U30925 ( .IN1(n27150), .IN2(n28266), .IN3(n27181), .IN4(n28268), .Q(
        n26951) );
  OA22X1 U30926 ( .IN1(n27186), .IN2(n28272), .IN3(n27175), .IN4(n28271), .Q(
        n26950) );
  OA22X1 U30927 ( .IN1(n27184), .IN2(n28265), .IN3(n27183), .IN4(n28267), .Q(
        n26949) );
  NAND4X0 U30928 ( .IN1(n26952), .IN2(n26951), .IN3(n26950), .IN4(n26949), 
        .QN(s4_data_o[11]) );
  OA22X1 U30929 ( .IN1(n27173), .IN2(n28280), .IN3(n27175), .IN4(n28282), .Q(
        n26956) );
  OA22X1 U30930 ( .IN1(n27186), .IN2(n28278), .IN3(n27168), .IN4(n28283), .Q(
        n26955) );
  OA22X1 U30931 ( .IN1(n27182), .IN2(n28281), .IN3(n27188), .IN4(n28277), .Q(
        n26954) );
  OA22X1 U30932 ( .IN1(n27150), .IN2(n28284), .IN3(n27176), .IN4(n28279), .Q(
        n26953) );
  NAND4X0 U30933 ( .IN1(n26956), .IN2(n26955), .IN3(n26954), .IN4(n26953), 
        .QN(s4_data_o[12]) );
  OA22X1 U30934 ( .IN1(n27184), .IN2(n28296), .IN3(n27181), .IN4(n28289), .Q(
        n26960) );
  OA22X1 U30935 ( .IN1(n27187), .IN2(n28292), .IN3(n27176), .IN4(n28291), .Q(
        n26959) );
  OA22X1 U30936 ( .IN1(n27185), .IN2(n28290), .IN3(n27174), .IN4(n28294), .Q(
        n26958) );
  OA22X1 U30937 ( .IN1(n27167), .IN2(n28293), .IN3(n27188), .IN4(n28295), .Q(
        n26957) );
  NAND4X0 U30938 ( .IN1(n26960), .IN2(n26959), .IN3(n26958), .IN4(n26957), 
        .QN(s4_data_o[13]) );
  OA22X1 U30939 ( .IN1(n27173), .IN2(n28308), .IN3(n27175), .IN4(n28305), .Q(
        n26964) );
  OA22X1 U30940 ( .IN1(n27185), .IN2(n28306), .IN3(n27167), .IN4(n28302), .Q(
        n26963) );
  OA22X1 U30941 ( .IN1(n27176), .IN2(n28301), .IN3(n27188), .IN4(n28303), .Q(
        n26962) );
  OA22X1 U30942 ( .IN1(n27174), .IN2(n28304), .IN3(n27168), .IN4(n28307), .Q(
        n26961) );
  NAND4X0 U30943 ( .IN1(n26964), .IN2(n26963), .IN3(n26962), .IN4(n26961), 
        .QN(s4_data_o[14]) );
  OA22X1 U30944 ( .IN1(n27168), .IN2(n28320), .IN3(n27167), .IN4(n28318), .Q(
        n26968) );
  OA22X1 U30945 ( .IN1(n27186), .IN2(n28315), .IN3(n27173), .IN4(n28314), .Q(
        n26967) );
  OA22X1 U30946 ( .IN1(n27176), .IN2(n28317), .IN3(n27188), .IN4(n28319), .Q(
        n26966) );
  OA22X1 U30947 ( .IN1(n27185), .IN2(n28316), .IN3(n27187), .IN4(n28313), .Q(
        n26965) );
  NAND4X0 U30948 ( .IN1(n26968), .IN2(n26967), .IN3(n26966), .IN4(n26965), 
        .QN(s4_data_o[15]) );
  OA22X1 U30949 ( .IN1(n27186), .IN2(n28332), .IN3(n27188), .IN4(n28327), .Q(
        n26972) );
  OA22X1 U30950 ( .IN1(n27150), .IN2(n28330), .IN3(n27167), .IN4(n28325), .Q(
        n26971) );
  OA22X1 U30951 ( .IN1(n27168), .IN2(n28329), .IN3(n27176), .IN4(n28328), .Q(
        n26970) );
  OA22X1 U30952 ( .IN1(n27184), .IN2(n28331), .IN3(n27187), .IN4(n28326), .Q(
        n26969) );
  NAND4X0 U30953 ( .IN1(n26972), .IN2(n26971), .IN3(n26970), .IN4(n26969), 
        .QN(s4_data_o[16]) );
  OA22X1 U30954 ( .IN1(n27174), .IN2(n28344), .IN3(n27176), .IN4(n28343), .Q(
        n26976) );
  OA22X1 U30955 ( .IN1(n27182), .IN2(n28339), .IN3(n27188), .IN4(n28341), .Q(
        n26975) );
  OA22X1 U30956 ( .IN1(n27173), .IN2(n28342), .IN3(n27168), .IN4(n28337), .Q(
        n26974) );
  OA22X1 U30957 ( .IN1(n27185), .IN2(n28340), .IN3(n27175), .IN4(n28338), .Q(
        n26973) );
  NAND4X0 U30958 ( .IN1(n26976), .IN2(n26975), .IN3(n26974), .IN4(n26973), 
        .QN(s4_data_o[17]) );
  OA22X1 U30959 ( .IN1(n27150), .IN2(n28352), .IN3(n27174), .IN4(n28356), .Q(
        n26980) );
  OA22X1 U30960 ( .IN1(n27173), .IN2(n28350), .IN3(n27167), .IN4(n28349), .Q(
        n26979) );
  OA22X1 U30961 ( .IN1(n27176), .IN2(n28351), .IN3(n27188), .IN4(n28353), .Q(
        n26978) );
  OA22X1 U30962 ( .IN1(n27187), .IN2(n28355), .IN3(n27181), .IN4(n28354), .Q(
        n26977) );
  NAND4X0 U30963 ( .IN1(n26980), .IN2(n26979), .IN3(n26978), .IN4(n26977), 
        .QN(s4_data_o[18]) );
  OA22X1 U30964 ( .IN1(n27167), .IN2(n28361), .IN3(n27188), .IN4(n28367), .Q(
        n26984) );
  OA22X1 U30965 ( .IN1(n27150), .IN2(n28366), .IN3(n27187), .IN4(n28363), .Q(
        n26983) );
  OA22X1 U30966 ( .IN1(n27184), .IN2(n28362), .IN3(n27181), .IN4(n28365), .Q(
        n26982) );
  OA22X1 U30967 ( .IN1(n27174), .IN2(n28364), .IN3(n27176), .IN4(n28368), .Q(
        n26981) );
  NAND4X0 U30968 ( .IN1(n26984), .IN2(n26983), .IN3(n26982), .IN4(n26981), 
        .QN(s4_data_o[19]) );
  OA22X1 U30969 ( .IN1(n27173), .IN2(n28374), .IN3(n27167), .IN4(n28380), .Q(
        n26988) );
  OA22X1 U30970 ( .IN1(n27185), .IN2(n28378), .IN3(n27175), .IN4(n28373), .Q(
        n26987) );
  OA22X1 U30971 ( .IN1(n27186), .IN2(n28377), .IN3(n27176), .IN4(n28379), .Q(
        n26986) );
  OA22X1 U30972 ( .IN1(n27168), .IN2(n28376), .IN3(n27188), .IN4(n28375), .Q(
        n26985) );
  NAND4X0 U30973 ( .IN1(n26988), .IN2(n26987), .IN3(n26986), .IN4(n26985), 
        .QN(s4_data_o[20]) );
  OA22X1 U30974 ( .IN1(n27182), .IN2(n28385), .IN3(n27188), .IN4(n28391), .Q(
        n26992) );
  OA22X1 U30975 ( .IN1(n27174), .IN2(n28386), .IN3(n27168), .IN4(n28387), .Q(
        n26991) );
  OA22X1 U30976 ( .IN1(n27184), .IN2(n28390), .IN3(n27176), .IN4(n28389), .Q(
        n26990) );
  OA22X1 U30977 ( .IN1(n27150), .IN2(n28392), .IN3(n27175), .IN4(n28388), .Q(
        n26989) );
  NAND4X0 U30978 ( .IN1(n26992), .IN2(n26991), .IN3(n26990), .IN4(n26989), 
        .QN(s4_data_o[21]) );
  OA22X1 U30979 ( .IN1(n27150), .IN2(n28400), .IN3(n27176), .IN4(n28401), .Q(
        n26996) );
  OA22X1 U30980 ( .IN1(n27173), .IN2(n28404), .IN3(n27188), .IN4(n28397), .Q(
        n26995) );
  OA22X1 U30981 ( .IN1(n27187), .IN2(n28403), .IN3(n27182), .IN4(n28399), .Q(
        n26994) );
  OA22X1 U30982 ( .IN1(n27186), .IN2(n28402), .IN3(n27181), .IN4(n28398), .Q(
        n26993) );
  NAND4X0 U30983 ( .IN1(n26996), .IN2(n26995), .IN3(n26994), .IN4(n26993), 
        .QN(s4_data_o[22]) );
  OA22X1 U30984 ( .IN1(n27186), .IN2(n28415), .IN3(n27137), .IN4(n28411), .Q(
        n27000) );
  OA22X1 U30985 ( .IN1(n27184), .IN2(n28414), .IN3(n27176), .IN4(n28409), .Q(
        n26999) );
  OA22X1 U30986 ( .IN1(n27150), .IN2(n28416), .IN3(n27168), .IN4(n28410), .Q(
        n26998) );
  OA22X1 U30987 ( .IN1(n27187), .IN2(n28413), .IN3(n27167), .IN4(n28412), .Q(
        n26997) );
  NAND4X0 U30988 ( .IN1(n27000), .IN2(n26999), .IN3(n26998), .IN4(n26997), 
        .QN(s4_data_o[23]) );
  OA22X1 U30989 ( .IN1(n27187), .IN2(n28421), .IN3(n27137), .IN4(n28423), .Q(
        n27004) );
  OA22X1 U30990 ( .IN1(n27173), .IN2(n28422), .IN3(n27168), .IN4(n28425), .Q(
        n27003) );
  OA22X1 U30991 ( .IN1(n27182), .IN2(n28428), .IN3(n27176), .IN4(n28427), .Q(
        n27002) );
  OA22X1 U30992 ( .IN1(n27185), .IN2(n28426), .IN3(n27174), .IN4(n28424), .Q(
        n27001) );
  NAND4X0 U30993 ( .IN1(n27004), .IN2(n27003), .IN3(n27002), .IN4(n27001), 
        .QN(s4_data_o[24]) );
  OA22X1 U30994 ( .IN1(n27185), .IN2(n28438), .IN3(n27174), .IN4(n28440), .Q(
        n27008) );
  OA22X1 U30995 ( .IN1(n27182), .IN2(n28437), .IN3(n27176), .IN4(n28436), .Q(
        n27007) );
  OA22X1 U30996 ( .IN1(n27184), .IN2(n28434), .IN3(n27181), .IN4(n28433), .Q(
        n27006) );
  OA22X1 U30997 ( .IN1(n27187), .IN2(n28439), .IN3(n27137), .IN4(n28435), .Q(
        n27005) );
  NAND4X0 U30998 ( .IN1(n27008), .IN2(n27007), .IN3(n27006), .IN4(n27005), 
        .QN(s4_data_o[25]) );
  OA22X1 U30999 ( .IN1(n27183), .IN2(n28447), .IN3(n27137), .IN4(n28445), .Q(
        n27012) );
  OA22X1 U31000 ( .IN1(n27187), .IN2(n28446), .IN3(n27167), .IN4(n28448), .Q(
        n27011) );
  OA22X1 U31001 ( .IN1(n27150), .IN2(n28452), .IN3(n27174), .IN4(n28451), .Q(
        n27010) );
  OA22X1 U31002 ( .IN1(n27184), .IN2(n28450), .IN3(n27181), .IN4(n28449), .Q(
        n27009) );
  NAND4X0 U31003 ( .IN1(n27012), .IN2(n27011), .IN3(n27010), .IN4(n27009), 
        .QN(s4_data_o[26]) );
  OA22X1 U31004 ( .IN1(n27174), .IN2(n28461), .IN3(n27182), .IN4(n28463), .Q(
        n27016) );
  OA22X1 U31005 ( .IN1(n27168), .IN2(n28457), .IN3(n27176), .IN4(n28460), .Q(
        n27015) );
  OA22X1 U31006 ( .IN1(n27185), .IN2(n28462), .IN3(n27187), .IN4(n28458), .Q(
        n27014) );
  OA22X1 U31007 ( .IN1(n27173), .IN2(n28464), .IN3(n27137), .IN4(n28459), .Q(
        n27013) );
  NAND4X0 U31008 ( .IN1(n27016), .IN2(n27015), .IN3(n27014), .IN4(n27013), 
        .QN(s4_data_o[27]) );
  OA22X1 U31009 ( .IN1(n27185), .IN2(n28474), .IN3(n27176), .IN4(n28469), .Q(
        n27020) );
  OA22X1 U31010 ( .IN1(n27168), .IN2(n28471), .IN3(n27137), .IN4(n28473), .Q(
        n27019) );
  OA22X1 U31011 ( .IN1(n27174), .IN2(n28476), .IN3(n27182), .IN4(n28475), .Q(
        n27018) );
  OA22X1 U31012 ( .IN1(n27173), .IN2(n28472), .IN3(n27187), .IN4(n28470), .Q(
        n27017) );
  NAND4X0 U31013 ( .IN1(n27020), .IN2(n27019), .IN3(n27018), .IN4(n27017), 
        .QN(s4_data_o[28]) );
  OA22X1 U31014 ( .IN1(n27186), .IN2(n28482), .IN3(n27168), .IN4(n28487), .Q(
        n27024) );
  OA22X1 U31015 ( .IN1(n27184), .IN2(n28488), .IN3(n27175), .IN4(n28486), .Q(
        n27023) );
  OA22X1 U31016 ( .IN1(n27182), .IN2(n28483), .IN3(n27176), .IN4(n28485), .Q(
        n27022) );
  OA22X1 U31017 ( .IN1(n27150), .IN2(n28484), .IN3(n27137), .IN4(n28481), .Q(
        n27021) );
  NAND4X0 U31018 ( .IN1(n27024), .IN2(n27023), .IN3(n27022), .IN4(n27021), 
        .QN(s4_data_o[29]) );
  OA22X1 U31019 ( .IN1(n27175), .IN2(n28496), .IN3(n27137), .IN4(n28499), .Q(
        n27028) );
  OA22X1 U31020 ( .IN1(n27150), .IN2(n28494), .IN3(n27176), .IN4(n28500), .Q(
        n27027) );
  OA22X1 U31021 ( .IN1(n27184), .IN2(n28497), .IN3(n27167), .IN4(n28495), .Q(
        n27026) );
  OA22X1 U31022 ( .IN1(n27174), .IN2(n28498), .IN3(n27168), .IN4(n28493), .Q(
        n27025) );
  NAND4X0 U31023 ( .IN1(n27028), .IN2(n27027), .IN3(n27026), .IN4(n27025), 
        .QN(s4_data_o[30]) );
  OA22X1 U31024 ( .IN1(n27168), .IN2(n28512), .IN3(n27137), .IN4(n28507), .Q(
        n27032) );
  OA22X1 U31025 ( .IN1(n27173), .IN2(n28506), .IN3(n27176), .IN4(n28511), .Q(
        n27031) );
  OA22X1 U31026 ( .IN1(n27186), .IN2(n28509), .IN3(n27187), .IN4(n28505), .Q(
        n27030) );
  OA22X1 U31027 ( .IN1(n27185), .IN2(n28510), .IN3(n27167), .IN4(n28508), .Q(
        n27029) );
  NAND4X0 U31028 ( .IN1(n27032), .IN2(n27031), .IN3(n27030), .IN4(n27029), 
        .QN(s4_data_o[31]) );
  OA22X1 U31029 ( .IN1(n27185), .IN2(n28518), .IN3(n27137), .IN4(n28519), .Q(
        n27036) );
  OA22X1 U31030 ( .IN1(n27168), .IN2(n28523), .IN3(n27183), .IN4(n28521), .Q(
        n27035) );
  OA22X1 U31031 ( .IN1(n27187), .IN2(n28524), .IN3(n27182), .IN4(n28520), .Q(
        n27034) );
  OA22X1 U31032 ( .IN1(n27186), .IN2(n28517), .IN3(n27184), .IN4(n28522), .Q(
        n27033) );
  NAND4X0 U31033 ( .IN1(n27036), .IN2(n27035), .IN3(n27034), .IN4(n27033), 
        .QN(s4_sel_o[0]) );
  OA22X1 U31034 ( .IN1(n27174), .IN2(n28532), .IN3(n27183), .IN4(n28531), .Q(
        n27040) );
  OA22X1 U31035 ( .IN1(n27167), .IN2(n28533), .IN3(n27137), .IN4(n28529), .Q(
        n27039) );
  OA22X1 U31036 ( .IN1(n27150), .IN2(n28534), .IN3(n27175), .IN4(n28536), .Q(
        n27038) );
  OA22X1 U31037 ( .IN1(n27173), .IN2(n28530), .IN3(n27181), .IN4(n28535), .Q(
        n27037) );
  NAND4X0 U31038 ( .IN1(n27040), .IN2(n27039), .IN3(n27038), .IN4(n27037), 
        .QN(s4_sel_o[1]) );
  OA22X1 U31039 ( .IN1(n27175), .IN2(n28548), .IN3(n27183), .IN4(n28545), .Q(
        n27044) );
  OA22X1 U31040 ( .IN1(n27150), .IN2(n28544), .IN3(n27137), .IN4(n28541), .Q(
        n27043) );
  OA22X1 U31041 ( .IN1(n27168), .IN2(n28547), .IN3(n27182), .IN4(n28542), .Q(
        n27042) );
  OA22X1 U31042 ( .IN1(n27174), .IN2(n28546), .IN3(n27184), .IN4(n28543), .Q(
        n27041) );
  NAND4X0 U31043 ( .IN1(n27044), .IN2(n27043), .IN3(n27042), .IN4(n27041), 
        .QN(s4_sel_o[2]) );
  OA22X1 U31044 ( .IN1(n27175), .IN2(n28557), .IN3(n27181), .IN4(n28556), .Q(
        n27048) );
  OA22X1 U31045 ( .IN1(n27150), .IN2(n28558), .IN3(n27167), .IN4(n28560), .Q(
        n27047) );
  OA22X1 U31046 ( .IN1(n27173), .IN2(n28553), .IN3(n27137), .IN4(n28555), .Q(
        n27046) );
  OA22X1 U31047 ( .IN1(n27186), .IN2(n28554), .IN3(n27183), .IN4(n28559), .Q(
        n27045) );
  NAND4X0 U31048 ( .IN1(n27048), .IN2(n27047), .IN3(n27046), .IN4(n27045), 
        .QN(s4_sel_o[3]) );
  OA22X1 U31049 ( .IN1(n27186), .IN2(n28570), .IN3(n27175), .IN4(n28566), .Q(
        n27052) );
  OA22X1 U31050 ( .IN1(n27173), .IN2(n28571), .IN3(n27183), .IN4(n28565), .Q(
        n27051) );
  OA22X1 U31051 ( .IN1(n27168), .IN2(n28568), .IN3(n27167), .IN4(n28567), .Q(
        n27050) );
  OA22X1 U31052 ( .IN1(n27150), .IN2(n28572), .IN3(n27137), .IN4(n28569), .Q(
        n27049) );
  NAND4X0 U31053 ( .IN1(n27052), .IN2(n27051), .IN3(n27050), .IN4(n27049), 
        .QN(s4_addr_o[0]) );
  OA22X1 U31054 ( .IN1(n27150), .IN2(n28580), .IN3(n27168), .IN4(n28579), .Q(
        n27056) );
  OA22X1 U31055 ( .IN1(n27173), .IN2(n28582), .IN3(n27182), .IN4(n28584), .Q(
        n27055) );
  OA22X1 U31056 ( .IN1(n27183), .IN2(n28577), .IN3(n27137), .IN4(n28583), .Q(
        n27054) );
  OA22X1 U31057 ( .IN1(n27186), .IN2(n28578), .IN3(n27175), .IN4(n28581), .Q(
        n27053) );
  NAND4X0 U31058 ( .IN1(n27056), .IN2(n27055), .IN3(n27054), .IN4(n27053), 
        .QN(s4_addr_o[1]) );
  OA22X1 U31059 ( .IN1(n28592), .IN2(n27175), .IN3(n28596), .IN4(n27188), .Q(
        n27060) );
  OA22X1 U31060 ( .IN1(n28591), .IN2(n27150), .IN3(n28595), .IN4(n27183), .Q(
        n27059) );
  OA22X1 U31061 ( .IN1(n28590), .IN2(n27181), .IN3(n28593), .IN4(n27182), .Q(
        n27058) );
  OA22X1 U31062 ( .IN1(n28594), .IN2(n27184), .IN3(n28589), .IN4(n27174), .Q(
        n27057) );
  NAND4X0 U31063 ( .IN1(n27060), .IN2(n27059), .IN3(n27058), .IN4(n27057), 
        .QN(s4_addr_o[2]) );
  OA22X1 U31064 ( .IN1(n28604), .IN2(n27173), .IN3(n28606), .IN4(n27181), .Q(
        n27064) );
  OA22X1 U31065 ( .IN1(n28605), .IN2(n27174), .IN3(n28603), .IN4(n27183), .Q(
        n27063) );
  OA22X1 U31066 ( .IN1(n28602), .IN2(n27182), .IN3(n28601), .IN4(n27185), .Q(
        n27062) );
  OA22X1 U31067 ( .IN1(n28608), .IN2(n27188), .IN3(n28607), .IN4(n27175), .Q(
        n27061) );
  NAND4X0 U31068 ( .IN1(n27064), .IN2(n27063), .IN3(n27062), .IN4(n27061), 
        .QN(s4_addr_o[3]) );
  OA22X1 U31069 ( .IN1(n28617), .IN2(n27185), .IN3(n28613), .IN4(n27184), .Q(
        n27068) );
  OA22X1 U31070 ( .IN1(n28619), .IN2(n27188), .IN3(n28615), .IN4(n27181), .Q(
        n27067) );
  OA22X1 U31071 ( .IN1(n28618), .IN2(n27187), .IN3(n28614), .IN4(n27167), .Q(
        n27066) );
  OA22X1 U31072 ( .IN1(n28616), .IN2(n27186), .IN3(n28620), .IN4(n27183), .Q(
        n27065) );
  NAND4X0 U31073 ( .IN1(n27068), .IN2(n27067), .IN3(n27066), .IN4(n27065), 
        .QN(s4_addr_o[4]) );
  OA22X1 U31074 ( .IN1(n28628), .IN2(n27176), .IN3(n28629), .IN4(n27185), .Q(
        n27072) );
  OA22X1 U31075 ( .IN1(n28632), .IN2(n27184), .IN3(n28625), .IN4(n27188), .Q(
        n27071) );
  OA22X1 U31076 ( .IN1(n28627), .IN2(n27182), .IN3(n28630), .IN4(n27174), .Q(
        n27070) );
  OA22X1 U31077 ( .IN1(n28626), .IN2(n27175), .IN3(n28631), .IN4(n27181), .Q(
        n27069) );
  NAND4X0 U31078 ( .IN1(n27072), .IN2(n27071), .IN3(n27070), .IN4(n27069), 
        .QN(s4_addr_o[5]) );
  OA22X1 U31079 ( .IN1(n27173), .IN2(n28644), .IN3(n27183), .IN4(n28641), .Q(
        n27076) );
  OA22X1 U31080 ( .IN1(n27168), .IN2(n28638), .IN3(n27137), .IN4(n28639), .Q(
        n27075) );
  OA22X1 U31081 ( .IN1(n27186), .IN2(n28640), .IN3(n27187), .IN4(n28643), .Q(
        n27074) );
  OA22X1 U31082 ( .IN1(n27150), .IN2(n28642), .IN3(n27167), .IN4(n28637), .Q(
        n27073) );
  NAND4X0 U31083 ( .IN1(n27076), .IN2(n27075), .IN3(n27074), .IN4(n27073), 
        .QN(s4_addr_o[6]) );
  OA22X1 U31084 ( .IN1(n27150), .IN2(n28654), .IN3(n27182), .IN4(n28649), .Q(
        n27080) );
  OA22X1 U31085 ( .IN1(n27183), .IN2(n28651), .IN3(n27137), .IN4(n28655), .Q(
        n27079) );
  OA22X1 U31086 ( .IN1(n27186), .IN2(n28652), .IN3(n27184), .IN4(n28656), .Q(
        n27078) );
  OA22X1 U31087 ( .IN1(n27187), .IN2(n28653), .IN3(n27181), .IN4(n28650), .Q(
        n27077) );
  NAND4X0 U31088 ( .IN1(n27080), .IN2(n27079), .IN3(n27078), .IN4(n27077), 
        .QN(s4_addr_o[7]) );
  OA22X1 U31089 ( .IN1(n27168), .IN2(n28668), .IN3(n27137), .IN4(n28667), .Q(
        n27084) );
  OA22X1 U31090 ( .IN1(n27187), .IN2(n28665), .IN3(n27182), .IN4(n28662), .Q(
        n27083) );
  OA22X1 U31091 ( .IN1(n27150), .IN2(n28664), .IN3(n27174), .IN4(n28663), .Q(
        n27082) );
  OA22X1 U31092 ( .IN1(n27173), .IN2(n28666), .IN3(n27183), .IN4(n28661), .Q(
        n27081) );
  NAND4X0 U31093 ( .IN1(n27084), .IN2(n27083), .IN3(n27082), .IN4(n27081), 
        .QN(s4_addr_o[8]) );
  OA22X1 U31094 ( .IN1(n27186), .IN2(n28679), .IN3(n27167), .IN4(n28678), .Q(
        n27088) );
  OA22X1 U31095 ( .IN1(n27173), .IN2(n28674), .IN3(n27183), .IN4(n28675), .Q(
        n27087) );
  OA22X1 U31096 ( .IN1(n27150), .IN2(n28680), .IN3(n27175), .IN4(n28676), .Q(
        n27086) );
  OA22X1 U31097 ( .IN1(n27168), .IN2(n28673), .IN3(n27137), .IN4(n28677), .Q(
        n27085) );
  NAND4X0 U31098 ( .IN1(n27088), .IN2(n27087), .IN3(n27086), .IN4(n27085), 
        .QN(s4_addr_o[9]) );
  OA22X1 U31099 ( .IN1(n27186), .IN2(n28686), .IN3(n27184), .IN4(n28688), .Q(
        n27092) );
  OA22X1 U31100 ( .IN1(n27168), .IN2(n28685), .IN3(n27167), .IN4(n28691), .Q(
        n27091) );
  OA22X1 U31101 ( .IN1(n27150), .IN2(n28692), .IN3(n27137), .IN4(n28689), .Q(
        n27090) );
  OA22X1 U31102 ( .IN1(n27187), .IN2(n28687), .IN3(n27183), .IN4(n28690), .Q(
        n27089) );
  NAND4X0 U31103 ( .IN1(n27092), .IN2(n27091), .IN3(n27090), .IN4(n27089), 
        .QN(s4_addr_o[10]) );
  OA22X1 U31104 ( .IN1(n27186), .IN2(n28698), .IN3(n27183), .IN4(n28700), .Q(
        n27096) );
  OA22X1 U31105 ( .IN1(n27181), .IN2(n28701), .IN3(n27182), .IN4(n28703), .Q(
        n27095) );
  OA22X1 U31106 ( .IN1(n27173), .IN2(n28697), .IN3(n27175), .IN4(n28704), .Q(
        n27094) );
  OA22X1 U31107 ( .IN1(n27150), .IN2(n28702), .IN3(n27137), .IN4(n28699), .Q(
        n27093) );
  NAND4X0 U31108 ( .IN1(n27096), .IN2(n27095), .IN3(n27094), .IN4(n27093), 
        .QN(s4_addr_o[11]) );
  OA22X1 U31109 ( .IN1(n27168), .IN2(n28709), .IN3(n27137), .IN4(n28713), .Q(
        n27100) );
  OA22X1 U31110 ( .IN1(n27186), .IN2(n28710), .IN3(n27173), .IN4(n28712), .Q(
        n27099) );
  OA22X1 U31111 ( .IN1(n27187), .IN2(n28716), .IN3(n27183), .IN4(n28711), .Q(
        n27098) );
  OA22X1 U31112 ( .IN1(n27150), .IN2(n28714), .IN3(n27167), .IN4(n28715), .Q(
        n27097) );
  NAND4X0 U31113 ( .IN1(n27100), .IN2(n27099), .IN3(n27098), .IN4(n27097), 
        .QN(s4_addr_o[12]) );
  OA22X1 U31114 ( .IN1(n27150), .IN2(n28722), .IN3(n27183), .IN4(n28725), .Q(
        n27104) );
  OA22X1 U31115 ( .IN1(n27175), .IN2(n28724), .IN3(n27168), .IN4(n28723), .Q(
        n27103) );
  OA22X1 U31116 ( .IN1(n27186), .IN2(n28728), .IN3(n27137), .IN4(n28727), .Q(
        n27102) );
  OA22X1 U31117 ( .IN1(n27173), .IN2(n28726), .IN3(n27182), .IN4(n28721), .Q(
        n27101) );
  NAND4X0 U31118 ( .IN1(n27104), .IN2(n27103), .IN3(n27102), .IN4(n27101), 
        .QN(s4_addr_o[13]) );
  OA22X1 U31119 ( .IN1(n27150), .IN2(n28734), .IN3(n27184), .IN4(n28736), .Q(
        n27108) );
  OA22X1 U31120 ( .IN1(n27183), .IN2(n28733), .IN3(n27137), .IN4(n28739), .Q(
        n27107) );
  OA22X1 U31121 ( .IN1(n27186), .IN2(n28738), .IN3(n27181), .IN4(n28740), .Q(
        n27106) );
  OA22X1 U31122 ( .IN1(n27187), .IN2(n28735), .IN3(n27182), .IN4(n28737), .Q(
        n27105) );
  NAND4X0 U31123 ( .IN1(n27108), .IN2(n27107), .IN3(n27106), .IN4(n27105), 
        .QN(s4_addr_o[14]) );
  OA22X1 U31124 ( .IN1(n27186), .IN2(n28748), .IN3(n27184), .IN4(n28750), .Q(
        n27112) );
  OA22X1 U31125 ( .IN1(n27176), .IN2(n28749), .IN3(n27137), .IN4(n28745), .Q(
        n27111) );
  OA22X1 U31126 ( .IN1(n27187), .IN2(n28752), .IN3(n27168), .IN4(n28747), .Q(
        n27110) );
  OA22X1 U31127 ( .IN1(n27150), .IN2(n28746), .IN3(n27167), .IN4(n28751), .Q(
        n27109) );
  NAND4X0 U31128 ( .IN1(n27112), .IN2(n27111), .IN3(n27110), .IN4(n27109), 
        .QN(s4_addr_o[15]) );
  OA22X1 U31129 ( .IN1(n27183), .IN2(n28764), .IN3(n27137), .IN4(n28763), .Q(
        n27116) );
  OA22X1 U31130 ( .IN1(n27186), .IN2(n28762), .IN3(n27184), .IN4(n28760), .Q(
        n27115) );
  OA22X1 U31131 ( .IN1(n27168), .IN2(n28759), .IN3(n27167), .IN4(n28757), .Q(
        n27114) );
  OA22X1 U31132 ( .IN1(n27150), .IN2(n28758), .IN3(n27187), .IN4(n28761), .Q(
        n27113) );
  NAND4X0 U31133 ( .IN1(n27116), .IN2(n27115), .IN3(n27114), .IN4(n27113), 
        .QN(s4_addr_o[16]) );
  OA22X1 U31134 ( .IN1(n27173), .IN2(n28774), .IN3(n27137), .IN4(n28769), .Q(
        n27120) );
  OA22X1 U31135 ( .IN1(n27186), .IN2(n28776), .IN3(n27167), .IN4(n28771), .Q(
        n27119) );
  OA22X1 U31136 ( .IN1(n27181), .IN2(n28775), .IN3(n27183), .IN4(n28770), .Q(
        n27118) );
  OA22X1 U31137 ( .IN1(n27185), .IN2(n28772), .IN3(n27187), .IN4(n28773), .Q(
        n27117) );
  NAND4X0 U31138 ( .IN1(n27120), .IN2(n27119), .IN3(n27118), .IN4(n27117), 
        .QN(s4_addr_o[17]) );
  OA22X1 U31139 ( .IN1(n27173), .IN2(n28787), .IN3(n27183), .IN4(n28785), .Q(
        n27124) );
  OA22X1 U31140 ( .IN1(n27187), .IN2(n28782), .IN3(n27137), .IN4(n28781), .Q(
        n27123) );
  OA22X1 U31141 ( .IN1(n27168), .IN2(n28784), .IN3(n27182), .IN4(n28783), .Q(
        n27122) );
  OA22X1 U31142 ( .IN1(n27150), .IN2(n28786), .IN3(n27174), .IN4(n28788), .Q(
        n27121) );
  NAND4X0 U31143 ( .IN1(n27124), .IN2(n27123), .IN3(n27122), .IN4(n27121), 
        .QN(s4_addr_o[18]) );
  OA22X1 U31144 ( .IN1(n27185), .IN2(n28796), .IN3(n27183), .IN4(n28793), .Q(
        n27128) );
  OA22X1 U31145 ( .IN1(n27182), .IN2(n28795), .IN3(n27137), .IN4(n28799), .Q(
        n27127) );
  OA22X1 U31146 ( .IN1(n27186), .IN2(n28800), .IN3(n27168), .IN4(n28797), .Q(
        n27126) );
  OA22X1 U31147 ( .IN1(n27173), .IN2(n28798), .IN3(n27175), .IN4(n28794), .Q(
        n27125) );
  NAND4X0 U31148 ( .IN1(n27128), .IN2(n27127), .IN3(n27126), .IN4(n27125), 
        .QN(s4_addr_o[19]) );
  OA22X1 U31149 ( .IN1(n27150), .IN2(n28812), .IN3(n27184), .IN4(n28807), .Q(
        n27132) );
  OA22X1 U31150 ( .IN1(n27181), .IN2(n28806), .IN3(n27137), .IN4(n28805), .Q(
        n27131) );
  OA22X1 U31151 ( .IN1(n27182), .IN2(n28811), .IN3(n27183), .IN4(n28809), .Q(
        n27130) );
  OA22X1 U31152 ( .IN1(n27174), .IN2(n28808), .IN3(n27187), .IN4(n28810), .Q(
        n27129) );
  NAND4X0 U31153 ( .IN1(n27132), .IN2(n27131), .IN3(n27130), .IN4(n27129), 
        .QN(s4_addr_o[20]) );
  OA22X1 U31154 ( .IN1(n27185), .IN2(n28822), .IN3(n27167), .IN4(n28823), .Q(
        n27136) );
  OA22X1 U31155 ( .IN1(n27173), .IN2(n28820), .IN3(n27175), .IN4(n28819), .Q(
        n27135) );
  OA22X1 U31156 ( .IN1(n27168), .IN2(n28821), .IN3(n27137), .IN4(n28817), .Q(
        n27134) );
  OA22X1 U31157 ( .IN1(n27186), .IN2(n28824), .IN3(n27183), .IN4(n28818), .Q(
        n27133) );
  NAND4X0 U31158 ( .IN1(n27136), .IN2(n27135), .IN3(n27134), .IN4(n27133), 
        .QN(s4_addr_o[21]) );
  OA22X1 U31159 ( .IN1(n27181), .IN2(n28836), .IN3(n27183), .IN4(n28837), .Q(
        n27141) );
  OA22X1 U31160 ( .IN1(n27173), .IN2(n28831), .IN3(n27167), .IN4(n28834), .Q(
        n27140) );
  OA22X1 U31161 ( .IN1(n27150), .IN2(n28833), .IN3(n27175), .IN4(n28838), .Q(
        n27139) );
  OA22X1 U31162 ( .IN1(n27174), .IN2(n28832), .IN3(n27137), .IN4(n28829), .Q(
        n27138) );
  NAND4X0 U31163 ( .IN1(n27141), .IN2(n27140), .IN3(n27139), .IN4(n27138), 
        .QN(s4_addr_o[22]) );
  OA22X1 U31164 ( .IN1(n27185), .IN2(n28848), .IN3(n27184), .IN4(n28843), .Q(
        n27145) );
  OA22X1 U31165 ( .IN1(n27168), .IN2(n28852), .IN3(n27188), .IN4(n28851), .Q(
        n27144) );
  OA22X1 U31166 ( .IN1(n27182), .IN2(n28849), .IN3(n27183), .IN4(n28846), .Q(
        n27143) );
  OA22X1 U31167 ( .IN1(n27186), .IN2(n28845), .IN3(n27175), .IN4(n28850), .Q(
        n27142) );
  NAND4X0 U31168 ( .IN1(n27145), .IN2(n27144), .IN3(n27143), .IN4(n27142), 
        .QN(s4_addr_o[23]) );
  OA22X1 U31169 ( .IN1(n28864), .IN2(n27174), .IN3(n28860), .IN4(n27188), .Q(
        n27149) );
  OA22X1 U31170 ( .IN1(n28859), .IN2(n27182), .IN3(n28863), .IN4(n27185), .Q(
        n27148) );
  OA22X1 U31171 ( .IN1(n28865), .IN2(n27176), .IN3(n28861), .IN4(n27181), .Q(
        n27147) );
  OA22X1 U31172 ( .IN1(n28858), .IN2(n27173), .IN3(n28857), .IN4(n27187), .Q(
        n27146) );
  NAND4X0 U31173 ( .IN1(n27149), .IN2(n27148), .IN3(n27147), .IN4(n27146), 
        .QN(s4_addr_o[24]) );
  OA22X1 U31174 ( .IN1(n28873), .IN2(n27184), .IN3(n28872), .IN4(n27181), .Q(
        n27154) );
  OA22X1 U31175 ( .IN1(n28870), .IN2(n27150), .IN3(n28874), .IN4(n27175), .Q(
        n27153) );
  OA22X1 U31176 ( .IN1(n28877), .IN2(n27186), .IN3(n28875), .IN4(n27188), .Q(
        n27152) );
  OA22X1 U31177 ( .IN1(n28871), .IN2(n27176), .IN3(n28876), .IN4(n27167), .Q(
        n27151) );
  NAND4X0 U31178 ( .IN1(n27154), .IN2(n27153), .IN3(n27152), .IN4(n27151), 
        .QN(s4_addr_o[25]) );
  OA22X1 U31179 ( .IN1(n28885), .IN2(n27173), .IN3(n28882), .IN4(n27187), .Q(
        n27158) );
  OA22X1 U31180 ( .IN1(n28883), .IN2(n27176), .IN3(n28884), .IN4(n27185), .Q(
        n27157) );
  OA22X1 U31181 ( .IN1(n28887), .IN2(n27174), .IN3(n28889), .IN4(n27188), .Q(
        n27156) );
  OA22X1 U31182 ( .IN1(n28888), .IN2(n27182), .IN3(n28886), .IN4(n27181), .Q(
        n27155) );
  NAND4X0 U31183 ( .IN1(n27158), .IN2(n27157), .IN3(n27156), .IN4(n27155), 
        .QN(s4_addr_o[26]) );
  OA22X1 U31184 ( .IN1(n28901), .IN2(n27187), .IN3(n28900), .IN4(n27168), .Q(
        n27162) );
  OA22X1 U31185 ( .IN1(n28898), .IN2(n27188), .IN3(n28896), .IN4(n27182), .Q(
        n27161) );
  OA22X1 U31186 ( .IN1(n28897), .IN2(n27176), .IN3(n28894), .IN4(n27185), .Q(
        n27160) );
  OA22X1 U31187 ( .IN1(n28899), .IN2(n27184), .IN3(n28895), .IN4(n27174), .Q(
        n27159) );
  NAND4X0 U31188 ( .IN1(n27162), .IN2(n27161), .IN3(n27160), .IN4(n27159), 
        .QN(s4_addr_o[27]) );
  OA22X1 U31189 ( .IN1(n28907), .IN2(n27176), .IN3(n28906), .IN4(n27181), .Q(
        n27166) );
  OA22X1 U31190 ( .IN1(n28910), .IN2(n27182), .IN3(n28908), .IN4(n27187), .Q(
        n27165) );
  OA22X1 U31191 ( .IN1(n28913), .IN2(n27188), .IN3(n28912), .IN4(n27185), .Q(
        n27164) );
  OA22X1 U31192 ( .IN1(n28909), .IN2(n27173), .IN3(n28911), .IN4(n27174), .Q(
        n27163) );
  NAND4X0 U31193 ( .IN1(n27166), .IN2(n27165), .IN3(n27164), .IN4(n27163), 
        .QN(s4_addr_o[28]) );
  OA22X1 U31194 ( .IN1(n28921), .IN2(n27188), .IN3(n28920), .IN4(n27167), .Q(
        n27172) );
  OA22X1 U31195 ( .IN1(n28924), .IN2(n27186), .IN3(n28923), .IN4(n27168), .Q(
        n27171) );
  OA22X1 U31196 ( .IN1(n28926), .IN2(n27184), .IN3(n28922), .IN4(n27183), .Q(
        n27170) );
  OA22X1 U31197 ( .IN1(n28925), .IN2(n27185), .IN3(n28919), .IN4(n27175), .Q(
        n27169) );
  NAND4X0 U31198 ( .IN1(n27172), .IN2(n27171), .IN3(n27170), .IN4(n27169), 
        .QN(s4_addr_o[29]) );
  OA22X1 U31199 ( .IN1(n28936), .IN2(n27182), .IN3(n28931), .IN4(n27185), .Q(
        n27180) );
  OA22X1 U31200 ( .IN1(n28932), .IN2(n27173), .IN3(n28939), .IN4(n27181), .Q(
        n27179) );
  OA22X1 U31201 ( .IN1(n28935), .IN2(n27174), .IN3(n28933), .IN4(n27188), .Q(
        n27178) );
  OA22X1 U31202 ( .IN1(n28937), .IN2(n27176), .IN3(n28940), .IN4(n27175), .Q(
        n27177) );
  NAND4X0 U31203 ( .IN1(n27180), .IN2(n27179), .IN3(n27178), .IN4(n27177), 
        .QN(s4_addr_o[30]) );
  OA22X1 U31204 ( .IN1(n28954), .IN2(n27182), .IN3(n28946), .IN4(n27181), .Q(
        n27192) );
  OA22X1 U31205 ( .IN1(n28948), .IN2(n27184), .IN3(n28956), .IN4(n27183), .Q(
        n27191) );
  OA22X1 U31206 ( .IN1(n28952), .IN2(n27186), .IN3(n28950), .IN4(n27185), .Q(
        n27190) );
  OA22X1 U31207 ( .IN1(n28960), .IN2(n27188), .IN3(n28958), .IN4(n27187), .Q(
        n27189) );
  NAND4X0 U31208 ( .IN1(n27192), .IN2(n27191), .IN3(n27190), .IN4(n27189), 
        .QN(s4_addr_o[31]) );
  OA22X1 U31209 ( .IN1(n29273), .IN2(n27194), .IN3(n29349), .IN4(n27193), .Q(
        n27205) );
  OA22X1 U31210 ( .IN1(n29235), .IN2(n27196), .IN3(n29311), .IN4(n27195), .Q(
        n27204) );
  INVX0 U31211 ( .INP(n27197), .ZN(n27199) );
  OA22X1 U31212 ( .IN1(n29254), .IN2(n27199), .IN3(n29292), .IN4(n27198), .Q(
        n27203) );
  OA22X1 U31213 ( .IN1(n29368), .IN2(n27201), .IN3(n29330), .IN4(n27200), .Q(
        n27202) );
  NAND4X0 U31214 ( .IN1(n27205), .IN2(n27204), .IN3(n27203), .IN4(n27202), 
        .QN(s3_stb_o) );
  INVX0 U31215 ( .INP(n29027), .ZN(n27487) );
  INVX0 U31216 ( .INP(n29019), .ZN(n27489) );
  OA22X1 U31217 ( .IN1(n27487), .IN2(n28128), .IN3(n27489), .IN4(n28125), .Q(
        n27209) );
  INVX0 U31218 ( .INP(n29021), .ZN(n27481) );
  INVX0 U31219 ( .INP(n29022), .ZN(n27456) );
  OA22X1 U31220 ( .IN1(n27481), .IN2(n28123), .IN3(n27456), .IN4(n28122), .Q(
        n27208) );
  INVX0 U31221 ( .INP(n29028), .ZN(n27473) );
  INVX0 U31222 ( .INP(n27443), .ZN(n29020) );
  INVX0 U31223 ( .INP(n29020), .ZN(n27491) );
  OA22X1 U31224 ( .IN1(n27473), .IN2(n28126), .IN3(n27491), .IN4(n28121), .Q(
        n27207) );
  OA22X1 U31225 ( .IN1(n27438), .IN2(n28124), .IN3(n27492), .IN4(n28127), .Q(
        n27206) );
  NAND4X0 U31226 ( .IN1(n27209), .IN2(n27208), .IN3(n27207), .IN4(n27206), 
        .QN(s3_we_o) );
  INVX0 U31227 ( .INP(n29030), .ZN(n27486) );
  OA22X1 U31228 ( .IN1(n27486), .IN2(n28134), .IN3(n27456), .IN4(n28138), .Q(
        n27213) );
  INVX0 U31229 ( .INP(n29021), .ZN(n27493) );
  OA22X1 U31230 ( .IN1(n27493), .IN2(n28133), .IN3(n27473), .IN4(n28139), .Q(
        n27212) );
  INVX0 U31231 ( .INP(n29019), .ZN(n27478) );
  OA22X1 U31232 ( .IN1(n27478), .IN2(n28136), .IN3(n27443), .IN4(n28135), .Q(
        n27211) );
  OA22X1 U31233 ( .IN1(n27480), .IN2(n28140), .IN3(n27492), .IN4(n28137), .Q(
        n27210) );
  NAND4X0 U31234 ( .IN1(n27213), .IN2(n27212), .IN3(n27211), .IN4(n27210), 
        .QN(s3_data_o[0]) );
  INVX0 U31235 ( .INP(n29028), .ZN(n27488) );
  OA22X1 U31236 ( .IN1(n27488), .IN2(n28145), .IN3(n27443), .IN4(n28147), .Q(
        n27217) );
  OA22X1 U31237 ( .IN1(n27480), .IN2(n28146), .IN3(n27492), .IN4(n28151), .Q(
        n27216) );
  OA22X1 U31238 ( .IN1(n27481), .IN2(n28148), .IN3(n27489), .IN4(n28152), .Q(
        n27215) );
  OA22X1 U31239 ( .IN1(n27486), .IN2(n28150), .IN3(n27456), .IN4(n28149), .Q(
        n27214) );
  NAND4X0 U31240 ( .IN1(n27217), .IN2(n27216), .IN3(n27215), .IN4(n27214), 
        .QN(s3_data_o[1]) );
  OA22X1 U31241 ( .IN1(n27480), .IN2(n28164), .IN3(n27456), .IN4(n28158), .Q(
        n27221) );
  OA22X1 U31242 ( .IN1(n27493), .IN2(n28163), .IN3(n27492), .IN4(n28157), .Q(
        n27220) );
  OA22X1 U31243 ( .IN1(n27473), .IN2(n28159), .IN3(n27489), .IN4(n28162), .Q(
        n27219) );
  OA22X1 U31244 ( .IN1(n27438), .IN2(n28160), .IN3(n27443), .IN4(n28161), .Q(
        n27218) );
  NAND4X0 U31245 ( .IN1(n27221), .IN2(n27220), .IN3(n27219), .IN4(n27218), 
        .QN(s3_data_o[2]) );
  INVX0 U31246 ( .INP(n27492), .ZN(n29029) );
  INVX0 U31247 ( .INP(n29029), .ZN(n27479) );
  OA22X1 U31248 ( .IN1(n27479), .IN2(n28169), .IN3(n27443), .IN4(n28173), .Q(
        n27225) );
  OA22X1 U31249 ( .IN1(n27486), .IN2(n28172), .IN3(n27456), .IN4(n28171), .Q(
        n27224) );
  OA22X1 U31250 ( .IN1(n27481), .IN2(n28176), .IN3(n27489), .IN4(n28175), .Q(
        n27223) );
  OA22X1 U31251 ( .IN1(n27480), .IN2(n28174), .IN3(n27473), .IN4(n28170), .Q(
        n27222) );
  NAND4X0 U31252 ( .IN1(n27225), .IN2(n27224), .IN3(n27223), .IN4(n27222), 
        .QN(s3_data_o[3]) );
  OA22X1 U31253 ( .IN1(n27493), .IN2(n28186), .IN3(n27443), .IN4(n28181), .Q(
        n27229) );
  OA22X1 U31254 ( .IN1(n27487), .IN2(n28184), .IN3(n27489), .IN4(n28183), .Q(
        n27228) );
  OA22X1 U31255 ( .IN1(n27486), .IN2(n28182), .IN3(n27456), .IN4(n28185), .Q(
        n27227) );
  OA22X1 U31256 ( .IN1(n27488), .IN2(n28188), .IN3(n27492), .IN4(n28187), .Q(
        n27226) );
  NAND4X0 U31257 ( .IN1(n27229), .IN2(n27228), .IN3(n27227), .IN4(n27226), 
        .QN(s3_data_o[4]) );
  OA22X1 U31258 ( .IN1(n27480), .IN2(n28200), .IN3(n27489), .IN4(n28197), .Q(
        n27233) );
  OA22X1 U31259 ( .IN1(n27438), .IN2(n28196), .IN3(n27456), .IN4(n28198), .Q(
        n27232) );
  OA22X1 U31260 ( .IN1(n27473), .IN2(n28193), .IN3(n27492), .IN4(n28195), .Q(
        n27231) );
  OA22X1 U31261 ( .IN1(n27481), .IN2(n28194), .IN3(n27443), .IN4(n28199), .Q(
        n27230) );
  NAND4X0 U31262 ( .IN1(n27233), .IN2(n27232), .IN3(n27231), .IN4(n27230), 
        .QN(s3_data_o[5]) );
  OA22X1 U31263 ( .IN1(n27488), .IN2(n28212), .IN3(n27456), .IN4(n28211), .Q(
        n27237) );
  OA22X1 U31264 ( .IN1(n27478), .IN2(n28205), .IN3(n27492), .IN4(n28210), .Q(
        n27236) );
  OA22X1 U31265 ( .IN1(n27486), .IN2(n28208), .IN3(n27443), .IN4(n28209), .Q(
        n27235) );
  OA22X1 U31266 ( .IN1(n27487), .IN2(n28207), .IN3(n27481), .IN4(n28206), .Q(
        n27234) );
  NAND4X0 U31267 ( .IN1(n27237), .IN2(n27236), .IN3(n27235), .IN4(n27234), 
        .QN(s3_data_o[6]) );
  OA22X1 U31268 ( .IN1(n27481), .IN2(n28224), .IN3(n27491), .IN4(n28221), .Q(
        n27241) );
  OA22X1 U31269 ( .IN1(n27489), .IN2(n28223), .IN3(n27492), .IN4(n28222), .Q(
        n27240) );
  OA22X1 U31270 ( .IN1(n27438), .IN2(n28220), .IN3(n27456), .IN4(n28217), .Q(
        n27239) );
  OA22X1 U31271 ( .IN1(n27480), .IN2(n28219), .IN3(n27473), .IN4(n28218), .Q(
        n27238) );
  NAND4X0 U31272 ( .IN1(n27241), .IN2(n27240), .IN3(n27239), .IN4(n27238), 
        .QN(s3_data_o[7]) );
  OA22X1 U31273 ( .IN1(n27487), .IN2(n28232), .IN3(n27491), .IN4(n28235), .Q(
        n27245) );
  INVX0 U31274 ( .INP(n29022), .ZN(n27490) );
  OA22X1 U31275 ( .IN1(n27490), .IN2(n28236), .IN3(n27489), .IN4(n28229), .Q(
        n27244) );
  OA22X1 U31276 ( .IN1(n27486), .IN2(n28230), .IN3(n27481), .IN4(n28231), .Q(
        n27243) );
  OA22X1 U31277 ( .IN1(n27473), .IN2(n28234), .IN3(n27492), .IN4(n28233), .Q(
        n27242) );
  NAND4X0 U31278 ( .IN1(n27245), .IN2(n27244), .IN3(n27243), .IN4(n27242), 
        .QN(s3_data_o[8]) );
  OA22X1 U31279 ( .IN1(n27478), .IN2(n28245), .IN3(n27491), .IN4(n28247), .Q(
        n27249) );
  OA22X1 U31280 ( .IN1(n27438), .IN2(n28242), .IN3(n27456), .IN4(n28241), .Q(
        n27248) );
  OA22X1 U31281 ( .IN1(n27493), .IN2(n28246), .IN3(n27479), .IN4(n28243), .Q(
        n27247) );
  OA22X1 U31282 ( .IN1(n27480), .IN2(n28244), .IN3(n27473), .IN4(n28248), .Q(
        n27246) );
  NAND4X0 U31283 ( .IN1(n27249), .IN2(n27248), .IN3(n27247), .IN4(n27246), 
        .QN(s3_data_o[9]) );
  OA22X1 U31284 ( .IN1(n27488), .IN2(n28256), .IN3(n27479), .IN4(n28253), .Q(
        n27253) );
  OA22X1 U31285 ( .IN1(n27456), .IN2(n28254), .IN3(n27489), .IN4(n28255), .Q(
        n27252) );
  OA22X1 U31286 ( .IN1(n27486), .IN2(n28258), .IN3(n27491), .IN4(n28259), .Q(
        n27251) );
  OA22X1 U31287 ( .IN1(n27487), .IN2(n28257), .IN3(n27481), .IN4(n28260), .Q(
        n27250) );
  NAND4X0 U31288 ( .IN1(n27253), .IN2(n27252), .IN3(n27251), .IN4(n27250), 
        .QN(s3_data_o[10]) );
  OA22X1 U31289 ( .IN1(n27490), .IN2(n28268), .IN3(n27491), .IN4(n28269), .Q(
        n27257) );
  OA22X1 U31290 ( .IN1(n27481), .IN2(n28265), .IN3(n27473), .IN4(n28271), .Q(
        n27256) );
  OA22X1 U31291 ( .IN1(n27480), .IN2(n28272), .IN3(n27479), .IN4(n28267), .Q(
        n27255) );
  OA22X1 U31292 ( .IN1(n27438), .IN2(n28266), .IN3(n27489), .IN4(n28270), .Q(
        n27254) );
  NAND4X0 U31293 ( .IN1(n27257), .IN2(n27256), .IN3(n27255), .IN4(n27254), 
        .QN(s3_data_o[11]) );
  OA22X1 U31294 ( .IN1(n27487), .IN2(n28278), .IN3(n27489), .IN4(n28281), .Q(
        n27261) );
  OA22X1 U31295 ( .IN1(n27493), .IN2(n28280), .IN3(n27473), .IN4(n28282), .Q(
        n27260) );
  OA22X1 U31296 ( .IN1(n27479), .IN2(n28279), .IN3(n27491), .IN4(n28277), .Q(
        n27259) );
  OA22X1 U31297 ( .IN1(n27486), .IN2(n28284), .IN3(n27456), .IN4(n28283), .Q(
        n27258) );
  NAND4X0 U31298 ( .IN1(n27261), .IN2(n27260), .IN3(n27259), .IN4(n27258), 
        .QN(s3_data_o[12]) );
  OA22X1 U31299 ( .IN1(n27488), .IN2(n28292), .IN3(n27491), .IN4(n28295), .Q(
        n27265) );
  OA22X1 U31300 ( .IN1(n27481), .IN2(n28296), .IN3(n27489), .IN4(n28293), .Q(
        n27264) );
  OA22X1 U31301 ( .IN1(n27456), .IN2(n28289), .IN3(n27479), .IN4(n28291), .Q(
        n27263) );
  OA22X1 U31302 ( .IN1(n27438), .IN2(n28290), .IN3(n27480), .IN4(n28294), .Q(
        n27262) );
  NAND4X0 U31303 ( .IN1(n27265), .IN2(n27264), .IN3(n27263), .IN4(n27262), 
        .QN(s3_data_o[13]) );
  OA22X1 U31304 ( .IN1(n27480), .IN2(n28304), .IN3(n27491), .IN4(n28303), .Q(
        n27269) );
  OA22X1 U31305 ( .IN1(n27493), .IN2(n28308), .IN3(n27473), .IN4(n28305), .Q(
        n27268) );
  OA22X1 U31306 ( .IN1(n27486), .IN2(n28306), .IN3(n27479), .IN4(n28301), .Q(
        n27267) );
  OA22X1 U31307 ( .IN1(n27490), .IN2(n28307), .IN3(n27489), .IN4(n28302), .Q(
        n27266) );
  NAND4X0 U31308 ( .IN1(n27269), .IN2(n27268), .IN3(n27267), .IN4(n27266), 
        .QN(s3_data_o[14]) );
  OA22X1 U31309 ( .IN1(n27438), .IN2(n28316), .IN3(n27491), .IN4(n28319), .Q(
        n27273) );
  OA22X1 U31310 ( .IN1(n27456), .IN2(n28320), .IN3(n27479), .IN4(n28317), .Q(
        n27272) );
  OA22X1 U31311 ( .IN1(n27488), .IN2(n28313), .IN3(n27489), .IN4(n28318), .Q(
        n27271) );
  OA22X1 U31312 ( .IN1(n27487), .IN2(n28315), .IN3(n27481), .IN4(n28314), .Q(
        n27270) );
  NAND4X0 U31313 ( .IN1(n27273), .IN2(n27272), .IN3(n27271), .IN4(n27270), 
        .QN(s3_data_o[15]) );
  OA22X1 U31314 ( .IN1(n27480), .IN2(n28332), .IN3(n27479), .IN4(n28328), .Q(
        n27277) );
  OA22X1 U31315 ( .IN1(n27478), .IN2(n28325), .IN3(n27491), .IN4(n28327), .Q(
        n27276) );
  OA22X1 U31316 ( .IN1(n27438), .IN2(n28330), .IN3(n27481), .IN4(n28331), .Q(
        n27275) );
  OA22X1 U31317 ( .IN1(n27473), .IN2(n28326), .IN3(n27456), .IN4(n28329), .Q(
        n27274) );
  NAND4X0 U31318 ( .IN1(n27277), .IN2(n27276), .IN3(n27275), .IN4(n27274), 
        .QN(s3_data_o[16]) );
  OA22X1 U31319 ( .IN1(n27486), .IN2(n28340), .IN3(n27481), .IN4(n28342), .Q(
        n27281) );
  OA22X1 U31320 ( .IN1(n27488), .IN2(n28338), .IN3(n27479), .IN4(n28343), .Q(
        n27280) );
  OA22X1 U31321 ( .IN1(n27490), .IN2(n28337), .IN3(n27489), .IN4(n28339), .Q(
        n27279) );
  OA22X1 U31322 ( .IN1(n27487), .IN2(n28344), .IN3(n27491), .IN4(n28341), .Q(
        n27278) );
  NAND4X0 U31323 ( .IN1(n27281), .IN2(n27280), .IN3(n27279), .IN4(n27278), 
        .QN(s3_data_o[17]) );
  OA22X1 U31324 ( .IN1(n27490), .IN2(n28354), .IN3(n27479), .IN4(n28351), .Q(
        n27285) );
  OA22X1 U31325 ( .IN1(n27438), .IN2(n28352), .IN3(n27489), .IN4(n28349), .Q(
        n27284) );
  OA22X1 U31326 ( .IN1(n27493), .IN2(n28350), .IN3(n27473), .IN4(n28355), .Q(
        n27283) );
  OA22X1 U31327 ( .IN1(n27480), .IN2(n28356), .IN3(n27491), .IN4(n28353), .Q(
        n27282) );
  NAND4X0 U31328 ( .IN1(n27285), .IN2(n27284), .IN3(n27283), .IN4(n27282), 
        .QN(s3_data_o[18]) );
  OA22X1 U31329 ( .IN1(n27487), .IN2(n28364), .IN3(n27479), .IN4(n28368), .Q(
        n27289) );
  OA22X1 U31330 ( .IN1(n27438), .IN2(n28366), .IN3(n27473), .IN4(n28363), .Q(
        n27288) );
  OA22X1 U31331 ( .IN1(n27493), .IN2(n28362), .IN3(n27489), .IN4(n28361), .Q(
        n27287) );
  OA22X1 U31332 ( .IN1(n27490), .IN2(n28365), .IN3(n27491), .IN4(n28367), .Q(
        n27286) );
  NAND4X0 U31333 ( .IN1(n27289), .IN2(n27288), .IN3(n27287), .IN4(n27286), 
        .QN(s3_data_o[19]) );
  OA22X1 U31334 ( .IN1(n27481), .IN2(n28374), .IN3(n27456), .IN4(n28376), .Q(
        n27293) );
  OA22X1 U31335 ( .IN1(n27438), .IN2(n28378), .IN3(n27491), .IN4(n28375), .Q(
        n27292) );
  OA22X1 U31336 ( .IN1(n27487), .IN2(n28377), .IN3(n27473), .IN4(n28373), .Q(
        n27291) );
  OA22X1 U31337 ( .IN1(n27489), .IN2(n28380), .IN3(n27479), .IN4(n28379), .Q(
        n27290) );
  NAND4X0 U31338 ( .IN1(n27293), .IN2(n27292), .IN3(n27291), .IN4(n27290), 
        .QN(s3_data_o[20]) );
  OA22X1 U31339 ( .IN1(n27481), .IN2(n28390), .IN3(n27479), .IN4(n28389), .Q(
        n27297) );
  OA22X1 U31340 ( .IN1(n27487), .IN2(n28386), .IN3(n27489), .IN4(n28385), .Q(
        n27296) );
  OA22X1 U31341 ( .IN1(n27438), .IN2(n28392), .IN3(n27491), .IN4(n28391), .Q(
        n27295) );
  OA22X1 U31342 ( .IN1(n27488), .IN2(n28388), .IN3(n27456), .IN4(n28387), .Q(
        n27294) );
  NAND4X0 U31343 ( .IN1(n27297), .IN2(n27296), .IN3(n27295), .IN4(n27294), 
        .QN(s3_data_o[21]) );
  OA22X1 U31344 ( .IN1(n27488), .IN2(n28403), .IN3(n27491), .IN4(n28397), .Q(
        n27301) );
  OA22X1 U31345 ( .IN1(n27481), .IN2(n28404), .IN3(n27489), .IN4(n28399), .Q(
        n27300) );
  OA22X1 U31346 ( .IN1(n27487), .IN2(n28402), .IN3(n27479), .IN4(n28401), .Q(
        n27299) );
  OA22X1 U31347 ( .IN1(n27438), .IN2(n28400), .IN3(n27456), .IN4(n28398), .Q(
        n27298) );
  NAND4X0 U31348 ( .IN1(n27301), .IN2(n27300), .IN3(n27299), .IN4(n27298), 
        .QN(s3_data_o[22]) );
  OA22X1 U31349 ( .IN1(n27487), .IN2(n28415), .IN3(n27481), .IN4(n28414), .Q(
        n27305) );
  OA22X1 U31350 ( .IN1(n27438), .IN2(n28416), .IN3(n27456), .IN4(n28410), .Q(
        n27304) );
  OA22X1 U31351 ( .IN1(n27488), .IN2(n28413), .IN3(n27443), .IN4(n28411), .Q(
        n27303) );
  OA22X1 U31352 ( .IN1(n27478), .IN2(n28412), .IN3(n27479), .IN4(n28409), .Q(
        n27302) );
  NAND4X0 U31353 ( .IN1(n27305), .IN2(n27304), .IN3(n27303), .IN4(n27302), 
        .QN(s3_data_o[23]) );
  OA22X1 U31354 ( .IN1(n27487), .IN2(n28424), .IN3(n27493), .IN4(n28422), .Q(
        n27309) );
  OA22X1 U31355 ( .IN1(n27478), .IN2(n28428), .IN3(n27479), .IN4(n28427), .Q(
        n27308) );
  OA22X1 U31356 ( .IN1(n27438), .IN2(n28426), .IN3(n27456), .IN4(n28425), .Q(
        n27307) );
  OA22X1 U31357 ( .IN1(n27488), .IN2(n28421), .IN3(n27443), .IN4(n28423), .Q(
        n27306) );
  NAND4X0 U31358 ( .IN1(n27309), .IN2(n27308), .IN3(n27307), .IN4(n27306), 
        .QN(s3_data_o[24]) );
  OA22X1 U31359 ( .IN1(n27479), .IN2(n28436), .IN3(n27443), .IN4(n28435), .Q(
        n27313) );
  OA22X1 U31360 ( .IN1(n27438), .IN2(n28438), .IN3(n27456), .IN4(n28433), .Q(
        n27312) );
  OA22X1 U31361 ( .IN1(n27487), .IN2(n28440), .IN3(n27473), .IN4(n28439), .Q(
        n27311) );
  OA22X1 U31362 ( .IN1(n27493), .IN2(n28434), .IN3(n27489), .IN4(n28437), .Q(
        n27310) );
  NAND4X0 U31363 ( .IN1(n27313), .IN2(n27312), .IN3(n27311), .IN4(n27310), 
        .QN(s3_data_o[25]) );
  OA22X1 U31364 ( .IN1(n27487), .IN2(n28451), .IN3(n27481), .IN4(n28450), .Q(
        n27317) );
  OA22X1 U31365 ( .IN1(n27488), .IN2(n28446), .IN3(n27443), .IN4(n28445), .Q(
        n27316) );
  OA22X1 U31366 ( .IN1(n27489), .IN2(n28448), .IN3(n27479), .IN4(n28447), .Q(
        n27315) );
  OA22X1 U31367 ( .IN1(n27438), .IN2(n28452), .IN3(n27456), .IN4(n28449), .Q(
        n27314) );
  NAND4X0 U31368 ( .IN1(n27317), .IN2(n27316), .IN3(n27315), .IN4(n27314), 
        .QN(s3_data_o[26]) );
  OA22X1 U31369 ( .IN1(n27487), .IN2(n28461), .IN3(n27481), .IN4(n28464), .Q(
        n27321) );
  OA22X1 U31370 ( .IN1(n27488), .IN2(n28458), .IN3(n27443), .IN4(n28459), .Q(
        n27320) );
  OA22X1 U31371 ( .IN1(n27478), .IN2(n28463), .IN3(n27492), .IN4(n28460), .Q(
        n27319) );
  OA22X1 U31372 ( .IN1(n27438), .IN2(n28462), .IN3(n27490), .IN4(n28457), .Q(
        n27318) );
  NAND4X0 U31373 ( .IN1(n27321), .IN2(n27320), .IN3(n27319), .IN4(n27318), 
        .QN(s3_data_o[27]) );
  OA22X1 U31374 ( .IN1(n27487), .IN2(n28476), .IN3(n27492), .IN4(n28469), .Q(
        n27325) );
  OA22X1 U31375 ( .IN1(n27481), .IN2(n28472), .IN3(n27473), .IN4(n28470), .Q(
        n27324) );
  OA22X1 U31376 ( .IN1(n27490), .IN2(n28471), .IN3(n27489), .IN4(n28475), .Q(
        n27323) );
  OA22X1 U31377 ( .IN1(n27438), .IN2(n28474), .IN3(n27443), .IN4(n28473), .Q(
        n27322) );
  NAND4X0 U31378 ( .IN1(n27325), .IN2(n27324), .IN3(n27323), .IN4(n27322), 
        .QN(s3_data_o[28]) );
  OA22X1 U31379 ( .IN1(n27490), .IN2(n28487), .IN3(n27478), .IN4(n28483), .Q(
        n27329) );
  OA22X1 U31380 ( .IN1(n27438), .IN2(n28484), .IN3(n27443), .IN4(n28481), .Q(
        n27328) );
  OA22X1 U31381 ( .IN1(n27481), .IN2(n28488), .IN3(n27492), .IN4(n28485), .Q(
        n27327) );
  OA22X1 U31382 ( .IN1(n27487), .IN2(n28482), .IN3(n27488), .IN4(n28486), .Q(
        n27326) );
  NAND4X0 U31383 ( .IN1(n27329), .IN2(n27328), .IN3(n27327), .IN4(n27326), 
        .QN(s3_data_o[29]) );
  OA22X1 U31384 ( .IN1(n27473), .IN2(n28496), .IN3(n27443), .IN4(n28499), .Q(
        n27333) );
  OA22X1 U31385 ( .IN1(n27438), .IN2(n28494), .IN3(n27492), .IN4(n28500), .Q(
        n27332) );
  OA22X1 U31386 ( .IN1(n27487), .IN2(n28498), .IN3(n27489), .IN4(n28495), .Q(
        n27331) );
  OA22X1 U31387 ( .IN1(n27493), .IN2(n28497), .IN3(n27456), .IN4(n28493), .Q(
        n27330) );
  NAND4X0 U31388 ( .IN1(n27333), .IN2(n27332), .IN3(n27331), .IN4(n27330), 
        .QN(s3_data_o[30]) );
  OA22X1 U31389 ( .IN1(n27490), .IN2(n28512), .IN3(n27443), .IN4(n28507), .Q(
        n27337) );
  OA22X1 U31390 ( .IN1(n27438), .IN2(n28510), .IN3(n27481), .IN4(n28506), .Q(
        n27336) );
  OA22X1 U31391 ( .IN1(n27487), .IN2(n28509), .IN3(n27489), .IN4(n28508), .Q(
        n27335) );
  OA22X1 U31392 ( .IN1(n27473), .IN2(n28505), .IN3(n27492), .IN4(n28511), .Q(
        n27334) );
  NAND4X0 U31393 ( .IN1(n27337), .IN2(n27336), .IN3(n27335), .IN4(n27334), 
        .QN(s3_data_o[31]) );
  OA22X1 U31394 ( .IN1(n27493), .IN2(n28522), .IN3(n27492), .IN4(n28521), .Q(
        n27341) );
  OA22X1 U31395 ( .IN1(n27478), .IN2(n28520), .IN3(n27443), .IN4(n28519), .Q(
        n27340) );
  OA22X1 U31396 ( .IN1(n27486), .IN2(n28518), .IN3(n27490), .IN4(n28523), .Q(
        n27339) );
  OA22X1 U31397 ( .IN1(n27487), .IN2(n28517), .IN3(n27473), .IN4(n28524), .Q(
        n27338) );
  NAND4X0 U31398 ( .IN1(n27341), .IN2(n27340), .IN3(n27339), .IN4(n27338), 
        .QN(s3_sel_o[0]) );
  OA22X1 U31399 ( .IN1(n27473), .IN2(n28536), .IN3(n27456), .IN4(n28535), .Q(
        n27345) );
  OA22X1 U31400 ( .IN1(n27481), .IN2(n28530), .IN3(n27443), .IN4(n28529), .Q(
        n27344) );
  OA22X1 U31401 ( .IN1(n27478), .IN2(n28533), .IN3(n27492), .IN4(n28531), .Q(
        n27343) );
  OA22X1 U31402 ( .IN1(n27486), .IN2(n28534), .IN3(n27480), .IN4(n28532), .Q(
        n27342) );
  NAND4X0 U31403 ( .IN1(n27345), .IN2(n27344), .IN3(n27343), .IN4(n27342), 
        .QN(s3_sel_o[1]) );
  OA22X1 U31404 ( .IN1(n27487), .IN2(n28546), .IN3(n27443), .IN4(n28541), .Q(
        n27349) );
  OA22X1 U31405 ( .IN1(n27486), .IN2(n28544), .IN3(n27473), .IN4(n28548), .Q(
        n27348) );
  OA22X1 U31406 ( .IN1(n27493), .IN2(n28543), .IN3(n27478), .IN4(n28542), .Q(
        n27347) );
  OA22X1 U31407 ( .IN1(n27456), .IN2(n28547), .IN3(n27492), .IN4(n28545), .Q(
        n27346) );
  NAND4X0 U31408 ( .IN1(n27349), .IN2(n27348), .IN3(n27347), .IN4(n27346), 
        .QN(s3_sel_o[2]) );
  OA22X1 U31409 ( .IN1(n27478), .IN2(n28560), .IN3(n27443), .IN4(n28555), .Q(
        n27353) );
  OA22X1 U31410 ( .IN1(n27480), .IN2(n28554), .IN3(n27490), .IN4(n28556), .Q(
        n27352) );
  OA22X1 U31411 ( .IN1(n27486), .IN2(n28558), .IN3(n27492), .IN4(n28559), .Q(
        n27351) );
  OA22X1 U31412 ( .IN1(n27493), .IN2(n28553), .IN3(n27488), .IN4(n28557), .Q(
        n27350) );
  NAND4X0 U31413 ( .IN1(n27353), .IN2(n27352), .IN3(n27351), .IN4(n27350), 
        .QN(s3_sel_o[3]) );
  OA22X1 U31414 ( .IN1(n27478), .IN2(n28567), .IN3(n27492), .IN4(n28565), .Q(
        n27357) );
  OA22X1 U31415 ( .IN1(n27493), .IN2(n28571), .IN3(n27488), .IN4(n28566), .Q(
        n27356) );
  OA22X1 U31416 ( .IN1(n27486), .IN2(n28572), .IN3(n27443), .IN4(n28569), .Q(
        n27355) );
  OA22X1 U31417 ( .IN1(n27480), .IN2(n28570), .IN3(n27490), .IN4(n28568), .Q(
        n27354) );
  NAND4X0 U31418 ( .IN1(n27357), .IN2(n27356), .IN3(n27355), .IN4(n27354), 
        .QN(s3_addr_o[0]) );
  OA22X1 U31419 ( .IN1(n27480), .IN2(n28578), .IN3(n27478), .IN4(n28584), .Q(
        n27361) );
  OA22X1 U31420 ( .IN1(n27493), .IN2(n28582), .IN3(n27443), .IN4(n28583), .Q(
        n27360) );
  OA22X1 U31421 ( .IN1(n27473), .IN2(n28581), .IN3(n27490), .IN4(n28579), .Q(
        n27359) );
  OA22X1 U31422 ( .IN1(n27438), .IN2(n28580), .IN3(n27492), .IN4(n28577), .Q(
        n27358) );
  NAND4X0 U31423 ( .IN1(n27361), .IN2(n27360), .IN3(n27359), .IN4(n27358), 
        .QN(s3_addr_o[1]) );
  OA22X1 U31424 ( .IN1(n28591), .IN2(n27486), .IN3(n28589), .IN4(n27480), .Q(
        n27365) );
  OA22X1 U31425 ( .IN1(n28592), .IN2(n27473), .IN3(n28593), .IN4(n27478), .Q(
        n27364) );
  OA22X1 U31426 ( .IN1(n28594), .IN2(n27493), .IN3(n28595), .IN4(n27492), .Q(
        n27363) );
  OA22X1 U31427 ( .IN1(n28596), .IN2(n27491), .IN3(n28590), .IN4(n27456), .Q(
        n27362) );
  NAND4X0 U31428 ( .IN1(n27365), .IN2(n27364), .IN3(n27363), .IN4(n27362), 
        .QN(s3_addr_o[2]) );
  OA22X1 U31429 ( .IN1(n28608), .IN2(n27491), .IN3(n28607), .IN4(n27488), .Q(
        n27369) );
  OA22X1 U31430 ( .IN1(n28602), .IN2(n27489), .IN3(n28605), .IN4(n27480), .Q(
        n27368) );
  OA22X1 U31431 ( .IN1(n28606), .IN2(n27456), .IN3(n28601), .IN4(n27486), .Q(
        n27367) );
  OA22X1 U31432 ( .IN1(n28604), .IN2(n27481), .IN3(n28603), .IN4(n27492), .Q(
        n27366) );
  NAND4X0 U31433 ( .IN1(n27369), .IN2(n27368), .IN3(n27367), .IN4(n27366), 
        .QN(s3_addr_o[3]) );
  OA22X1 U31434 ( .IN1(n28618), .IN2(n27488), .IN3(n28614), .IN4(n27478), .Q(
        n27373) );
  OA22X1 U31435 ( .IN1(n28620), .IN2(n27479), .IN3(n28615), .IN4(n27456), .Q(
        n27372) );
  OA22X1 U31436 ( .IN1(n28616), .IN2(n27487), .IN3(n28619), .IN4(n27491), .Q(
        n27371) );
  OA22X1 U31437 ( .IN1(n28617), .IN2(n27438), .IN3(n28613), .IN4(n27481), .Q(
        n27370) );
  NAND4X0 U31438 ( .IN1(n27373), .IN2(n27372), .IN3(n27371), .IN4(n27370), 
        .QN(s3_addr_o[4]) );
  OA22X1 U31439 ( .IN1(n28627), .IN2(n27478), .IN3(n28625), .IN4(n27491), .Q(
        n27377) );
  OA22X1 U31440 ( .IN1(n28632), .IN2(n27493), .IN3(n28626), .IN4(n27488), .Q(
        n27376) );
  OA22X1 U31441 ( .IN1(n28630), .IN2(n27487), .IN3(n28629), .IN4(n27486), .Q(
        n27375) );
  OA22X1 U31442 ( .IN1(n28628), .IN2(n27479), .IN3(n28631), .IN4(n27490), .Q(
        n27374) );
  NAND4X0 U31443 ( .IN1(n27377), .IN2(n27376), .IN3(n27375), .IN4(n27374), 
        .QN(s3_addr_o[5]) );
  OA22X1 U31444 ( .IN1(n27438), .IN2(n28642), .IN3(n27478), .IN4(n28637), .Q(
        n27381) );
  OA22X1 U31445 ( .IN1(n27493), .IN2(n28644), .IN3(n27473), .IN4(n28643), .Q(
        n27380) );
  OA22X1 U31446 ( .IN1(n27480), .IN2(n28640), .IN3(n27492), .IN4(n28641), .Q(
        n27379) );
  OA22X1 U31447 ( .IN1(n27490), .IN2(n28638), .IN3(n27443), .IN4(n28639), .Q(
        n27378) );
  NAND4X0 U31448 ( .IN1(n27381), .IN2(n27380), .IN3(n27379), .IN4(n27378), 
        .QN(s3_addr_o[6]) );
  OA22X1 U31449 ( .IN1(n27473), .IN2(n28653), .IN3(n27443), .IN4(n28655), .Q(
        n27385) );
  OA22X1 U31450 ( .IN1(n27438), .IN2(n28654), .IN3(n27481), .IN4(n28656), .Q(
        n27384) );
  OA22X1 U31451 ( .IN1(n27480), .IN2(n28652), .IN3(n27489), .IN4(n28649), .Q(
        n27383) );
  OA22X1 U31452 ( .IN1(n27490), .IN2(n28650), .IN3(n27492), .IN4(n28651), .Q(
        n27382) );
  NAND4X0 U31453 ( .IN1(n27385), .IN2(n27384), .IN3(n27383), .IN4(n27382), 
        .QN(s3_addr_o[7]) );
  OA22X1 U31454 ( .IN1(n27487), .IN2(n28663), .IN3(n27478), .IN4(n28662), .Q(
        n27389) );
  OA22X1 U31455 ( .IN1(n27486), .IN2(n28664), .IN3(n27443), .IN4(n28667), .Q(
        n27388) );
  OA22X1 U31456 ( .IN1(n27493), .IN2(n28666), .IN3(n27490), .IN4(n28668), .Q(
        n27387) );
  OA22X1 U31457 ( .IN1(n27488), .IN2(n28665), .IN3(n27492), .IN4(n28661), .Q(
        n27386) );
  NAND4X0 U31458 ( .IN1(n27389), .IN2(n27388), .IN3(n27387), .IN4(n27386), 
        .QN(s3_addr_o[8]) );
  OA22X1 U31459 ( .IN1(n27493), .IN2(n28674), .IN3(n27478), .IN4(n28678), .Q(
        n27393) );
  OA22X1 U31460 ( .IN1(n27479), .IN2(n28675), .IN3(n27443), .IN4(n28677), .Q(
        n27392) );
  OA22X1 U31461 ( .IN1(n27486), .IN2(n28680), .IN3(n27480), .IN4(n28679), .Q(
        n27391) );
  OA22X1 U31462 ( .IN1(n27488), .IN2(n28676), .IN3(n27456), .IN4(n28673), .Q(
        n27390) );
  NAND4X0 U31463 ( .IN1(n27393), .IN2(n27392), .IN3(n27391), .IN4(n27390), 
        .QN(s3_addr_o[9]) );
  OA22X1 U31464 ( .IN1(n27438), .IN2(n28692), .IN3(n27481), .IN4(n28688), .Q(
        n27397) );
  OA22X1 U31465 ( .IN1(n27490), .IN2(n28685), .IN3(n27443), .IN4(n28689), .Q(
        n27396) );
  OA22X1 U31466 ( .IN1(n27480), .IN2(n28686), .IN3(n27489), .IN4(n28691), .Q(
        n27395) );
  OA22X1 U31467 ( .IN1(n27473), .IN2(n28687), .IN3(n27492), .IN4(n28690), .Q(
        n27394) );
  NAND4X0 U31468 ( .IN1(n27397), .IN2(n27396), .IN3(n27395), .IN4(n27394), 
        .QN(s3_addr_o[10]) );
  OA22X1 U31469 ( .IN1(n27493), .IN2(n28697), .IN3(n27478), .IN4(n28703), .Q(
        n27401) );
  OA22X1 U31470 ( .IN1(n27473), .IN2(n28704), .IN3(n27490), .IN4(n28701), .Q(
        n27400) );
  OA22X1 U31471 ( .IN1(n27480), .IN2(n28698), .IN3(n27443), .IN4(n28699), .Q(
        n27399) );
  OA22X1 U31472 ( .IN1(n27486), .IN2(n28702), .IN3(n27492), .IN4(n28700), .Q(
        n27398) );
  NAND4X0 U31473 ( .IN1(n27401), .IN2(n27400), .IN3(n27399), .IN4(n27398), 
        .QN(s3_addr_o[11]) );
  OA22X1 U31474 ( .IN1(n27488), .IN2(n28716), .IN3(n27490), .IN4(n28709), .Q(
        n27405) );
  OA22X1 U31475 ( .IN1(n27480), .IN2(n28710), .IN3(n27443), .IN4(n28713), .Q(
        n27404) );
  OA22X1 U31476 ( .IN1(n27493), .IN2(n28712), .IN3(n27489), .IN4(n28715), .Q(
        n27403) );
  OA22X1 U31477 ( .IN1(n27486), .IN2(n28714), .IN3(n27492), .IN4(n28711), .Q(
        n27402) );
  NAND4X0 U31478 ( .IN1(n27405), .IN2(n27404), .IN3(n27403), .IN4(n27402), 
        .QN(s3_addr_o[12]) );
  OA22X1 U31479 ( .IN1(n27487), .IN2(n28728), .IN3(n27443), .IN4(n28727), .Q(
        n27409) );
  OA22X1 U31480 ( .IN1(n27490), .IN2(n28723), .IN3(n27492), .IN4(n28725), .Q(
        n27408) );
  OA22X1 U31481 ( .IN1(n27438), .IN2(n28722), .IN3(n27481), .IN4(n28726), .Q(
        n27407) );
  OA22X1 U31482 ( .IN1(n27473), .IN2(n28724), .IN3(n27489), .IN4(n28721), .Q(
        n27406) );
  NAND4X0 U31483 ( .IN1(n27409), .IN2(n27408), .IN3(n27407), .IN4(n27406), 
        .QN(s3_addr_o[13]) );
  OA22X1 U31484 ( .IN1(n27487), .IN2(n28738), .IN3(n27478), .IN4(n28737), .Q(
        n27413) );
  OA22X1 U31485 ( .IN1(n27493), .IN2(n28736), .IN3(n27492), .IN4(n28733), .Q(
        n27412) );
  OA22X1 U31486 ( .IN1(n27488), .IN2(n28735), .IN3(n27443), .IN4(n28739), .Q(
        n27411) );
  OA22X1 U31487 ( .IN1(n27438), .IN2(n28734), .IN3(n27456), .IN4(n28740), .Q(
        n27410) );
  NAND4X0 U31488 ( .IN1(n27413), .IN2(n27412), .IN3(n27411), .IN4(n27410), 
        .QN(s3_addr_o[14]) );
  OA22X1 U31489 ( .IN1(n27487), .IN2(n28748), .IN3(n27456), .IN4(n28747), .Q(
        n27417) );
  OA22X1 U31490 ( .IN1(n27481), .IN2(n28750), .IN3(n27492), .IN4(n28749), .Q(
        n27416) );
  OA22X1 U31491 ( .IN1(n27473), .IN2(n28752), .IN3(n27478), .IN4(n28751), .Q(
        n27415) );
  OA22X1 U31492 ( .IN1(n27438), .IN2(n28746), .IN3(n27443), .IN4(n28745), .Q(
        n27414) );
  NAND4X0 U31493 ( .IN1(n27417), .IN2(n27416), .IN3(n27415), .IN4(n27414), 
        .QN(s3_addr_o[15]) );
  OA22X1 U31494 ( .IN1(n27486), .IN2(n28758), .IN3(n27443), .IN4(n28763), .Q(
        n27421) );
  OA22X1 U31495 ( .IN1(n27493), .IN2(n28760), .IN3(n27492), .IN4(n28764), .Q(
        n27420) );
  OA22X1 U31496 ( .IN1(n27480), .IN2(n28762), .IN3(n27489), .IN4(n28757), .Q(
        n27419) );
  OA22X1 U31497 ( .IN1(n27488), .IN2(n28761), .IN3(n27490), .IN4(n28759), .Q(
        n27418) );
  NAND4X0 U31498 ( .IN1(n27421), .IN2(n27420), .IN3(n27419), .IN4(n27418), 
        .QN(s3_addr_o[16]) );
  OA22X1 U31499 ( .IN1(n27487), .IN2(n28776), .IN3(n27456), .IN4(n28775), .Q(
        n27425) );
  OA22X1 U31500 ( .IN1(n27493), .IN2(n28774), .IN3(n27443), .IN4(n28769), .Q(
        n27424) );
  OA22X1 U31501 ( .IN1(n27486), .IN2(n28772), .IN3(n27488), .IN4(n28773), .Q(
        n27423) );
  OA22X1 U31502 ( .IN1(n27478), .IN2(n28771), .IN3(n27492), .IN4(n28770), .Q(
        n27422) );
  NAND4X0 U31503 ( .IN1(n27425), .IN2(n27424), .IN3(n27423), .IN4(n27422), 
        .QN(s3_addr_o[17]) );
  OA22X1 U31504 ( .IN1(n27480), .IN2(n28788), .IN3(n27478), .IN4(n28783), .Q(
        n27429) );
  OA22X1 U31505 ( .IN1(n27488), .IN2(n28782), .IN3(n27443), .IN4(n28781), .Q(
        n27428) );
  OA22X1 U31506 ( .IN1(n27438), .IN2(n28786), .IN3(n27490), .IN4(n28784), .Q(
        n27427) );
  OA22X1 U31507 ( .IN1(n27493), .IN2(n28787), .IN3(n27492), .IN4(n28785), .Q(
        n27426) );
  NAND4X0 U31508 ( .IN1(n27429), .IN2(n27428), .IN3(n27427), .IN4(n27426), 
        .QN(s3_addr_o[18]) );
  OA22X1 U31509 ( .IN1(n27488), .IN2(n28794), .IN3(n27489), .IN4(n28795), .Q(
        n27433) );
  OA22X1 U31510 ( .IN1(n27486), .IN2(n28796), .IN3(n27492), .IN4(n28793), .Q(
        n27432) );
  OA22X1 U31511 ( .IN1(n27456), .IN2(n28797), .IN3(n27443), .IN4(n28799), .Q(
        n27431) );
  OA22X1 U31512 ( .IN1(n27487), .IN2(n28800), .IN3(n27481), .IN4(n28798), .Q(
        n27430) );
  NAND4X0 U31513 ( .IN1(n27433), .IN2(n27432), .IN3(n27431), .IN4(n27430), 
        .QN(s3_addr_o[19]) );
  OA22X1 U31514 ( .IN1(n27487), .IN2(n28808), .IN3(n27443), .IN4(n28805), .Q(
        n27437) );
  OA22X1 U31515 ( .IN1(n27488), .IN2(n28810), .IN3(n27490), .IN4(n28806), .Q(
        n27436) );
  OA22X1 U31516 ( .IN1(n27493), .IN2(n28807), .IN3(n27489), .IN4(n28811), .Q(
        n27435) );
  OA22X1 U31517 ( .IN1(n27438), .IN2(n28812), .IN3(n27492), .IN4(n28809), .Q(
        n27434) );
  NAND4X0 U31518 ( .IN1(n27437), .IN2(n27436), .IN3(n27435), .IN4(n27434), 
        .QN(s3_addr_o[20]) );
  OA22X1 U31519 ( .IN1(n27480), .IN2(n28824), .IN3(n27481), .IN4(n28820), .Q(
        n27442) );
  OA22X1 U31520 ( .IN1(n27490), .IN2(n28821), .IN3(n27492), .IN4(n28818), .Q(
        n27441) );
  OA22X1 U31521 ( .IN1(n27438), .IN2(n28822), .IN3(n27443), .IN4(n28817), .Q(
        n27440) );
  OA22X1 U31522 ( .IN1(n27488), .IN2(n28819), .IN3(n27478), .IN4(n28823), .Q(
        n27439) );
  NAND4X0 U31523 ( .IN1(n27442), .IN2(n27441), .IN3(n27440), .IN4(n27439), 
        .QN(s3_addr_o[21]) );
  OA22X1 U31524 ( .IN1(n27480), .IN2(n28832), .IN3(n27492), .IN4(n28837), .Q(
        n27447) );
  OA22X1 U31525 ( .IN1(n27486), .IN2(n28833), .IN3(n27481), .IN4(n28831), .Q(
        n27446) );
  OA22X1 U31526 ( .IN1(n27456), .IN2(n28836), .IN3(n27478), .IN4(n28834), .Q(
        n27445) );
  OA22X1 U31527 ( .IN1(n27488), .IN2(n28838), .IN3(n27443), .IN4(n28829), .Q(
        n27444) );
  NAND4X0 U31528 ( .IN1(n27447), .IN2(n27446), .IN3(n27445), .IN4(n27444), 
        .QN(s3_addr_o[22]) );
  OA22X1 U31529 ( .IN1(n27490), .IN2(n28852), .IN3(n27491), .IN4(n28851), .Q(
        n27451) );
  OA22X1 U31530 ( .IN1(n27486), .IN2(n28848), .IN3(n27492), .IN4(n28846), .Q(
        n27450) );
  OA22X1 U31531 ( .IN1(n27493), .IN2(n28843), .IN3(n27478), .IN4(n28849), .Q(
        n27449) );
  OA22X1 U31532 ( .IN1(n27480), .IN2(n28845), .IN3(n27473), .IN4(n28850), .Q(
        n27448) );
  NAND4X0 U31533 ( .IN1(n27451), .IN2(n27450), .IN3(n27449), .IN4(n27448), 
        .QN(s3_addr_o[23]) );
  OA22X1 U31534 ( .IN1(n28864), .IN2(n27480), .IN3(n28859), .IN4(n27478), .Q(
        n27455) );
  OA22X1 U31535 ( .IN1(n28863), .IN2(n27486), .IN3(n28861), .IN4(n27490), .Q(
        n27454) );
  OA22X1 U31536 ( .IN1(n28860), .IN2(n27491), .IN3(n28857), .IN4(n27473), .Q(
        n27453) );
  OA22X1 U31537 ( .IN1(n28858), .IN2(n27481), .IN3(n28865), .IN4(n27479), .Q(
        n27452) );
  NAND4X0 U31538 ( .IN1(n27455), .IN2(n27454), .IN3(n27453), .IN4(n27452), 
        .QN(s3_addr_o[24]) );
  OA22X1 U31539 ( .IN1(n28871), .IN2(n27479), .IN3(n28876), .IN4(n27478), .Q(
        n27460) );
  OA22X1 U31540 ( .IN1(n28870), .IN2(n27486), .IN3(n28874), .IN4(n27488), .Q(
        n27459) );
  OA22X1 U31541 ( .IN1(n28877), .IN2(n27487), .IN3(n28872), .IN4(n27456), .Q(
        n27458) );
  OA22X1 U31542 ( .IN1(n28873), .IN2(n27493), .IN3(n28875), .IN4(n27491), .Q(
        n27457) );
  NAND4X0 U31543 ( .IN1(n27460), .IN2(n27459), .IN3(n27458), .IN4(n27457), 
        .QN(s3_addr_o[25]) );
  OA22X1 U31544 ( .IN1(n28882), .IN2(n27473), .IN3(n28886), .IN4(n27490), .Q(
        n27464) );
  OA22X1 U31545 ( .IN1(n28889), .IN2(n27491), .IN3(n28888), .IN4(n27478), .Q(
        n27463) );
  OA22X1 U31546 ( .IN1(n28885), .IN2(n27481), .IN3(n28883), .IN4(n27479), .Q(
        n27462) );
  OA22X1 U31547 ( .IN1(n28887), .IN2(n27480), .IN3(n28884), .IN4(n27486), .Q(
        n27461) );
  NAND4X0 U31548 ( .IN1(n27464), .IN2(n27463), .IN3(n27462), .IN4(n27461), 
        .QN(s3_addr_o[26]) );
  OA22X1 U31549 ( .IN1(n28899), .IN2(n27493), .IN3(n28895), .IN4(n27480), .Q(
        n27468) );
  OA22X1 U31550 ( .IN1(n28897), .IN2(n27479), .IN3(n28894), .IN4(n27486), .Q(
        n27467) );
  OA22X1 U31551 ( .IN1(n28901), .IN2(n27488), .IN3(n28900), .IN4(n27490), .Q(
        n27466) );
  OA22X1 U31552 ( .IN1(n28898), .IN2(n27491), .IN3(n28896), .IN4(n27478), .Q(
        n27465) );
  NAND4X0 U31553 ( .IN1(n27468), .IN2(n27467), .IN3(n27466), .IN4(n27465), 
        .QN(s3_addr_o[27]) );
  OA22X1 U31554 ( .IN1(n28907), .IN2(n27479), .IN3(n28912), .IN4(n27486), .Q(
        n27472) );
  OA22X1 U31555 ( .IN1(n28913), .IN2(n27491), .IN3(n28910), .IN4(n27478), .Q(
        n27471) );
  OA22X1 U31556 ( .IN1(n28911), .IN2(n27480), .IN3(n28906), .IN4(n27490), .Q(
        n27470) );
  OA22X1 U31557 ( .IN1(n28909), .IN2(n27481), .IN3(n28908), .IN4(n27473), .Q(
        n27469) );
  NAND4X0 U31558 ( .IN1(n27472), .IN2(n27471), .IN3(n27470), .IN4(n27469), 
        .QN(s3_addr_o[28]) );
  OA22X1 U31559 ( .IN1(n28920), .IN2(n27489), .IN3(n28919), .IN4(n27473), .Q(
        n27477) );
  OA22X1 U31560 ( .IN1(n28922), .IN2(n27479), .IN3(n28921), .IN4(n27491), .Q(
        n27476) );
  OA22X1 U31561 ( .IN1(n28924), .IN2(n27487), .IN3(n28925), .IN4(n27486), .Q(
        n27475) );
  OA22X1 U31562 ( .IN1(n28926), .IN2(n27493), .IN3(n28923), .IN4(n27490), .Q(
        n27474) );
  NAND4X0 U31563 ( .IN1(n27477), .IN2(n27476), .IN3(n27475), .IN4(n27474), 
        .QN(s3_addr_o[29]) );
  OA22X1 U31564 ( .IN1(n28933), .IN2(n27491), .IN3(n28940), .IN4(n27488), .Q(
        n27485) );
  OA22X1 U31565 ( .IN1(n28936), .IN2(n27478), .IN3(n28931), .IN4(n27486), .Q(
        n27484) );
  OA22X1 U31566 ( .IN1(n28937), .IN2(n27479), .IN3(n28939), .IN4(n27490), .Q(
        n27483) );
  OA22X1 U31567 ( .IN1(n28932), .IN2(n27481), .IN3(n28935), .IN4(n27480), .Q(
        n27482) );
  NAND4X0 U31568 ( .IN1(n27485), .IN2(n27484), .IN3(n27483), .IN4(n27482), 
        .QN(s3_addr_o[30]) );
  OA22X1 U31569 ( .IN1(n28952), .IN2(n27487), .IN3(n28950), .IN4(n27486), .Q(
        n27497) );
  OA22X1 U31570 ( .IN1(n28954), .IN2(n27489), .IN3(n28958), .IN4(n27488), .Q(
        n27496) );
  OA22X1 U31571 ( .IN1(n28960), .IN2(n27491), .IN3(n28946), .IN4(n27490), .Q(
        n27495) );
  OA22X1 U31572 ( .IN1(n28948), .IN2(n27493), .IN3(n28956), .IN4(n27492), .Q(
        n27494) );
  NAND4X0 U31573 ( .IN1(n27497), .IN2(n27496), .IN3(n27495), .IN4(n27494), 
        .QN(s3_addr_o[31]) );
  OA22X1 U31574 ( .IN1(n29349), .IN2(n27499), .IN3(n29235), .IN4(n27498), .Q(
        n27509) );
  OA22X1 U31575 ( .IN1(n29254), .IN2(n27501), .IN3(n29292), .IN4(n27500), .Q(
        n27508) );
  OA22X1 U31576 ( .IN1(n29273), .IN2(n27503), .IN3(n29330), .IN4(n27502), .Q(
        n27507) );
  OA22X1 U31577 ( .IN1(n29368), .IN2(n27505), .IN3(n29311), .IN4(n27504), .Q(
        n27506) );
  NAND4X0 U31578 ( .IN1(n27509), .IN2(n27508), .IN3(n27507), .IN4(n27506), 
        .QN(s2_stb_o) );
  INVX0 U31579 ( .INP(n29011), .ZN(n27781) );
  INVX0 U31580 ( .INP(n29012), .ZN(n27792) );
  OA22X1 U31581 ( .IN1(n27781), .IN2(n28126), .IN3(n27792), .IN4(n28122), .Q(
        n27513) );
  INVX0 U31582 ( .INP(n29002), .ZN(n27784) );
  OA22X1 U31583 ( .IN1(n27784), .IN2(n28124), .IN3(n27772), .IN4(n28127), .Q(
        n27512) );
  INVX0 U31584 ( .INP(n29010), .ZN(n27797) );
  INVX0 U31585 ( .INP(n27747), .ZN(n29004) );
  INVX0 U31586 ( .INP(n29004), .ZN(n27794) );
  OA22X1 U31587 ( .IN1(n27797), .IN2(n28125), .IN3(n27794), .IN4(n28121), .Q(
        n27511) );
  INVX0 U31588 ( .INP(n29009), .ZN(n27795) );
  INVX0 U31589 ( .INP(n29003), .ZN(n27742) );
  OA22X1 U31590 ( .IN1(n27795), .IN2(n28128), .IN3(n27742), .IN4(n28123), .Q(
        n27510) );
  NAND4X0 U31591 ( .IN1(n27513), .IN2(n27512), .IN3(n27511), .IN4(n27510), 
        .QN(s2_we_o) );
  INVX0 U31592 ( .INP(n29011), .ZN(n27796) );
  OA22X1 U31593 ( .IN1(n27796), .IN2(n28139), .IN3(n27792), .IN4(n28138), .Q(
        n27517) );
  INVX0 U31594 ( .INP(n27772), .ZN(n29001) );
  INVX0 U31595 ( .INP(n29001), .ZN(n27793) );
  OA22X1 U31596 ( .IN1(n27793), .IN2(n28137), .IN3(n27747), .IN4(n28135), .Q(
        n27516) );
  OA22X1 U31597 ( .IN1(n27784), .IN2(n28134), .IN3(n27742), .IN4(n28133), .Q(
        n27515) );
  INVX0 U31598 ( .INP(n29009), .ZN(n27785) );
  OA22X1 U31599 ( .IN1(n27785), .IN2(n28140), .IN3(n27797), .IN4(n28136), .Q(
        n27514) );
  NAND4X0 U31600 ( .IN1(n27517), .IN2(n27516), .IN3(n27515), .IN4(n27514), 
        .QN(s2_data_o[0]) );
  INVX0 U31601 ( .INP(n29010), .ZN(n27782) );
  OA22X1 U31602 ( .IN1(n27782), .IN2(n28152), .IN3(n27747), .IN4(n28147), .Q(
        n27521) );
  OA22X1 U31603 ( .IN1(n27781), .IN2(n28145), .IN3(n27792), .IN4(n28149), .Q(
        n27520) );
  INVX0 U31604 ( .INP(n29002), .ZN(n27790) );
  OA22X1 U31605 ( .IN1(n27790), .IN2(n28150), .IN3(n27772), .IN4(n28151), .Q(
        n27519) );
  OA22X1 U31606 ( .IN1(n27785), .IN2(n28146), .IN3(n27742), .IN4(n28148), .Q(
        n27518) );
  NAND4X0 U31607 ( .IN1(n27521), .IN2(n27520), .IN3(n27519), .IN4(n27518), 
        .QN(s2_data_o[1]) );
  OA22X1 U31608 ( .IN1(n27742), .IN2(n28163), .IN3(n27772), .IN4(n28157), .Q(
        n27525) );
  OA22X1 U31609 ( .IN1(n27795), .IN2(n28164), .IN3(n27797), .IN4(n28162), .Q(
        n27524) );
  OA22X1 U31610 ( .IN1(n27792), .IN2(n28158), .IN3(n27747), .IN4(n28161), .Q(
        n27523) );
  OA22X1 U31611 ( .IN1(n27790), .IN2(n28160), .IN3(n27781), .IN4(n28159), .Q(
        n27522) );
  NAND4X0 U31612 ( .IN1(n27525), .IN2(n27524), .IN3(n27523), .IN4(n27522), 
        .QN(s2_data_o[2]) );
  INVX0 U31613 ( .INP(n29012), .ZN(n27783) );
  OA22X1 U31614 ( .IN1(n27783), .IN2(n28171), .IN3(n27747), .IN4(n28173), .Q(
        n27529) );
  OA22X1 U31615 ( .IN1(n27790), .IN2(n28172), .IN3(n27781), .IN4(n28170), .Q(
        n27528) );
  OA22X1 U31616 ( .IN1(n27782), .IN2(n28175), .IN3(n27772), .IN4(n28169), .Q(
        n27527) );
  OA22X1 U31617 ( .IN1(n27785), .IN2(n28174), .IN3(n27742), .IN4(n28176), .Q(
        n27526) );
  NAND4X0 U31618 ( .IN1(n27529), .IN2(n27528), .IN3(n27527), .IN4(n27526), 
        .QN(s2_data_o[3]) );
  OA22X1 U31619 ( .IN1(n27782), .IN2(n28183), .IN3(n27747), .IN4(n28181), .Q(
        n27533) );
  OA22X1 U31620 ( .IN1(n27790), .IN2(n28182), .IN3(n27792), .IN4(n28185), .Q(
        n27532) );
  OA22X1 U31621 ( .IN1(n27785), .IN2(n28184), .IN3(n27781), .IN4(n28188), .Q(
        n27531) );
  OA22X1 U31622 ( .IN1(n27742), .IN2(n28186), .IN3(n27772), .IN4(n28187), .Q(
        n27530) );
  NAND4X0 U31623 ( .IN1(n27533), .IN2(n27532), .IN3(n27531), .IN4(n27530), 
        .QN(s2_data_o[4]) );
  OA22X1 U31624 ( .IN1(n27796), .IN2(n28193), .IN3(n27797), .IN4(n28197), .Q(
        n27537) );
  OA22X1 U31625 ( .IN1(n27792), .IN2(n28198), .IN3(n27747), .IN4(n28199), .Q(
        n27536) );
  OA22X1 U31626 ( .IN1(n27795), .IN2(n28200), .IN3(n27772), .IN4(n28195), .Q(
        n27535) );
  OA22X1 U31627 ( .IN1(n27790), .IN2(n28196), .IN3(n27742), .IN4(n28194), .Q(
        n27534) );
  NAND4X0 U31628 ( .IN1(n27537), .IN2(n27536), .IN3(n27535), .IN4(n27534), 
        .QN(s2_data_o[5]) );
  OA22X1 U31629 ( .IN1(n27790), .IN2(n28208), .IN3(n27785), .IN4(n28207), .Q(
        n27541) );
  INVX0 U31630 ( .INP(n29003), .ZN(n27791) );
  OA22X1 U31631 ( .IN1(n27791), .IN2(n28206), .IN3(n27772), .IN4(n28210), .Q(
        n27540) );
  OA22X1 U31632 ( .IN1(n27781), .IN2(n28212), .IN3(n27797), .IN4(n28205), .Q(
        n27539) );
  OA22X1 U31633 ( .IN1(n27783), .IN2(n28211), .IN3(n27747), .IN4(n28209), .Q(
        n27538) );
  NAND4X0 U31634 ( .IN1(n27541), .IN2(n27540), .IN3(n27539), .IN4(n27538), 
        .QN(s2_data_o[6]) );
  OA22X1 U31635 ( .IN1(n27796), .IN2(n28218), .IN3(n27794), .IN4(n28221), .Q(
        n27545) );
  OA22X1 U31636 ( .IN1(n27795), .IN2(n28219), .IN3(n27742), .IN4(n28224), .Q(
        n27544) );
  OA22X1 U31637 ( .IN1(n27782), .IN2(n28223), .IN3(n27772), .IN4(n28222), .Q(
        n27543) );
  OA22X1 U31638 ( .IN1(n27790), .IN2(n28220), .IN3(n27792), .IN4(n28217), .Q(
        n27542) );
  NAND4X0 U31639 ( .IN1(n27545), .IN2(n27544), .IN3(n27543), .IN4(n27542), 
        .QN(s2_data_o[7]) );
  OA22X1 U31640 ( .IN1(n27793), .IN2(n28233), .IN3(n27794), .IN4(n28235), .Q(
        n27549) );
  OA22X1 U31641 ( .IN1(n27785), .IN2(n28232), .IN3(n27797), .IN4(n28229), .Q(
        n27548) );
  OA22X1 U31642 ( .IN1(n27790), .IN2(n28230), .IN3(n27742), .IN4(n28231), .Q(
        n27547) );
  OA22X1 U31643 ( .IN1(n27781), .IN2(n28234), .IN3(n27792), .IN4(n28236), .Q(
        n27546) );
  NAND4X0 U31644 ( .IN1(n27549), .IN2(n27548), .IN3(n27547), .IN4(n27546), 
        .QN(s2_data_o[8]) );
  OA22X1 U31645 ( .IN1(n27785), .IN2(n28244), .IN3(n27742), .IN4(n28246), .Q(
        n27553) );
  OA22X1 U31646 ( .IN1(n27796), .IN2(n28248), .IN3(n27797), .IN4(n28245), .Q(
        n27552) );
  OA22X1 U31647 ( .IN1(n27792), .IN2(n28241), .IN3(n27794), .IN4(n28247), .Q(
        n27551) );
  OA22X1 U31648 ( .IN1(n27784), .IN2(n28242), .IN3(n27772), .IN4(n28243), .Q(
        n27550) );
  NAND4X0 U31649 ( .IN1(n27553), .IN2(n27552), .IN3(n27551), .IN4(n27550), 
        .QN(s2_data_o[9]) );
  OA22X1 U31650 ( .IN1(n27742), .IN2(n28260), .IN3(n27781), .IN4(n28256), .Q(
        n27557) );
  OA22X1 U31651 ( .IN1(n27784), .IN2(n28258), .IN3(n27793), .IN4(n28253), .Q(
        n27556) );
  OA22X1 U31652 ( .IN1(n27783), .IN2(n28254), .IN3(n27797), .IN4(n28255), .Q(
        n27555) );
  OA22X1 U31653 ( .IN1(n27795), .IN2(n28257), .IN3(n27794), .IN4(n28259), .Q(
        n27554) );
  NAND4X0 U31654 ( .IN1(n27557), .IN2(n27556), .IN3(n27555), .IN4(n27554), 
        .QN(s2_data_o[10]) );
  OA22X1 U31655 ( .IN1(n27796), .IN2(n28271), .IN3(n27794), .IN4(n28269), .Q(
        n27561) );
  OA22X1 U31656 ( .IN1(n27790), .IN2(n28266), .IN3(n27793), .IN4(n28267), .Q(
        n27560) );
  OA22X1 U31657 ( .IN1(n27742), .IN2(n28265), .IN3(n27792), .IN4(n28268), .Q(
        n27559) );
  OA22X1 U31658 ( .IN1(n27785), .IN2(n28272), .IN3(n27797), .IN4(n28270), .Q(
        n27558) );
  NAND4X0 U31659 ( .IN1(n27561), .IN2(n27560), .IN3(n27559), .IN4(n27558), 
        .QN(s2_data_o[11]) );
  OA22X1 U31660 ( .IN1(n27796), .IN2(n28282), .IN3(n27793), .IN4(n28279), .Q(
        n27565) );
  OA22X1 U31661 ( .IN1(n27790), .IN2(n28284), .IN3(n27794), .IN4(n28277), .Q(
        n27564) );
  OA22X1 U31662 ( .IN1(n27792), .IN2(n28283), .IN3(n27797), .IN4(n28281), .Q(
        n27563) );
  OA22X1 U31663 ( .IN1(n27785), .IN2(n28278), .IN3(n27742), .IN4(n28280), .Q(
        n27562) );
  NAND4X0 U31664 ( .IN1(n27565), .IN2(n27564), .IN3(n27563), .IN4(n27562), 
        .QN(s2_data_o[12]) );
  OA22X1 U31665 ( .IN1(n27795), .IN2(n28294), .IN3(n27742), .IN4(n28296), .Q(
        n27569) );
  OA22X1 U31666 ( .IN1(n27796), .IN2(n28292), .IN3(n27797), .IN4(n28293), .Q(
        n27568) );
  OA22X1 U31667 ( .IN1(n27784), .IN2(n28290), .IN3(n27794), .IN4(n28295), .Q(
        n27567) );
  OA22X1 U31668 ( .IN1(n27783), .IN2(n28289), .IN3(n27793), .IN4(n28291), .Q(
        n27566) );
  NAND4X0 U31669 ( .IN1(n27569), .IN2(n27568), .IN3(n27567), .IN4(n27566), 
        .QN(s2_data_o[13]) );
  OA22X1 U31670 ( .IN1(n27782), .IN2(n28302), .IN3(n27794), .IN4(n28303), .Q(
        n27573) );
  OA22X1 U31671 ( .IN1(n27742), .IN2(n28308), .IN3(n27781), .IN4(n28305), .Q(
        n27572) );
  OA22X1 U31672 ( .IN1(n27790), .IN2(n28306), .IN3(n27792), .IN4(n28307), .Q(
        n27571) );
  OA22X1 U31673 ( .IN1(n27795), .IN2(n28304), .IN3(n27793), .IN4(n28301), .Q(
        n27570) );
  NAND4X0 U31674 ( .IN1(n27573), .IN2(n27572), .IN3(n27571), .IN4(n27570), 
        .QN(s2_data_o[14]) );
  OA22X1 U31675 ( .IN1(n27742), .IN2(n28314), .IN3(n27782), .IN4(n28318), .Q(
        n27577) );
  OA22X1 U31676 ( .IN1(n27785), .IN2(n28315), .IN3(n27793), .IN4(n28317), .Q(
        n27576) );
  OA22X1 U31677 ( .IN1(n27784), .IN2(n28316), .IN3(n27792), .IN4(n28320), .Q(
        n27575) );
  OA22X1 U31678 ( .IN1(n27796), .IN2(n28313), .IN3(n27794), .IN4(n28319), .Q(
        n27574) );
  NAND4X0 U31679 ( .IN1(n27577), .IN2(n27576), .IN3(n27575), .IN4(n27574), 
        .QN(s2_data_o[15]) );
  OA22X1 U31680 ( .IN1(n27785), .IN2(n28332), .IN3(n27781), .IN4(n28326), .Q(
        n27581) );
  OA22X1 U31681 ( .IN1(n27793), .IN2(n28328), .IN3(n27794), .IN4(n28327), .Q(
        n27580) );
  OA22X1 U31682 ( .IN1(n27784), .IN2(n28330), .IN3(n27782), .IN4(n28325), .Q(
        n27579) );
  OA22X1 U31683 ( .IN1(n27791), .IN2(n28331), .IN3(n27792), .IN4(n28329), .Q(
        n27578) );
  NAND4X0 U31684 ( .IN1(n27581), .IN2(n27580), .IN3(n27579), .IN4(n27578), 
        .QN(s2_data_o[16]) );
  OA22X1 U31685 ( .IN1(n27791), .IN2(n28342), .IN3(n27797), .IN4(n28339), .Q(
        n27585) );
  OA22X1 U31686 ( .IN1(n27790), .IN2(n28340), .IN3(n27785), .IN4(n28344), .Q(
        n27584) );
  OA22X1 U31687 ( .IN1(n27796), .IN2(n28338), .IN3(n27792), .IN4(n28337), .Q(
        n27583) );
  OA22X1 U31688 ( .IN1(n27772), .IN2(n28343), .IN3(n27794), .IN4(n28341), .Q(
        n27582) );
  NAND4X0 U31689 ( .IN1(n27585), .IN2(n27584), .IN3(n27583), .IN4(n27582), 
        .QN(s2_data_o[17]) );
  OA22X1 U31690 ( .IN1(n27790), .IN2(n28352), .IN3(n27797), .IN4(n28349), .Q(
        n27589) );
  OA22X1 U31691 ( .IN1(n27795), .IN2(n28356), .IN3(n27792), .IN4(n28354), .Q(
        n27588) );
  OA22X1 U31692 ( .IN1(n27742), .IN2(n28350), .IN3(n27794), .IN4(n28353), .Q(
        n27587) );
  OA22X1 U31693 ( .IN1(n27796), .IN2(n28355), .IN3(n27793), .IN4(n28351), .Q(
        n27586) );
  NAND4X0 U31694 ( .IN1(n27589), .IN2(n27588), .IN3(n27587), .IN4(n27586), 
        .QN(s2_data_o[18]) );
  OA22X1 U31695 ( .IN1(n27742), .IN2(n28362), .IN3(n27793), .IN4(n28368), .Q(
        n27593) );
  OA22X1 U31696 ( .IN1(n27796), .IN2(n28363), .IN3(n27794), .IN4(n28367), .Q(
        n27592) );
  OA22X1 U31697 ( .IN1(n27784), .IN2(n28366), .IN3(n27797), .IN4(n28361), .Q(
        n27591) );
  OA22X1 U31698 ( .IN1(n27785), .IN2(n28364), .IN3(n27792), .IN4(n28365), .Q(
        n27590) );
  NAND4X0 U31699 ( .IN1(n27593), .IN2(n27592), .IN3(n27591), .IN4(n27590), 
        .QN(s2_data_o[19]) );
  OA22X1 U31700 ( .IN1(n27795), .IN2(n28377), .IN3(n27781), .IN4(n28373), .Q(
        n27597) );
  OA22X1 U31701 ( .IN1(n27782), .IN2(n28380), .IN3(n27793), .IN4(n28379), .Q(
        n27596) );
  OA22X1 U31702 ( .IN1(n27790), .IN2(n28378), .IN3(n27792), .IN4(n28376), .Q(
        n27595) );
  OA22X1 U31703 ( .IN1(n27742), .IN2(n28374), .IN3(n27794), .IN4(n28375), .Q(
        n27594) );
  NAND4X0 U31704 ( .IN1(n27597), .IN2(n27596), .IN3(n27595), .IN4(n27594), 
        .QN(s2_data_o[20]) );
  OA22X1 U31705 ( .IN1(n27796), .IN2(n28388), .IN3(n27792), .IN4(n28387), .Q(
        n27601) );
  OA22X1 U31706 ( .IN1(n27795), .IN2(n28386), .IN3(n27742), .IN4(n28390), .Q(
        n27600) );
  OA22X1 U31707 ( .IN1(n27782), .IN2(n28385), .IN3(n27793), .IN4(n28389), .Q(
        n27599) );
  OA22X1 U31708 ( .IN1(n27790), .IN2(n28392), .IN3(n27794), .IN4(n28391), .Q(
        n27598) );
  NAND4X0 U31709 ( .IN1(n27601), .IN2(n27600), .IN3(n27599), .IN4(n27598), 
        .QN(s2_data_o[21]) );
  OA22X1 U31710 ( .IN1(n27790), .IN2(n28400), .IN3(n27785), .IN4(n28402), .Q(
        n27605) );
  OA22X1 U31711 ( .IN1(n27796), .IN2(n28403), .IN3(n27794), .IN4(n28397), .Q(
        n27604) );
  OA22X1 U31712 ( .IN1(n27782), .IN2(n28399), .IN3(n27793), .IN4(n28401), .Q(
        n27603) );
  OA22X1 U31713 ( .IN1(n27742), .IN2(n28404), .IN3(n27792), .IN4(n28398), .Q(
        n27602) );
  NAND4X0 U31714 ( .IN1(n27605), .IN2(n27604), .IN3(n27603), .IN4(n27602), 
        .QN(s2_data_o[22]) );
  OA22X1 U31715 ( .IN1(n27785), .IN2(n28415), .IN3(n27747), .IN4(n28411), .Q(
        n27609) );
  OA22X1 U31716 ( .IN1(n27791), .IN2(n28414), .IN3(n27781), .IN4(n28413), .Q(
        n27608) );
  OA22X1 U31717 ( .IN1(n27792), .IN2(n28410), .IN3(n27793), .IN4(n28409), .Q(
        n27607) );
  OA22X1 U31718 ( .IN1(n27784), .IN2(n28416), .IN3(n27782), .IN4(n28412), .Q(
        n27606) );
  NAND4X0 U31719 ( .IN1(n27609), .IN2(n27608), .IN3(n27607), .IN4(n27606), 
        .QN(s2_data_o[23]) );
  OA22X1 U31720 ( .IN1(n27742), .IN2(n28422), .IN3(n27793), .IN4(n28427), .Q(
        n27613) );
  OA22X1 U31721 ( .IN1(n27784), .IN2(n28426), .IN3(n27796), .IN4(n28421), .Q(
        n27612) );
  OA22X1 U31722 ( .IN1(n27783), .IN2(n28425), .IN3(n27747), .IN4(n28423), .Q(
        n27611) );
  OA22X1 U31723 ( .IN1(n27785), .IN2(n28424), .IN3(n27797), .IN4(n28428), .Q(
        n27610) );
  NAND4X0 U31724 ( .IN1(n27613), .IN2(n27612), .IN3(n27611), .IN4(n27610), 
        .QN(s2_data_o[24]) );
  OA22X1 U31725 ( .IN1(n27791), .IN2(n28434), .IN3(n27781), .IN4(n28439), .Q(
        n27617) );
  OA22X1 U31726 ( .IN1(n27790), .IN2(n28438), .IN3(n27792), .IN4(n28433), .Q(
        n27616) );
  OA22X1 U31727 ( .IN1(n27795), .IN2(n28440), .IN3(n27793), .IN4(n28436), .Q(
        n27615) );
  OA22X1 U31728 ( .IN1(n27782), .IN2(n28437), .IN3(n27747), .IN4(n28435), .Q(
        n27614) );
  NAND4X0 U31729 ( .IN1(n27617), .IN2(n27616), .IN3(n27615), .IN4(n27614), 
        .QN(s2_data_o[25]) );
  OA22X1 U31730 ( .IN1(n27784), .IN2(n28452), .IN3(n27747), .IN4(n28445), .Q(
        n27621) );
  OA22X1 U31731 ( .IN1(n27795), .IN2(n28451), .IN3(n27782), .IN4(n28448), .Q(
        n27620) );
  OA22X1 U31732 ( .IN1(n27796), .IN2(n28446), .IN3(n27792), .IN4(n28449), .Q(
        n27619) );
  OA22X1 U31733 ( .IN1(n27742), .IN2(n28450), .IN3(n27793), .IN4(n28447), .Q(
        n27618) );
  NAND4X0 U31734 ( .IN1(n27621), .IN2(n27620), .IN3(n27619), .IN4(n27618), 
        .QN(s2_data_o[26]) );
  OA22X1 U31735 ( .IN1(n27782), .IN2(n28463), .IN3(n27793), .IN4(n28460), .Q(
        n27625) );
  OA22X1 U31736 ( .IN1(n27784), .IN2(n28462), .IN3(n27747), .IN4(n28459), .Q(
        n27624) );
  OA22X1 U31737 ( .IN1(n27791), .IN2(n28464), .IN3(n27781), .IN4(n28458), .Q(
        n27623) );
  OA22X1 U31738 ( .IN1(n27785), .IN2(n28461), .IN3(n27783), .IN4(n28457), .Q(
        n27622) );
  NAND4X0 U31739 ( .IN1(n27625), .IN2(n27624), .IN3(n27623), .IN4(n27622), 
        .QN(s2_data_o[27]) );
  OA22X1 U31740 ( .IN1(n27790), .IN2(n28474), .IN3(n27791), .IN4(n28472), .Q(
        n27629) );
  OA22X1 U31741 ( .IN1(n27796), .IN2(n28470), .IN3(n27747), .IN4(n28473), .Q(
        n27628) );
  OA22X1 U31742 ( .IN1(n27783), .IN2(n28471), .IN3(n27782), .IN4(n28475), .Q(
        n27627) );
  OA22X1 U31743 ( .IN1(n27795), .IN2(n28476), .IN3(n27772), .IN4(n28469), .Q(
        n27626) );
  NAND4X0 U31744 ( .IN1(n27629), .IN2(n27628), .IN3(n27627), .IN4(n27626), 
        .QN(s2_data_o[28]) );
  OA22X1 U31745 ( .IN1(n27783), .IN2(n28487), .IN3(n27797), .IN4(n28483), .Q(
        n27633) );
  OA22X1 U31746 ( .IN1(n27796), .IN2(n28486), .IN3(n27772), .IN4(n28485), .Q(
        n27632) );
  OA22X1 U31747 ( .IN1(n27790), .IN2(n28484), .IN3(n27747), .IN4(n28481), .Q(
        n27631) );
  OA22X1 U31748 ( .IN1(n27795), .IN2(n28482), .IN3(n27791), .IN4(n28488), .Q(
        n27630) );
  NAND4X0 U31749 ( .IN1(n27633), .IN2(n27632), .IN3(n27631), .IN4(n27630), 
        .QN(s2_data_o[29]) );
  OA22X1 U31750 ( .IN1(n27742), .IN2(n28497), .IN3(n27772), .IN4(n28500), .Q(
        n27637) );
  OA22X1 U31751 ( .IN1(n27782), .IN2(n28495), .IN3(n27747), .IN4(n28499), .Q(
        n27636) );
  OA22X1 U31752 ( .IN1(n27790), .IN2(n28494), .IN3(n27781), .IN4(n28496), .Q(
        n27635) );
  OA22X1 U31753 ( .IN1(n27785), .IN2(n28498), .IN3(n27792), .IN4(n28493), .Q(
        n27634) );
  NAND4X0 U31754 ( .IN1(n27637), .IN2(n27636), .IN3(n27635), .IN4(n27634), 
        .QN(s2_data_o[30]) );
  OA22X1 U31755 ( .IN1(n27795), .IN2(n28509), .IN3(n27772), .IN4(n28511), .Q(
        n27641) );
  OA22X1 U31756 ( .IN1(n27796), .IN2(n28505), .IN3(n27747), .IN4(n28507), .Q(
        n27640) );
  OA22X1 U31757 ( .IN1(n27784), .IN2(n28510), .IN3(n27783), .IN4(n28512), .Q(
        n27639) );
  OA22X1 U31758 ( .IN1(n27791), .IN2(n28506), .IN3(n27797), .IN4(n28508), .Q(
        n27638) );
  NAND4X0 U31759 ( .IN1(n27641), .IN2(n27640), .IN3(n27639), .IN4(n27638), 
        .QN(s2_data_o[31]) );
  OA22X1 U31760 ( .IN1(n27784), .IN2(n28518), .IN3(n27785), .IN4(n28517), .Q(
        n27645) );
  OA22X1 U31761 ( .IN1(n27782), .IN2(n28520), .IN3(n27772), .IN4(n28521), .Q(
        n27644) );
  OA22X1 U31762 ( .IN1(n27783), .IN2(n28523), .IN3(n27747), .IN4(n28519), .Q(
        n27643) );
  OA22X1 U31763 ( .IN1(n27791), .IN2(n28522), .IN3(n27796), .IN4(n28524), .Q(
        n27642) );
  NAND4X0 U31764 ( .IN1(n27645), .IN2(n27644), .IN3(n27643), .IN4(n27642), 
        .QN(s2_sel_o[0]) );
  OA22X1 U31765 ( .IN1(n27790), .IN2(n28534), .IN3(n27792), .IN4(n28535), .Q(
        n27649) );
  OA22X1 U31766 ( .IN1(n27795), .IN2(n28532), .IN3(n27781), .IN4(n28536), .Q(
        n27648) );
  OA22X1 U31767 ( .IN1(n27791), .IN2(n28530), .IN3(n27772), .IN4(n28531), .Q(
        n27647) );
  OA22X1 U31768 ( .IN1(n27782), .IN2(n28533), .IN3(n27747), .IN4(n28529), .Q(
        n27646) );
  NAND4X0 U31769 ( .IN1(n27649), .IN2(n27648), .IN3(n27647), .IN4(n27646), 
        .QN(s2_sel_o[1]) );
  OA22X1 U31770 ( .IN1(n27783), .IN2(n28547), .IN3(n27772), .IN4(n28545), .Q(
        n27653) );
  OA22X1 U31771 ( .IN1(n27791), .IN2(n28543), .IN3(n27797), .IN4(n28542), .Q(
        n27652) );
  OA22X1 U31772 ( .IN1(n27784), .IN2(n28544), .IN3(n27796), .IN4(n28548), .Q(
        n27651) );
  OA22X1 U31773 ( .IN1(n27795), .IN2(n28546), .IN3(n27747), .IN4(n28541), .Q(
        n27650) );
  NAND4X0 U31774 ( .IN1(n27653), .IN2(n27652), .IN3(n27651), .IN4(n27650), 
        .QN(s2_sel_o[2]) );
  OA22X1 U31775 ( .IN1(n27784), .IN2(n28558), .IN3(n27772), .IN4(n28559), .Q(
        n27657) );
  OA22X1 U31776 ( .IN1(n27792), .IN2(n28556), .IN3(n27747), .IN4(n28555), .Q(
        n27656) );
  OA22X1 U31777 ( .IN1(n27742), .IN2(n28553), .IN3(n27781), .IN4(n28557), .Q(
        n27655) );
  OA22X1 U31778 ( .IN1(n27795), .IN2(n28554), .IN3(n27797), .IN4(n28560), .Q(
        n27654) );
  NAND4X0 U31779 ( .IN1(n27657), .IN2(n27656), .IN3(n27655), .IN4(n27654), 
        .QN(s2_sel_o[3]) );
  OA22X1 U31780 ( .IN1(n27791), .IN2(n28571), .IN3(n27781), .IN4(n28566), .Q(
        n27661) );
  OA22X1 U31781 ( .IN1(n27782), .IN2(n28567), .IN3(n27772), .IN4(n28565), .Q(
        n27660) );
  OA22X1 U31782 ( .IN1(n27795), .IN2(n28570), .IN3(n27747), .IN4(n28569), .Q(
        n27659) );
  OA22X1 U31783 ( .IN1(n27784), .IN2(n28572), .IN3(n27783), .IN4(n28568), .Q(
        n27658) );
  NAND4X0 U31784 ( .IN1(n27661), .IN2(n27660), .IN3(n27659), .IN4(n27658), 
        .QN(s2_addr_o[0]) );
  OA22X1 U31785 ( .IN1(n27795), .IN2(n28578), .IN3(n27742), .IN4(n28582), .Q(
        n27665) );
  OA22X1 U31786 ( .IN1(n27784), .IN2(n28580), .IN3(n27781), .IN4(n28581), .Q(
        n27664) );
  OA22X1 U31787 ( .IN1(n27782), .IN2(n28584), .IN3(n27772), .IN4(n28577), .Q(
        n27663) );
  OA22X1 U31788 ( .IN1(n27783), .IN2(n28579), .IN3(n27747), .IN4(n28583), .Q(
        n27662) );
  NAND4X0 U31789 ( .IN1(n27665), .IN2(n27664), .IN3(n27663), .IN4(n27662), 
        .QN(s2_addr_o[1]) );
  OA22X1 U31790 ( .IN1(n28596), .IN2(n27794), .IN3(n28593), .IN4(n27797), .Q(
        n27669) );
  OA22X1 U31791 ( .IN1(n28594), .IN2(n27791), .IN3(n28595), .IN4(n27772), .Q(
        n27668) );
  OA22X1 U31792 ( .IN1(n28592), .IN2(n27796), .IN3(n28589), .IN4(n27785), .Q(
        n27667) );
  OA22X1 U31793 ( .IN1(n28591), .IN2(n27784), .IN3(n28590), .IN4(n27792), .Q(
        n27666) );
  NAND4X0 U31794 ( .IN1(n27669), .IN2(n27668), .IN3(n27667), .IN4(n27666), 
        .QN(s2_addr_o[2]) );
  OA22X1 U31795 ( .IN1(n28601), .IN2(n27790), .IN3(n28607), .IN4(n27781), .Q(
        n27673) );
  OA22X1 U31796 ( .IN1(n28602), .IN2(n27782), .IN3(n28605), .IN4(n27785), .Q(
        n27672) );
  OA22X1 U31797 ( .IN1(n28606), .IN2(n27792), .IN3(n28603), .IN4(n27772), .Q(
        n27671) );
  OA22X1 U31798 ( .IN1(n28604), .IN2(n27791), .IN3(n28608), .IN4(n27794), .Q(
        n27670) );
  NAND4X0 U31799 ( .IN1(n27673), .IN2(n27672), .IN3(n27671), .IN4(n27670), 
        .QN(s2_addr_o[3]) );
  OA22X1 U31800 ( .IN1(n28618), .IN2(n27781), .IN3(n28615), .IN4(n27792), .Q(
        n27677) );
  OA22X1 U31801 ( .IN1(n28619), .IN2(n27794), .IN3(n28614), .IN4(n27782), .Q(
        n27676) );
  OA22X1 U31802 ( .IN1(n28617), .IN2(n27784), .IN3(n28613), .IN4(n27791), .Q(
        n27675) );
  OA22X1 U31803 ( .IN1(n28616), .IN2(n27785), .IN3(n28620), .IN4(n27772), .Q(
        n27674) );
  NAND4X0 U31804 ( .IN1(n27677), .IN2(n27676), .IN3(n27675), .IN4(n27674), 
        .QN(s2_addr_o[4]) );
  OA22X1 U31805 ( .IN1(n28628), .IN2(n27793), .IN3(n28630), .IN4(n27785), .Q(
        n27681) );
  OA22X1 U31806 ( .IN1(n28632), .IN2(n27791), .IN3(n28626), .IN4(n27781), .Q(
        n27680) );
  OA22X1 U31807 ( .IN1(n28627), .IN2(n27797), .IN3(n28629), .IN4(n27790), .Q(
        n27679) );
  OA22X1 U31808 ( .IN1(n28631), .IN2(n27783), .IN3(n28625), .IN4(n27794), .Q(
        n27678) );
  NAND4X0 U31809 ( .IN1(n27681), .IN2(n27680), .IN3(n27679), .IN4(n27678), 
        .QN(s2_addr_o[5]) );
  OA22X1 U31810 ( .IN1(n27742), .IN2(n28644), .IN3(n27772), .IN4(n28641), .Q(
        n27685) );
  OA22X1 U31811 ( .IN1(n27795), .IN2(n28640), .IN3(n27782), .IN4(n28637), .Q(
        n27684) );
  OA22X1 U31812 ( .IN1(n27784), .IN2(n28642), .IN3(n27781), .IN4(n28643), .Q(
        n27683) );
  OA22X1 U31813 ( .IN1(n27783), .IN2(n28638), .IN3(n27747), .IN4(n28639), .Q(
        n27682) );
  NAND4X0 U31814 ( .IN1(n27685), .IN2(n27684), .IN3(n27683), .IN4(n27682), 
        .QN(s2_addr_o[6]) );
  OA22X1 U31815 ( .IN1(n27783), .IN2(n28650), .IN3(n27782), .IN4(n28649), .Q(
        n27689) );
  OA22X1 U31816 ( .IN1(n27796), .IN2(n28653), .IN3(n27772), .IN4(n28651), .Q(
        n27688) );
  OA22X1 U31817 ( .IN1(n27795), .IN2(n28652), .IN3(n27747), .IN4(n28655), .Q(
        n27687) );
  OA22X1 U31818 ( .IN1(n27784), .IN2(n28654), .IN3(n27742), .IN4(n28656), .Q(
        n27686) );
  NAND4X0 U31819 ( .IN1(n27689), .IN2(n27688), .IN3(n27687), .IN4(n27686), 
        .QN(s2_addr_o[7]) );
  OA22X1 U31820 ( .IN1(n27793), .IN2(n28661), .IN3(n27747), .IN4(n28667), .Q(
        n27693) );
  OA22X1 U31821 ( .IN1(n27796), .IN2(n28665), .IN3(n27782), .IN4(n28662), .Q(
        n27692) );
  OA22X1 U31822 ( .IN1(n27784), .IN2(n28664), .IN3(n27783), .IN4(n28668), .Q(
        n27691) );
  OA22X1 U31823 ( .IN1(n27795), .IN2(n28663), .IN3(n27742), .IN4(n28666), .Q(
        n27690) );
  NAND4X0 U31824 ( .IN1(n27693), .IN2(n27692), .IN3(n27691), .IN4(n27690), 
        .QN(s2_addr_o[8]) );
  OA22X1 U31825 ( .IN1(n27781), .IN2(n28676), .IN3(n27747), .IN4(n28677), .Q(
        n27697) );
  OA22X1 U31826 ( .IN1(n27784), .IN2(n28680), .IN3(n27791), .IN4(n28674), .Q(
        n27696) );
  OA22X1 U31827 ( .IN1(n27782), .IN2(n28678), .IN3(n27772), .IN4(n28675), .Q(
        n27695) );
  OA22X1 U31828 ( .IN1(n27795), .IN2(n28679), .IN3(n27792), .IN4(n28673), .Q(
        n27694) );
  NAND4X0 U31829 ( .IN1(n27697), .IN2(n27696), .IN3(n27695), .IN4(n27694), 
        .QN(s2_addr_o[9]) );
  OA22X1 U31830 ( .IN1(n27784), .IN2(n28692), .IN3(n27785), .IN4(n28686), .Q(
        n27701) );
  OA22X1 U31831 ( .IN1(n27796), .IN2(n28687), .IN3(n27797), .IN4(n28691), .Q(
        n27700) );
  OA22X1 U31832 ( .IN1(n27793), .IN2(n28690), .IN3(n27747), .IN4(n28689), .Q(
        n27699) );
  OA22X1 U31833 ( .IN1(n27791), .IN2(n28688), .IN3(n27783), .IN4(n28685), .Q(
        n27698) );
  NAND4X0 U31834 ( .IN1(n27701), .IN2(n27700), .IN3(n27699), .IN4(n27698), 
        .QN(s2_addr_o[10]) );
  OA22X1 U31835 ( .IN1(n27781), .IN2(n28704), .IN3(n27782), .IN4(n28703), .Q(
        n27705) );
  OA22X1 U31836 ( .IN1(n27784), .IN2(n28702), .IN3(n27785), .IN4(n28698), .Q(
        n27704) );
  OA22X1 U31837 ( .IN1(n27742), .IN2(n28697), .IN3(n27792), .IN4(n28701), .Q(
        n27703) );
  OA22X1 U31838 ( .IN1(n27772), .IN2(n28700), .IN3(n27747), .IN4(n28699), .Q(
        n27702) );
  NAND4X0 U31839 ( .IN1(n27705), .IN2(n27704), .IN3(n27703), .IN4(n27702), 
        .QN(s2_addr_o[11]) );
  OA22X1 U31840 ( .IN1(n27796), .IN2(n28716), .IN3(n27747), .IN4(n28713), .Q(
        n27709) );
  OA22X1 U31841 ( .IN1(n27784), .IN2(n28714), .IN3(n27783), .IN4(n28709), .Q(
        n27708) );
  OA22X1 U31842 ( .IN1(n27791), .IN2(n28712), .IN3(n27772), .IN4(n28711), .Q(
        n27707) );
  OA22X1 U31843 ( .IN1(n27795), .IN2(n28710), .IN3(n27797), .IN4(n28715), .Q(
        n27706) );
  NAND4X0 U31844 ( .IN1(n27709), .IN2(n27708), .IN3(n27707), .IN4(n27706), 
        .QN(s2_addr_o[12]) );
  OA22X1 U31845 ( .IN1(n27781), .IN2(n28724), .IN3(n27772), .IN4(n28725), .Q(
        n27713) );
  OA22X1 U31846 ( .IN1(n27742), .IN2(n28726), .IN3(n27797), .IN4(n28721), .Q(
        n27712) );
  OA22X1 U31847 ( .IN1(n27795), .IN2(n28728), .IN3(n27747), .IN4(n28727), .Q(
        n27711) );
  OA22X1 U31848 ( .IN1(n27784), .IN2(n28722), .IN3(n27783), .IN4(n28723), .Q(
        n27710) );
  NAND4X0 U31849 ( .IN1(n27713), .IN2(n27712), .IN3(n27711), .IN4(n27710), 
        .QN(s2_addr_o[13]) );
  OA22X1 U31850 ( .IN1(n27797), .IN2(n28737), .IN3(n27747), .IN4(n28739), .Q(
        n27717) );
  OA22X1 U31851 ( .IN1(n27790), .IN2(n28734), .IN3(n27796), .IN4(n28735), .Q(
        n27716) );
  OA22X1 U31852 ( .IN1(n27795), .IN2(n28738), .IN3(n27772), .IN4(n28733), .Q(
        n27715) );
  OA22X1 U31853 ( .IN1(n27791), .IN2(n28736), .IN3(n27792), .IN4(n28740), .Q(
        n27714) );
  NAND4X0 U31854 ( .IN1(n27717), .IN2(n27716), .IN3(n27715), .IN4(n27714), 
        .QN(s2_addr_o[14]) );
  OA22X1 U31855 ( .IN1(n27796), .IN2(n28752), .IN3(n27747), .IN4(n28745), .Q(
        n27721) );
  OA22X1 U31856 ( .IN1(n27790), .IN2(n28746), .IN3(n27785), .IN4(n28748), .Q(
        n27720) );
  OA22X1 U31857 ( .IN1(n27782), .IN2(n28751), .IN3(n27772), .IN4(n28749), .Q(
        n27719) );
  OA22X1 U31858 ( .IN1(n27742), .IN2(n28750), .IN3(n27783), .IN4(n28747), .Q(
        n27718) );
  NAND4X0 U31859 ( .IN1(n27721), .IN2(n27720), .IN3(n27719), .IN4(n27718), 
        .QN(s2_addr_o[15]) );
  OA22X1 U31860 ( .IN1(n27796), .IN2(n28761), .IN3(n27797), .IN4(n28757), .Q(
        n27725) );
  OA22X1 U31861 ( .IN1(n27784), .IN2(n28758), .IN3(n27747), .IN4(n28763), .Q(
        n27724) );
  OA22X1 U31862 ( .IN1(n27791), .IN2(n28760), .IN3(n27772), .IN4(n28764), .Q(
        n27723) );
  OA22X1 U31863 ( .IN1(n27795), .IN2(n28762), .IN3(n27792), .IN4(n28759), .Q(
        n27722) );
  NAND4X0 U31864 ( .IN1(n27725), .IN2(n27724), .IN3(n27723), .IN4(n27722), 
        .QN(s2_addr_o[16]) );
  OA22X1 U31865 ( .IN1(n27785), .IN2(n28776), .IN3(n27781), .IN4(n28773), .Q(
        n27729) );
  OA22X1 U31866 ( .IN1(n27742), .IN2(n28774), .IN3(n27783), .IN4(n28775), .Q(
        n27728) );
  OA22X1 U31867 ( .IN1(n27782), .IN2(n28771), .IN3(n27747), .IN4(n28769), .Q(
        n27727) );
  OA22X1 U31868 ( .IN1(n27784), .IN2(n28772), .IN3(n27772), .IN4(n28770), .Q(
        n27726) );
  NAND4X0 U31869 ( .IN1(n27729), .IN2(n27728), .IN3(n27727), .IN4(n27726), 
        .QN(s2_addr_o[17]) );
  OA22X1 U31870 ( .IN1(n27781), .IN2(n28782), .IN3(n27797), .IN4(n28783), .Q(
        n27733) );
  OA22X1 U31871 ( .IN1(n27783), .IN2(n28784), .IN3(n27747), .IN4(n28781), .Q(
        n27732) );
  OA22X1 U31872 ( .IN1(n27790), .IN2(n28786), .IN3(n27742), .IN4(n28787), .Q(
        n27731) );
  OA22X1 U31873 ( .IN1(n27795), .IN2(n28788), .IN3(n27772), .IN4(n28785), .Q(
        n27730) );
  NAND4X0 U31874 ( .IN1(n27733), .IN2(n27732), .IN3(n27731), .IN4(n27730), 
        .QN(s2_addr_o[18]) );
  OA22X1 U31875 ( .IN1(n27784), .IN2(n28796), .IN3(n27797), .IN4(n28795), .Q(
        n27737) );
  OA22X1 U31876 ( .IN1(n27796), .IN2(n28794), .IN3(n27792), .IN4(n28797), .Q(
        n27736) );
  OA22X1 U31877 ( .IN1(n27791), .IN2(n28798), .IN3(n27772), .IN4(n28793), .Q(
        n27735) );
  OA22X1 U31878 ( .IN1(n27785), .IN2(n28800), .IN3(n27747), .IN4(n28799), .Q(
        n27734) );
  NAND4X0 U31879 ( .IN1(n27737), .IN2(n27736), .IN3(n27735), .IN4(n27734), 
        .QN(s2_addr_o[19]) );
  OA22X1 U31880 ( .IN1(n27795), .IN2(n28808), .IN3(n27797), .IN4(n28811), .Q(
        n27741) );
  OA22X1 U31881 ( .IN1(n27790), .IN2(n28812), .IN3(n27747), .IN4(n28805), .Q(
        n27740) );
  OA22X1 U31882 ( .IN1(n27742), .IN2(n28807), .IN3(n27781), .IN4(n28810), .Q(
        n27739) );
  OA22X1 U31883 ( .IN1(n27783), .IN2(n28806), .IN3(n27772), .IN4(n28809), .Q(
        n27738) );
  NAND4X0 U31884 ( .IN1(n27741), .IN2(n27740), .IN3(n27739), .IN4(n27738), 
        .QN(s2_addr_o[20]) );
  OA22X1 U31885 ( .IN1(n27784), .IN2(n28822), .IN3(n27742), .IN4(n28820), .Q(
        n27746) );
  OA22X1 U31886 ( .IN1(n27797), .IN2(n28823), .IN3(n27747), .IN4(n28817), .Q(
        n27745) );
  OA22X1 U31887 ( .IN1(n27781), .IN2(n28819), .IN3(n27772), .IN4(n28818), .Q(
        n27744) );
  OA22X1 U31888 ( .IN1(n27785), .IN2(n28824), .IN3(n27783), .IN4(n28821), .Q(
        n27743) );
  NAND4X0 U31889 ( .IN1(n27746), .IN2(n27745), .IN3(n27744), .IN4(n27743), 
        .QN(s2_addr_o[21]) );
  OA22X1 U31890 ( .IN1(n27783), .IN2(n28836), .IN3(n27747), .IN4(n28829), .Q(
        n27751) );
  OA22X1 U31891 ( .IN1(n27791), .IN2(n28831), .IN3(n27781), .IN4(n28838), .Q(
        n27750) );
  OA22X1 U31892 ( .IN1(n27784), .IN2(n28833), .IN3(n27797), .IN4(n28834), .Q(
        n27749) );
  OA22X1 U31893 ( .IN1(n27795), .IN2(n28832), .IN3(n27772), .IN4(n28837), .Q(
        n27748) );
  NAND4X0 U31894 ( .IN1(n27751), .IN2(n27750), .IN3(n27749), .IN4(n27748), 
        .QN(s2_addr_o[22]) );
  OA22X1 U31895 ( .IN1(n27796), .IN2(n28850), .IN3(n27783), .IN4(n28852), .Q(
        n27755) );
  OA22X1 U31896 ( .IN1(n27785), .IN2(n28845), .IN3(n27797), .IN4(n28849), .Q(
        n27754) );
  OA22X1 U31897 ( .IN1(n27791), .IN2(n28843), .IN3(n27794), .IN4(n28851), .Q(
        n27753) );
  OA22X1 U31898 ( .IN1(n27790), .IN2(n28848), .IN3(n27772), .IN4(n28846), .Q(
        n27752) );
  NAND4X0 U31899 ( .IN1(n27755), .IN2(n27754), .IN3(n27753), .IN4(n27752), 
        .QN(s2_addr_o[23]) );
  OA22X1 U31900 ( .IN1(n28864), .IN2(n27795), .IN3(n28863), .IN4(n27790), .Q(
        n27759) );
  OA22X1 U31901 ( .IN1(n28865), .IN2(n27793), .IN3(n28861), .IN4(n27783), .Q(
        n27758) );
  OA22X1 U31902 ( .IN1(n28858), .IN2(n27791), .IN3(n28860), .IN4(n27794), .Q(
        n27757) );
  OA22X1 U31903 ( .IN1(n28859), .IN2(n27782), .IN3(n28857), .IN4(n27781), .Q(
        n27756) );
  NAND4X0 U31904 ( .IN1(n27759), .IN2(n27758), .IN3(n27757), .IN4(n27756), 
        .QN(s2_addr_o[24]) );
  OA22X1 U31905 ( .IN1(n28875), .IN2(n27794), .IN3(n28874), .IN4(n27796), .Q(
        n27763) );
  OA22X1 U31906 ( .IN1(n28873), .IN2(n27791), .IN3(n28877), .IN4(n27785), .Q(
        n27762) );
  OA22X1 U31907 ( .IN1(n28871), .IN2(n27793), .IN3(n28876), .IN4(n27797), .Q(
        n27761) );
  OA22X1 U31908 ( .IN1(n28870), .IN2(n27790), .IN3(n28872), .IN4(n27783), .Q(
        n27760) );
  NAND4X0 U31909 ( .IN1(n27763), .IN2(n27762), .IN3(n27761), .IN4(n27760), 
        .QN(s2_addr_o[25]) );
  OA22X1 U31910 ( .IN1(n28883), .IN2(n27793), .IN3(n28886), .IN4(n27783), .Q(
        n27767) );
  OA22X1 U31911 ( .IN1(n28888), .IN2(n27797), .IN3(n28884), .IN4(n27790), .Q(
        n27766) );
  OA22X1 U31912 ( .IN1(n28885), .IN2(n27791), .IN3(n28887), .IN4(n27785), .Q(
        n27765) );
  OA22X1 U31913 ( .IN1(n28889), .IN2(n27794), .IN3(n28882), .IN4(n27796), .Q(
        n27764) );
  NAND4X0 U31914 ( .IN1(n27767), .IN2(n27766), .IN3(n27765), .IN4(n27764), 
        .QN(s2_addr_o[26]) );
  OA22X1 U31915 ( .IN1(n28897), .IN2(n27793), .IN3(n28896), .IN4(n27782), .Q(
        n27771) );
  OA22X1 U31916 ( .IN1(n28898), .IN2(n27794), .IN3(n28900), .IN4(n27783), .Q(
        n27770) );
  OA22X1 U31917 ( .IN1(n28895), .IN2(n27785), .IN3(n28894), .IN4(n27790), .Q(
        n27769) );
  OA22X1 U31918 ( .IN1(n28899), .IN2(n27791), .IN3(n28901), .IN4(n27781), .Q(
        n27768) );
  NAND4X0 U31919 ( .IN1(n27771), .IN2(n27770), .IN3(n27769), .IN4(n27768), 
        .QN(s2_addr_o[27]) );
  OA22X1 U31920 ( .IN1(n28913), .IN2(n27794), .IN3(n28908), .IN4(n27781), .Q(
        n27776) );
  OA22X1 U31921 ( .IN1(n28911), .IN2(n27795), .IN3(n28912), .IN4(n27790), .Q(
        n27775) );
  OA22X1 U31922 ( .IN1(n28909), .IN2(n27791), .IN3(n28907), .IN4(n27772), .Q(
        n27774) );
  OA22X1 U31923 ( .IN1(n28910), .IN2(n27782), .IN3(n28906), .IN4(n27783), .Q(
        n27773) );
  NAND4X0 U31924 ( .IN1(n27776), .IN2(n27775), .IN3(n27774), .IN4(n27773), 
        .QN(s2_addr_o[28]) );
  OA22X1 U31925 ( .IN1(n28922), .IN2(n27793), .IN3(n28925), .IN4(n27790), .Q(
        n27780) );
  OA22X1 U31926 ( .IN1(n28920), .IN2(n27797), .IN3(n28923), .IN4(n27783), .Q(
        n27779) );
  OA22X1 U31927 ( .IN1(n28926), .IN2(n27791), .IN3(n28919), .IN4(n27781), .Q(
        n27778) );
  OA22X1 U31928 ( .IN1(n28924), .IN2(n27785), .IN3(n28921), .IN4(n27794), .Q(
        n27777) );
  NAND4X0 U31929 ( .IN1(n27780), .IN2(n27779), .IN3(n27778), .IN4(n27777), 
        .QN(s2_addr_o[29]) );
  OA22X1 U31930 ( .IN1(n28936), .IN2(n27782), .IN3(n28940), .IN4(n27781), .Q(
        n27789) );
  OA22X1 U31931 ( .IN1(n28931), .IN2(n27784), .IN3(n28939), .IN4(n27783), .Q(
        n27788) );
  OA22X1 U31932 ( .IN1(n28932), .IN2(n27791), .IN3(n28935), .IN4(n27785), .Q(
        n27787) );
  OA22X1 U31933 ( .IN1(n28937), .IN2(n27793), .IN3(n28933), .IN4(n27794), .Q(
        n27786) );
  NAND4X0 U31934 ( .IN1(n27789), .IN2(n27788), .IN3(n27787), .IN4(n27786), 
        .QN(s2_addr_o[30]) );
  OA22X1 U31935 ( .IN1(n28948), .IN2(n27791), .IN3(n28950), .IN4(n27790), .Q(
        n27801) );
  OA22X1 U31936 ( .IN1(n28956), .IN2(n27793), .IN3(n28946), .IN4(n27792), .Q(
        n27800) );
  OA22X1 U31937 ( .IN1(n28952), .IN2(n27795), .IN3(n28960), .IN4(n27794), .Q(
        n27799) );
  OA22X1 U31938 ( .IN1(n28954), .IN2(n27797), .IN3(n28958), .IN4(n27796), .Q(
        n27798) );
  NAND4X0 U31939 ( .IN1(n27801), .IN2(n27800), .IN3(n27799), .IN4(n27798), 
        .QN(s2_addr_o[31]) );
  OA22X1 U31940 ( .IN1(n29330), .IN2(n27803), .IN3(n29292), .IN4(n27802), .Q(
        n27815) );
  INVX0 U31941 ( .INP(n27804), .ZN(n27806) );
  OA22X1 U31942 ( .IN1(n29254), .IN2(n27806), .IN3(n29311), .IN4(n27805), .Q(
        n27814) );
  INVX0 U31943 ( .INP(n27807), .ZN(n27808) );
  OA22X1 U31944 ( .IN1(n29368), .IN2(n27809), .IN3(n29235), .IN4(n27808), .Q(
        n27813) );
  OA22X1 U31945 ( .IN1(n29273), .IN2(n27811), .IN3(n29349), .IN4(n27810), .Q(
        n27812) );
  NAND4X0 U31946 ( .IN1(n27815), .IN2(n27814), .IN3(n27813), .IN4(n27812), 
        .QN(s1_stb_o) );
  INVX0 U31947 ( .INP(n28985), .ZN(n28097) );
  INVX0 U31948 ( .INP(n28992), .ZN(n28088) );
  OA22X1 U31949 ( .IN1(n28097), .IN2(n28123), .IN3(n28088), .IN4(n28122), .Q(
        n27819) );
  INVX0 U31950 ( .INP(n28090), .ZN(n28986) );
  INVX0 U31951 ( .INP(n28986), .ZN(n28100) );
  OA22X1 U31952 ( .IN1(n28100), .IN2(n28126), .IN3(n28078), .IN4(n28127), .Q(
        n27818) );
  INVX0 U31953 ( .INP(n28993), .ZN(n28091) );
  INVX0 U31954 ( .INP(n28991), .ZN(n28102) );
  OA22X1 U31955 ( .IN1(n28091), .IN2(n28128), .IN3(n28102), .IN4(n28125), .Q(
        n27817) );
  INVX0 U31956 ( .INP(n28057), .ZN(n28994) );
  INVX0 U31957 ( .INP(n28994), .ZN(n28099) );
  OA22X1 U31958 ( .IN1(n28098), .IN2(n28124), .IN3(n28099), .IN4(n28121), .Q(
        n27816) );
  NAND4X0 U31959 ( .IN1(n27819), .IN2(n27818), .IN3(n27817), .IN4(n27816), 
        .QN(s1_we_o) );
  INVX0 U31960 ( .INP(n28991), .ZN(n28079) );
  OA22X1 U31961 ( .IN1(n28079), .IN2(n28136), .IN3(n28078), .IN4(n28137), .Q(
        n27823) );
  OA22X1 U31962 ( .IN1(n28091), .IN2(n28140), .IN3(n28057), .IN4(n28135), .Q(
        n27822) );
  OA22X1 U31963 ( .IN1(n28098), .IN2(n28134), .IN3(n28097), .IN4(n28133), .Q(
        n27821) );
  INVX0 U31964 ( .INP(n28992), .ZN(n28096) );
  OA22X1 U31965 ( .IN1(n28100), .IN2(n28139), .IN3(n28096), .IN4(n28138), .Q(
        n27820) );
  NAND4X0 U31966 ( .IN1(n27823), .IN2(n27822), .IN3(n27821), .IN4(n27820), 
        .QN(s1_data_o[0]) );
  OA22X1 U31967 ( .IN1(n28103), .IN2(n28146), .IN3(n28078), .IN4(n28151), .Q(
        n27827) );
  OA22X1 U31968 ( .IN1(n28088), .IN2(n28149), .IN3(n28079), .IN4(n28152), .Q(
        n27826) );
  INVX0 U31969 ( .INP(n28984), .ZN(n28056) );
  OA22X1 U31970 ( .IN1(n28056), .IN2(n28150), .IN3(n28090), .IN4(n28145), .Q(
        n27825) );
  OA22X1 U31971 ( .IN1(n28089), .IN2(n28148), .IN3(n28057), .IN4(n28147), .Q(
        n27824) );
  NAND4X0 U31972 ( .IN1(n27827), .IN2(n27826), .IN3(n27825), .IN4(n27824), 
        .QN(s1_data_o[1]) );
  OA22X1 U31973 ( .IN1(n28091), .IN2(n28164), .IN3(n28097), .IN4(n28163), .Q(
        n27831) );
  OA22X1 U31974 ( .IN1(n28102), .IN2(n28162), .IN3(n28057), .IN4(n28161), .Q(
        n27830) );
  OA22X1 U31975 ( .IN1(n28096), .IN2(n28158), .IN3(n28078), .IN4(n28157), .Q(
        n27829) );
  OA22X1 U31976 ( .IN1(n28098), .IN2(n28160), .IN3(n28090), .IN4(n28159), .Q(
        n27828) );
  NAND4X0 U31977 ( .IN1(n27831), .IN2(n27830), .IN3(n27829), .IN4(n27828), 
        .QN(s1_data_o[2]) );
  OA22X1 U31978 ( .IN1(n28103), .IN2(n28174), .IN3(n28057), .IN4(n28173), .Q(
        n27835) );
  OA22X1 U31979 ( .IN1(n28056), .IN2(n28172), .IN3(n28097), .IN4(n28176), .Q(
        n27834) );
  OA22X1 U31980 ( .IN1(n28088), .IN2(n28171), .IN3(n28079), .IN4(n28175), .Q(
        n27833) );
  OA22X1 U31981 ( .IN1(n28100), .IN2(n28170), .IN3(n28078), .IN4(n28169), .Q(
        n27832) );
  NAND4X0 U31982 ( .IN1(n27835), .IN2(n27834), .IN3(n27833), .IN4(n27832), 
        .QN(s1_data_o[3]) );
  OA22X1 U31983 ( .IN1(n28091), .IN2(n28184), .IN3(n28057), .IN4(n28181), .Q(
        n27839) );
  OA22X1 U31984 ( .IN1(n28098), .IN2(n28182), .IN3(n28078), .IN4(n28187), .Q(
        n27838) );
  OA22X1 U31985 ( .IN1(n28097), .IN2(n28186), .IN3(n28079), .IN4(n28183), .Q(
        n27837) );
  OA22X1 U31986 ( .IN1(n28100), .IN2(n28188), .IN3(n28096), .IN4(n28185), .Q(
        n27836) );
  NAND4X0 U31987 ( .IN1(n27839), .IN2(n27838), .IN3(n27837), .IN4(n27836), 
        .QN(s1_data_o[4]) );
  OA22X1 U31988 ( .IN1(n28103), .IN2(n28200), .IN3(n28079), .IN4(n28197), .Q(
        n27843) );
  OA22X1 U31989 ( .IN1(n28100), .IN2(n28193), .IN3(n28078), .IN4(n28195), .Q(
        n27842) );
  OA22X1 U31990 ( .IN1(n28089), .IN2(n28194), .IN3(n28057), .IN4(n28199), .Q(
        n27841) );
  OA22X1 U31991 ( .IN1(n28056), .IN2(n28196), .IN3(n28096), .IN4(n28198), .Q(
        n27840) );
  NAND4X0 U31992 ( .IN1(n27843), .IN2(n27842), .IN3(n27841), .IN4(n27840), 
        .QN(s1_data_o[5]) );
  OA22X1 U31993 ( .IN1(n28098), .IN2(n28208), .IN3(n28078), .IN4(n28210), .Q(
        n27847) );
  OA22X1 U31994 ( .IN1(n28100), .IN2(n28212), .IN3(n28096), .IN4(n28211), .Q(
        n27846) );
  OA22X1 U31995 ( .IN1(n28089), .IN2(n28206), .IN3(n28079), .IN4(n28205), .Q(
        n27845) );
  OA22X1 U31996 ( .IN1(n28103), .IN2(n28207), .IN3(n28057), .IN4(n28209), .Q(
        n27844) );
  NAND4X0 U31997 ( .IN1(n27847), .IN2(n27846), .IN3(n27845), .IN4(n27844), 
        .QN(s1_data_o[6]) );
  OA22X1 U31998 ( .IN1(n28079), .IN2(n28223), .IN3(n28057), .IN4(n28221), .Q(
        n27851) );
  OA22X1 U31999 ( .IN1(n28091), .IN2(n28219), .IN3(n28090), .IN4(n28218), .Q(
        n27850) );
  OA22X1 U32000 ( .IN1(n28056), .IN2(n28220), .IN3(n28078), .IN4(n28222), .Q(
        n27849) );
  OA22X1 U32001 ( .IN1(n28089), .IN2(n28224), .IN3(n28096), .IN4(n28217), .Q(
        n27848) );
  NAND4X0 U32002 ( .IN1(n27851), .IN2(n27850), .IN3(n27849), .IN4(n27848), 
        .QN(s1_data_o[7]) );
  OA22X1 U32003 ( .IN1(n28100), .IN2(n28234), .IN3(n28079), .IN4(n28229), .Q(
        n27855) );
  INVX0 U32004 ( .INP(n28078), .ZN(n28983) );
  INVX0 U32005 ( .INP(n28983), .ZN(n28101) );
  OA22X1 U32006 ( .IN1(n28098), .IN2(n28230), .IN3(n28101), .IN4(n28233), .Q(
        n27854) );
  OA22X1 U32007 ( .IN1(n28096), .IN2(n28236), .IN3(n28099), .IN4(n28235), .Q(
        n27853) );
  OA22X1 U32008 ( .IN1(n28103), .IN2(n28232), .IN3(n28097), .IN4(n28231), .Q(
        n27852) );
  NAND4X0 U32009 ( .IN1(n27855), .IN2(n27854), .IN3(n27853), .IN4(n27852), 
        .QN(s1_data_o[8]) );
  OA22X1 U32010 ( .IN1(n28097), .IN2(n28246), .IN3(n28099), .IN4(n28247), .Q(
        n27859) );
  OA22X1 U32011 ( .IN1(n28056), .IN2(n28242), .IN3(n28079), .IN4(n28245), .Q(
        n27858) );
  OA22X1 U32012 ( .IN1(n28091), .IN2(n28244), .IN3(n28096), .IN4(n28241), .Q(
        n27857) );
  OA22X1 U32013 ( .IN1(n28090), .IN2(n28248), .IN3(n28101), .IN4(n28243), .Q(
        n27856) );
  NAND4X0 U32014 ( .IN1(n27859), .IN2(n27858), .IN3(n27857), .IN4(n27856), 
        .QN(s1_data_o[9]) );
  OA22X1 U32015 ( .IN1(n28098), .IN2(n28258), .IN3(n28096), .IN4(n28254), .Q(
        n27863) );
  OA22X1 U32016 ( .IN1(n28102), .IN2(n28255), .IN3(n28101), .IN4(n28253), .Q(
        n27862) );
  OA22X1 U32017 ( .IN1(n28103), .IN2(n28257), .IN3(n28099), .IN4(n28259), .Q(
        n27861) );
  OA22X1 U32018 ( .IN1(n28089), .IN2(n28260), .IN3(n28090), .IN4(n28256), .Q(
        n27860) );
  NAND4X0 U32019 ( .IN1(n27863), .IN2(n27862), .IN3(n27861), .IN4(n27860), 
        .QN(s1_data_o[10]) );
  OA22X1 U32020 ( .IN1(n28088), .IN2(n28268), .IN3(n28101), .IN4(n28267), .Q(
        n27867) );
  OA22X1 U32021 ( .IN1(n28079), .IN2(n28270), .IN3(n28099), .IN4(n28269), .Q(
        n27866) );
  OA22X1 U32022 ( .IN1(n28056), .IN2(n28266), .IN3(n28091), .IN4(n28272), .Q(
        n27865) );
  OA22X1 U32023 ( .IN1(n28089), .IN2(n28265), .IN3(n28090), .IN4(n28271), .Q(
        n27864) );
  NAND4X0 U32024 ( .IN1(n27867), .IN2(n27866), .IN3(n27865), .IN4(n27864), 
        .QN(s1_data_o[11]) );
  OA22X1 U32025 ( .IN1(n28096), .IN2(n28283), .IN3(n28079), .IN4(n28281), .Q(
        n27871) );
  OA22X1 U32026 ( .IN1(n28091), .IN2(n28278), .IN3(n28101), .IN4(n28279), .Q(
        n27870) );
  OA22X1 U32027 ( .IN1(n28097), .IN2(n28280), .IN3(n28090), .IN4(n28282), .Q(
        n27869) );
  OA22X1 U32028 ( .IN1(n28098), .IN2(n28284), .IN3(n28099), .IN4(n28277), .Q(
        n27868) );
  NAND4X0 U32029 ( .IN1(n27871), .IN2(n27870), .IN3(n27869), .IN4(n27868), 
        .QN(s1_data_o[12]) );
  OA22X1 U32030 ( .IN1(n28090), .IN2(n28292), .IN3(n28101), .IN4(n28291), .Q(
        n27875) );
  OA22X1 U32031 ( .IN1(n28056), .IN2(n28290), .IN3(n28089), .IN4(n28296), .Q(
        n27874) );
  OA22X1 U32032 ( .IN1(n28088), .IN2(n28289), .IN3(n28099), .IN4(n28295), .Q(
        n27873) );
  OA22X1 U32033 ( .IN1(n28103), .IN2(n28294), .IN3(n28079), .IN4(n28293), .Q(
        n27872) );
  NAND4X0 U32034 ( .IN1(n27875), .IN2(n27874), .IN3(n27873), .IN4(n27872), 
        .QN(s1_data_o[13]) );
  OA22X1 U32035 ( .IN1(n28056), .IN2(n28306), .IN3(n28079), .IN4(n28302), .Q(
        n27879) );
  OA22X1 U32036 ( .IN1(n28089), .IN2(n28308), .IN3(n28101), .IN4(n28301), .Q(
        n27878) );
  OA22X1 U32037 ( .IN1(n28103), .IN2(n28304), .IN3(n28096), .IN4(n28307), .Q(
        n27877) );
  OA22X1 U32038 ( .IN1(n28090), .IN2(n28305), .IN3(n28099), .IN4(n28303), .Q(
        n27876) );
  NAND4X0 U32039 ( .IN1(n27879), .IN2(n27878), .IN3(n27877), .IN4(n27876), 
        .QN(s1_data_o[14]) );
  OA22X1 U32040 ( .IN1(n28103), .IN2(n28315), .IN3(n28101), .IN4(n28317), .Q(
        n27883) );
  OA22X1 U32041 ( .IN1(n28056), .IN2(n28316), .IN3(n28096), .IN4(n28320), .Q(
        n27882) );
  OA22X1 U32042 ( .IN1(n28090), .IN2(n28313), .IN3(n28099), .IN4(n28319), .Q(
        n27881) );
  OA22X1 U32043 ( .IN1(n28089), .IN2(n28314), .IN3(n28079), .IN4(n28318), .Q(
        n27880) );
  NAND4X0 U32044 ( .IN1(n27883), .IN2(n27882), .IN3(n27881), .IN4(n27880), 
        .QN(s1_data_o[15]) );
  OA22X1 U32045 ( .IN1(n28089), .IN2(n28331), .IN3(n28096), .IN4(n28329), .Q(
        n27887) );
  OA22X1 U32046 ( .IN1(n28102), .IN2(n28325), .IN3(n28099), .IN4(n28327), .Q(
        n27886) );
  OA22X1 U32047 ( .IN1(n28090), .IN2(n28326), .IN3(n28101), .IN4(n28328), .Q(
        n27885) );
  OA22X1 U32048 ( .IN1(n28056), .IN2(n28330), .IN3(n28091), .IN4(n28332), .Q(
        n27884) );
  NAND4X0 U32049 ( .IN1(n27887), .IN2(n27886), .IN3(n27885), .IN4(n27884), 
        .QN(s1_data_o[16]) );
  OA22X1 U32050 ( .IN1(n28088), .IN2(n28337), .IN3(n28079), .IN4(n28339), .Q(
        n27891) );
  OA22X1 U32051 ( .IN1(n28101), .IN2(n28343), .IN3(n28099), .IN4(n28341), .Q(
        n27890) );
  OA22X1 U32052 ( .IN1(n28089), .IN2(n28342), .IN3(n28090), .IN4(n28338), .Q(
        n27889) );
  OA22X1 U32053 ( .IN1(n28056), .IN2(n28340), .IN3(n28091), .IN4(n28344), .Q(
        n27888) );
  NAND4X0 U32054 ( .IN1(n27891), .IN2(n27890), .IN3(n27889), .IN4(n27888), 
        .QN(s1_data_o[17]) );
  OA22X1 U32055 ( .IN1(n28056), .IN2(n28352), .IN3(n28097), .IN4(n28350), .Q(
        n27895) );
  OA22X1 U32056 ( .IN1(n28100), .IN2(n28355), .IN3(n28099), .IN4(n28353), .Q(
        n27894) );
  OA22X1 U32057 ( .IN1(n28103), .IN2(n28356), .IN3(n28101), .IN4(n28351), .Q(
        n27893) );
  OA22X1 U32058 ( .IN1(n28096), .IN2(n28354), .IN3(n28102), .IN4(n28349), .Q(
        n27892) );
  NAND4X0 U32059 ( .IN1(n27895), .IN2(n27894), .IN3(n27893), .IN4(n27892), 
        .QN(s1_data_o[18]) );
  OA22X1 U32060 ( .IN1(n28089), .IN2(n28362), .IN3(n28101), .IN4(n28368), .Q(
        n27899) );
  OA22X1 U32061 ( .IN1(n28088), .IN2(n28365), .IN3(n28099), .IN4(n28367), .Q(
        n27898) );
  OA22X1 U32062 ( .IN1(n28056), .IN2(n28366), .IN3(n28090), .IN4(n28363), .Q(
        n27897) );
  OA22X1 U32063 ( .IN1(n28091), .IN2(n28364), .IN3(n28102), .IN4(n28361), .Q(
        n27896) );
  NAND4X0 U32064 ( .IN1(n27899), .IN2(n27898), .IN3(n27897), .IN4(n27896), 
        .QN(s1_data_o[19]) );
  OA22X1 U32065 ( .IN1(n28090), .IN2(n28373), .IN3(n28101), .IN4(n28379), .Q(
        n27903) );
  OA22X1 U32066 ( .IN1(n28103), .IN2(n28377), .IN3(n28096), .IN4(n28376), .Q(
        n27902) );
  OA22X1 U32067 ( .IN1(n28102), .IN2(n28380), .IN3(n28099), .IN4(n28375), .Q(
        n27901) );
  OA22X1 U32068 ( .IN1(n28056), .IN2(n28378), .IN3(n28097), .IN4(n28374), .Q(
        n27900) );
  NAND4X0 U32069 ( .IN1(n27903), .IN2(n27902), .IN3(n27901), .IN4(n27900), 
        .QN(s1_data_o[20]) );
  OA22X1 U32070 ( .IN1(n28090), .IN2(n28388), .IN3(n28099), .IN4(n28391), .Q(
        n27907) );
  OA22X1 U32071 ( .IN1(n28079), .IN2(n28385), .IN3(n28101), .IN4(n28389), .Q(
        n27906) );
  OA22X1 U32072 ( .IN1(n28056), .IN2(n28392), .IN3(n28089), .IN4(n28390), .Q(
        n27905) );
  OA22X1 U32073 ( .IN1(n28103), .IN2(n28386), .IN3(n28096), .IN4(n28387), .Q(
        n27904) );
  NAND4X0 U32074 ( .IN1(n27907), .IN2(n27906), .IN3(n27905), .IN4(n27904), 
        .QN(s1_data_o[21]) );
  OA22X1 U32075 ( .IN1(n28088), .IN2(n28398), .IN3(n28079), .IN4(n28399), .Q(
        n27911) );
  OA22X1 U32076 ( .IN1(n28101), .IN2(n28401), .IN3(n28099), .IN4(n28397), .Q(
        n27910) );
  OA22X1 U32077 ( .IN1(n28056), .IN2(n28400), .IN3(n28090), .IN4(n28403), .Q(
        n27909) );
  OA22X1 U32078 ( .IN1(n28103), .IN2(n28402), .IN3(n28097), .IN4(n28404), .Q(
        n27908) );
  NAND4X0 U32079 ( .IN1(n27911), .IN2(n27910), .IN3(n27909), .IN4(n27908), 
        .QN(s1_data_o[22]) );
  OA22X1 U32080 ( .IN1(n28056), .IN2(n28416), .IN3(n28096), .IN4(n28410), .Q(
        n27915) );
  OA22X1 U32081 ( .IN1(n28090), .IN2(n28413), .IN3(n28079), .IN4(n28412), .Q(
        n27914) );
  OA22X1 U32082 ( .IN1(n28089), .IN2(n28414), .IN3(n28099), .IN4(n28411), .Q(
        n27913) );
  OA22X1 U32083 ( .IN1(n28103), .IN2(n28415), .IN3(n28101), .IN4(n28409), .Q(
        n27912) );
  NAND4X0 U32084 ( .IN1(n27915), .IN2(n27914), .IN3(n27913), .IN4(n27912), 
        .QN(s1_data_o[23]) );
  OA22X1 U32085 ( .IN1(n28089), .IN2(n28422), .IN3(n28096), .IN4(n28425), .Q(
        n27919) );
  OA22X1 U32086 ( .IN1(n28056), .IN2(n28426), .IN3(n28101), .IN4(n28427), .Q(
        n27918) );
  OA22X1 U32087 ( .IN1(n28090), .IN2(n28421), .IN3(n28057), .IN4(n28423), .Q(
        n27917) );
  OA22X1 U32088 ( .IN1(n28103), .IN2(n28424), .IN3(n28102), .IN4(n28428), .Q(
        n27916) );
  NAND4X0 U32089 ( .IN1(n27919), .IN2(n27918), .IN3(n27917), .IN4(n27916), 
        .QN(s1_data_o[24]) );
  OA22X1 U32090 ( .IN1(n28056), .IN2(n28438), .IN3(n28091), .IN4(n28440), .Q(
        n27923) );
  OA22X1 U32091 ( .IN1(n28089), .IN2(n28434), .IN3(n28057), .IN4(n28435), .Q(
        n27922) );
  OA22X1 U32092 ( .IN1(n28088), .IN2(n28433), .IN3(n28079), .IN4(n28437), .Q(
        n27921) );
  OA22X1 U32093 ( .IN1(n28090), .IN2(n28439), .IN3(n28101), .IN4(n28436), .Q(
        n27920) );
  NAND4X0 U32094 ( .IN1(n27923), .IN2(n27922), .IN3(n27921), .IN4(n27920), 
        .QN(s1_data_o[25]) );
  OA22X1 U32095 ( .IN1(n28102), .IN2(n28448), .IN3(n28078), .IN4(n28447), .Q(
        n27927) );
  OA22X1 U32096 ( .IN1(n28089), .IN2(n28450), .IN3(n28090), .IN4(n28446), .Q(
        n27926) );
  OA22X1 U32097 ( .IN1(n28056), .IN2(n28452), .IN3(n28091), .IN4(n28451), .Q(
        n27925) );
  OA22X1 U32098 ( .IN1(n28088), .IN2(n28449), .IN3(n28057), .IN4(n28445), .Q(
        n27924) );
  NAND4X0 U32099 ( .IN1(n27927), .IN2(n27926), .IN3(n27925), .IN4(n27924), 
        .QN(s1_data_o[26]) );
  OA22X1 U32100 ( .IN1(n28056), .IN2(n28462), .IN3(n28078), .IN4(n28460), .Q(
        n27931) );
  OA22X1 U32101 ( .IN1(n28089), .IN2(n28464), .IN3(n28057), .IN4(n28459), .Q(
        n27930) );
  OA22X1 U32102 ( .IN1(n28103), .IN2(n28461), .IN3(n28096), .IN4(n28457), .Q(
        n27929) );
  OA22X1 U32103 ( .IN1(n28090), .IN2(n28458), .IN3(n28102), .IN4(n28463), .Q(
        n27928) );
  NAND4X0 U32104 ( .IN1(n27931), .IN2(n27930), .IN3(n27929), .IN4(n27928), 
        .QN(s1_data_o[27]) );
  OA22X1 U32105 ( .IN1(n28098), .IN2(n28474), .IN3(n28091), .IN4(n28476), .Q(
        n27935) );
  OA22X1 U32106 ( .IN1(n28088), .IN2(n28471), .IN3(n28057), .IN4(n28473), .Q(
        n27934) );
  OA22X1 U32107 ( .IN1(n28102), .IN2(n28475), .IN3(n28078), .IN4(n28469), .Q(
        n27933) );
  OA22X1 U32108 ( .IN1(n28089), .IN2(n28472), .IN3(n28100), .IN4(n28470), .Q(
        n27932) );
  NAND4X0 U32109 ( .IN1(n27935), .IN2(n27934), .IN3(n27933), .IN4(n27932), 
        .QN(s1_data_o[28]) );
  OA22X1 U32110 ( .IN1(n28103), .IN2(n28482), .IN3(n28089), .IN4(n28488), .Q(
        n27939) );
  OA22X1 U32111 ( .IN1(n28098), .IN2(n28484), .IN3(n28096), .IN4(n28487), .Q(
        n27938) );
  OA22X1 U32112 ( .IN1(n28090), .IN2(n28486), .IN3(n28057), .IN4(n28481), .Q(
        n27937) );
  OA22X1 U32113 ( .IN1(n28102), .IN2(n28483), .IN3(n28078), .IN4(n28485), .Q(
        n27936) );
  NAND4X0 U32114 ( .IN1(n27939), .IN2(n27938), .IN3(n27937), .IN4(n27936), 
        .QN(s1_data_o[29]) );
  OA22X1 U32115 ( .IN1(n28089), .IN2(n28497), .IN3(n28102), .IN4(n28495), .Q(
        n27943) );
  OA22X1 U32116 ( .IN1(n28088), .IN2(n28493), .IN3(n28078), .IN4(n28500), .Q(
        n27942) );
  OA22X1 U32117 ( .IN1(n28098), .IN2(n28494), .IN3(n28057), .IN4(n28499), .Q(
        n27941) );
  OA22X1 U32118 ( .IN1(n28103), .IN2(n28498), .IN3(n28100), .IN4(n28496), .Q(
        n27940) );
  NAND4X0 U32119 ( .IN1(n27943), .IN2(n27942), .IN3(n27941), .IN4(n27940), 
        .QN(s1_data_o[30]) );
  OA22X1 U32120 ( .IN1(n28102), .IN2(n28508), .IN3(n28057), .IN4(n28507), .Q(
        n27947) );
  OA22X1 U32121 ( .IN1(n28097), .IN2(n28506), .IN3(n28096), .IN4(n28512), .Q(
        n27946) );
  OA22X1 U32122 ( .IN1(n28098), .IN2(n28510), .IN3(n28100), .IN4(n28505), .Q(
        n27945) );
  OA22X1 U32123 ( .IN1(n28103), .IN2(n28509), .IN3(n28078), .IN4(n28511), .Q(
        n27944) );
  NAND4X0 U32124 ( .IN1(n27947), .IN2(n27946), .IN3(n27945), .IN4(n27944), 
        .QN(s1_data_o[31]) );
  OA22X1 U32125 ( .IN1(n28088), .IN2(n28523), .IN3(n28078), .IN4(n28521), .Q(
        n27951) );
  OA22X1 U32126 ( .IN1(n28097), .IN2(n28522), .IN3(n28057), .IN4(n28519), .Q(
        n27950) );
  OA22X1 U32127 ( .IN1(n28090), .IN2(n28524), .IN3(n28079), .IN4(n28520), .Q(
        n27949) );
  OA22X1 U32128 ( .IN1(n28098), .IN2(n28518), .IN3(n28091), .IN4(n28517), .Q(
        n27948) );
  NAND4X0 U32129 ( .IN1(n27951), .IN2(n27950), .IN3(n27949), .IN4(n27948), 
        .QN(s1_sel_o[0]) );
  OA22X1 U32130 ( .IN1(n28088), .IN2(n28535), .IN3(n28057), .IN4(n28529), .Q(
        n27955) );
  OA22X1 U32131 ( .IN1(n28097), .IN2(n28530), .IN3(n28079), .IN4(n28533), .Q(
        n27954) );
  OA22X1 U32132 ( .IN1(n28098), .IN2(n28534), .IN3(n28078), .IN4(n28531), .Q(
        n27953) );
  OA22X1 U32133 ( .IN1(n28103), .IN2(n28532), .IN3(n28100), .IN4(n28536), .Q(
        n27952) );
  NAND4X0 U32134 ( .IN1(n27955), .IN2(n27954), .IN3(n27953), .IN4(n27952), 
        .QN(s1_sel_o[1]) );
  OA22X1 U32135 ( .IN1(n28090), .IN2(n28548), .IN3(n28088), .IN4(n28547), .Q(
        n27959) );
  OA22X1 U32136 ( .IN1(n28091), .IN2(n28546), .IN3(n28097), .IN4(n28543), .Q(
        n27958) );
  OA22X1 U32137 ( .IN1(n28098), .IN2(n28544), .IN3(n28102), .IN4(n28542), .Q(
        n27957) );
  OA22X1 U32138 ( .IN1(n28101), .IN2(n28545), .IN3(n28057), .IN4(n28541), .Q(
        n27956) );
  NAND4X0 U32139 ( .IN1(n27959), .IN2(n27958), .IN3(n27957), .IN4(n27956), 
        .QN(s1_sel_o[2]) );
  OA22X1 U32140 ( .IN1(n28102), .IN2(n28560), .IN3(n28078), .IN4(n28559), .Q(
        n27963) );
  OA22X1 U32141 ( .IN1(n28097), .IN2(n28553), .IN3(n28057), .IN4(n28555), .Q(
        n27962) );
  OA22X1 U32142 ( .IN1(n28090), .IN2(n28557), .IN3(n28096), .IN4(n28556), .Q(
        n27961) );
  OA22X1 U32143 ( .IN1(n28098), .IN2(n28558), .IN3(n28091), .IN4(n28554), .Q(
        n27960) );
  NAND4X0 U32144 ( .IN1(n27963), .IN2(n27962), .IN3(n27961), .IN4(n27960), 
        .QN(s1_sel_o[3]) );
  OA22X1 U32145 ( .IN1(n28091), .IN2(n28570), .IN3(n28078), .IN4(n28565), .Q(
        n27967) );
  OA22X1 U32146 ( .IN1(n28090), .IN2(n28566), .IN3(n28088), .IN4(n28568), .Q(
        n27966) );
  OA22X1 U32147 ( .IN1(n28056), .IN2(n28572), .IN3(n28057), .IN4(n28569), .Q(
        n27965) );
  OA22X1 U32148 ( .IN1(n28089), .IN2(n28571), .IN3(n28079), .IN4(n28567), .Q(
        n27964) );
  NAND4X0 U32149 ( .IN1(n27967), .IN2(n27966), .IN3(n27965), .IN4(n27964), 
        .QN(s1_addr_o[0]) );
  OA22X1 U32150 ( .IN1(n28102), .IN2(n28584), .IN3(n28078), .IN4(n28577), .Q(
        n27971) );
  OA22X1 U32151 ( .IN1(n28088), .IN2(n28579), .IN3(n28057), .IN4(n28583), .Q(
        n27970) );
  OA22X1 U32152 ( .IN1(n28091), .IN2(n28578), .IN3(n28100), .IN4(n28581), .Q(
        n27969) );
  OA22X1 U32153 ( .IN1(n28056), .IN2(n28580), .IN3(n28097), .IN4(n28582), .Q(
        n27968) );
  NAND4X0 U32154 ( .IN1(n27971), .IN2(n27970), .IN3(n27969), .IN4(n27968), 
        .QN(s1_addr_o[1]) );
  OA22X1 U32155 ( .IN1(n28592), .IN2(n28100), .IN3(n28590), .IN4(n28088), .Q(
        n27975) );
  OA22X1 U32156 ( .IN1(n28589), .IN2(n28091), .IN3(n28595), .IN4(n28078), .Q(
        n27974) );
  OA22X1 U32157 ( .IN1(n28594), .IN2(n28089), .IN3(n28593), .IN4(n28079), .Q(
        n27973) );
  OA22X1 U32158 ( .IN1(n28596), .IN2(n28099), .IN3(n28591), .IN4(n28056), .Q(
        n27972) );
  NAND4X0 U32159 ( .IN1(n27975), .IN2(n27974), .IN3(n27973), .IN4(n27972), 
        .QN(s1_addr_o[2]) );
  OA22X1 U32160 ( .IN1(n28604), .IN2(n28097), .IN3(n28601), .IN4(n28056), .Q(
        n27979) );
  OA22X1 U32161 ( .IN1(n28602), .IN2(n28079), .IN3(n28605), .IN4(n28103), .Q(
        n27978) );
  OA22X1 U32162 ( .IN1(n28603), .IN2(n28101), .IN3(n28607), .IN4(n28100), .Q(
        n27977) );
  OA22X1 U32163 ( .IN1(n28606), .IN2(n28088), .IN3(n28608), .IN4(n28099), .Q(
        n27976) );
  NAND4X0 U32164 ( .IN1(n27979), .IN2(n27978), .IN3(n27977), .IN4(n27976), 
        .QN(s1_addr_o[3]) );
  OA22X1 U32165 ( .IN1(n28616), .IN2(n28091), .IN3(n28615), .IN4(n28096), .Q(
        n27983) );
  OA22X1 U32166 ( .IN1(n28618), .IN2(n28100), .IN3(n28613), .IN4(n28097), .Q(
        n27982) );
  OA22X1 U32167 ( .IN1(n28620), .IN2(n28101), .IN3(n28617), .IN4(n28098), .Q(
        n27981) );
  OA22X1 U32168 ( .IN1(n28619), .IN2(n28099), .IN3(n28614), .IN4(n28079), .Q(
        n27980) );
  NAND4X0 U32169 ( .IN1(n27983), .IN2(n27982), .IN3(n27981), .IN4(n27980), 
        .QN(s1_addr_o[4]) );
  OA22X1 U32170 ( .IN1(n28628), .IN2(n28101), .IN3(n28626), .IN4(n28100), .Q(
        n27987) );
  OA22X1 U32171 ( .IN1(n28631), .IN2(n28096), .IN3(n28630), .IN4(n28091), .Q(
        n27986) );
  OA22X1 U32172 ( .IN1(n28632), .IN2(n28097), .IN3(n28627), .IN4(n28079), .Q(
        n27985) );
  OA22X1 U32173 ( .IN1(n28625), .IN2(n28099), .IN3(n28629), .IN4(n28098), .Q(
        n27984) );
  NAND4X0 U32174 ( .IN1(n27987), .IN2(n27986), .IN3(n27985), .IN4(n27984), 
        .QN(s1_addr_o[5]) );
  OA22X1 U32175 ( .IN1(n28056), .IN2(n28642), .IN3(n28091), .IN4(n28640), .Q(
        n27991) );
  OA22X1 U32176 ( .IN1(n28090), .IN2(n28643), .IN3(n28078), .IN4(n28641), .Q(
        n27990) );
  OA22X1 U32177 ( .IN1(n28088), .IN2(n28638), .IN3(n28057), .IN4(n28639), .Q(
        n27989) );
  OA22X1 U32178 ( .IN1(n28097), .IN2(n28644), .IN3(n28102), .IN4(n28637), .Q(
        n27988) );
  NAND4X0 U32179 ( .IN1(n27991), .IN2(n27990), .IN3(n27989), .IN4(n27988), 
        .QN(s1_addr_o[6]) );
  OA22X1 U32180 ( .IN1(n28091), .IN2(n28652), .IN3(n28097), .IN4(n28656), .Q(
        n27995) );
  OA22X1 U32181 ( .IN1(n28090), .IN2(n28653), .IN3(n28078), .IN4(n28651), .Q(
        n27994) );
  OA22X1 U32182 ( .IN1(n28102), .IN2(n28649), .IN3(n28057), .IN4(n28655), .Q(
        n27993) );
  OA22X1 U32183 ( .IN1(n28098), .IN2(n28654), .IN3(n28096), .IN4(n28650), .Q(
        n27992) );
  NAND4X0 U32184 ( .IN1(n27995), .IN2(n27994), .IN3(n27993), .IN4(n27992), 
        .QN(s1_addr_o[7]) );
  OA22X1 U32185 ( .IN1(n28088), .IN2(n28668), .IN3(n28057), .IN4(n28667), .Q(
        n27999) );
  OA22X1 U32186 ( .IN1(n28056), .IN2(n28664), .IN3(n28089), .IN4(n28666), .Q(
        n27998) );
  OA22X1 U32187 ( .IN1(n28091), .IN2(n28663), .IN3(n28078), .IN4(n28661), .Q(
        n27997) );
  OA22X1 U32188 ( .IN1(n28090), .IN2(n28665), .IN3(n28079), .IN4(n28662), .Q(
        n27996) );
  NAND4X0 U32189 ( .IN1(n27999), .IN2(n27998), .IN3(n27997), .IN4(n27996), 
        .QN(s1_addr_o[8]) );
  OA22X1 U32190 ( .IN1(n28088), .IN2(n28673), .IN3(n28057), .IN4(n28677), .Q(
        n28003) );
  OA22X1 U32191 ( .IN1(n28103), .IN2(n28679), .IN3(n28100), .IN4(n28676), .Q(
        n28002) );
  OA22X1 U32192 ( .IN1(n28097), .IN2(n28674), .IN3(n28078), .IN4(n28675), .Q(
        n28001) );
  OA22X1 U32193 ( .IN1(n28098), .IN2(n28680), .IN3(n28102), .IN4(n28678), .Q(
        n28000) );
  NAND4X0 U32194 ( .IN1(n28003), .IN2(n28002), .IN3(n28001), .IN4(n28000), 
        .QN(s1_addr_o[9]) );
  OA22X1 U32195 ( .IN1(n28090), .IN2(n28687), .IN3(n28057), .IN4(n28689), .Q(
        n28007) );
  OA22X1 U32196 ( .IN1(n28102), .IN2(n28691), .IN3(n28078), .IN4(n28690), .Q(
        n28006) );
  OA22X1 U32197 ( .IN1(n28056), .IN2(n28692), .IN3(n28091), .IN4(n28686), .Q(
        n28005) );
  OA22X1 U32198 ( .IN1(n28089), .IN2(n28688), .IN3(n28088), .IN4(n28685), .Q(
        n28004) );
  NAND4X0 U32199 ( .IN1(n28007), .IN2(n28006), .IN3(n28005), .IN4(n28004), 
        .QN(s1_addr_o[10]) );
  OA22X1 U32200 ( .IN1(n28089), .IN2(n28697), .IN3(n28057), .IN4(n28699), .Q(
        n28011) );
  OA22X1 U32201 ( .IN1(n28090), .IN2(n28704), .IN3(n28088), .IN4(n28701), .Q(
        n28010) );
  OA22X1 U32202 ( .IN1(n28103), .IN2(n28698), .IN3(n28078), .IN4(n28700), .Q(
        n28009) );
  OA22X1 U32203 ( .IN1(n28098), .IN2(n28702), .IN3(n28102), .IN4(n28703), .Q(
        n28008) );
  NAND4X0 U32204 ( .IN1(n28011), .IN2(n28010), .IN3(n28009), .IN4(n28008), 
        .QN(s1_addr_o[11]) );
  OA22X1 U32205 ( .IN1(n28090), .IN2(n28716), .IN3(n28079), .IN4(n28715), .Q(
        n28015) );
  OA22X1 U32206 ( .IN1(n28091), .IN2(n28710), .IN3(n28057), .IN4(n28713), .Q(
        n28014) );
  OA22X1 U32207 ( .IN1(n28088), .IN2(n28709), .IN3(n28078), .IN4(n28711), .Q(
        n28013) );
  OA22X1 U32208 ( .IN1(n28098), .IN2(n28714), .IN3(n28097), .IN4(n28712), .Q(
        n28012) );
  NAND4X0 U32209 ( .IN1(n28015), .IN2(n28014), .IN3(n28013), .IN4(n28012), 
        .QN(s1_addr_o[12]) );
  OA22X1 U32210 ( .IN1(n28097), .IN2(n28726), .IN3(n28079), .IN4(n28721), .Q(
        n28019) );
  OA22X1 U32211 ( .IN1(n28056), .IN2(n28722), .IN3(n28096), .IN4(n28723), .Q(
        n28018) );
  OA22X1 U32212 ( .IN1(n28101), .IN2(n28725), .IN3(n28057), .IN4(n28727), .Q(
        n28017) );
  OA22X1 U32213 ( .IN1(n28091), .IN2(n28728), .IN3(n28100), .IN4(n28724), .Q(
        n28016) );
  NAND4X0 U32214 ( .IN1(n28019), .IN2(n28018), .IN3(n28017), .IN4(n28016), 
        .QN(s1_addr_o[13]) );
  OA22X1 U32215 ( .IN1(n28090), .IN2(n28735), .IN3(n28057), .IN4(n28739), .Q(
        n28023) );
  OA22X1 U32216 ( .IN1(n28056), .IN2(n28734), .IN3(n28078), .IN4(n28733), .Q(
        n28022) );
  OA22X1 U32217 ( .IN1(n28089), .IN2(n28736), .IN3(n28088), .IN4(n28740), .Q(
        n28021) );
  OA22X1 U32218 ( .IN1(n28091), .IN2(n28738), .IN3(n28079), .IN4(n28737), .Q(
        n28020) );
  NAND4X0 U32219 ( .IN1(n28023), .IN2(n28022), .IN3(n28021), .IN4(n28020), 
        .QN(s1_addr_o[14]) );
  OA22X1 U32220 ( .IN1(n28056), .IN2(n28746), .IN3(n28096), .IN4(n28747), .Q(
        n28027) );
  OA22X1 U32221 ( .IN1(n28102), .IN2(n28751), .IN3(n28057), .IN4(n28745), .Q(
        n28026) );
  OA22X1 U32222 ( .IN1(n28103), .IN2(n28748), .IN3(n28100), .IN4(n28752), .Q(
        n28025) );
  OA22X1 U32223 ( .IN1(n28089), .IN2(n28750), .IN3(n28078), .IN4(n28749), .Q(
        n28024) );
  NAND4X0 U32224 ( .IN1(n28027), .IN2(n28026), .IN3(n28025), .IN4(n28024), 
        .QN(s1_addr_o[15]) );
  OA22X1 U32225 ( .IN1(n28096), .IN2(n28759), .IN3(n28057), .IN4(n28763), .Q(
        n28031) );
  OA22X1 U32226 ( .IN1(n28098), .IN2(n28758), .IN3(n28078), .IN4(n28764), .Q(
        n28030) );
  OA22X1 U32227 ( .IN1(n28089), .IN2(n28760), .IN3(n28100), .IN4(n28761), .Q(
        n28029) );
  OA22X1 U32228 ( .IN1(n28103), .IN2(n28762), .IN3(n28102), .IN4(n28757), .Q(
        n28028) );
  NAND4X0 U32229 ( .IN1(n28031), .IN2(n28030), .IN3(n28029), .IN4(n28028), 
        .QN(s1_addr_o[16]) );
  OA22X1 U32230 ( .IN1(n28103), .IN2(n28776), .IN3(n28097), .IN4(n28774), .Q(
        n28035) );
  OA22X1 U32231 ( .IN1(n28088), .IN2(n28775), .IN3(n28057), .IN4(n28769), .Q(
        n28034) );
  OA22X1 U32232 ( .IN1(n28102), .IN2(n28771), .IN3(n28078), .IN4(n28770), .Q(
        n28033) );
  OA22X1 U32233 ( .IN1(n28056), .IN2(n28772), .IN3(n28100), .IN4(n28773), .Q(
        n28032) );
  NAND4X0 U32234 ( .IN1(n28035), .IN2(n28034), .IN3(n28033), .IN4(n28032), 
        .QN(s1_addr_o[17]) );
  OA22X1 U32235 ( .IN1(n28091), .IN2(n28788), .IN3(n28102), .IN4(n28783), .Q(
        n28039) );
  OA22X1 U32236 ( .IN1(n28090), .IN2(n28782), .IN3(n28078), .IN4(n28785), .Q(
        n28038) );
  OA22X1 U32237 ( .IN1(n28097), .IN2(n28787), .IN3(n28096), .IN4(n28784), .Q(
        n28037) );
  OA22X1 U32238 ( .IN1(n28098), .IN2(n28786), .IN3(n28057), .IN4(n28781), .Q(
        n28036) );
  NAND4X0 U32239 ( .IN1(n28039), .IN2(n28038), .IN3(n28037), .IN4(n28036), 
        .QN(s1_addr_o[18]) );
  OA22X1 U32240 ( .IN1(n28098), .IN2(n28796), .IN3(n28102), .IN4(n28795), .Q(
        n28043) );
  OA22X1 U32241 ( .IN1(n28090), .IN2(n28794), .IN3(n28096), .IN4(n28797), .Q(
        n28042) );
  OA22X1 U32242 ( .IN1(n28091), .IN2(n28800), .IN3(n28097), .IN4(n28798), .Q(
        n28041) );
  OA22X1 U32243 ( .IN1(n28101), .IN2(n28793), .IN3(n28057), .IN4(n28799), .Q(
        n28040) );
  NAND4X0 U32244 ( .IN1(n28043), .IN2(n28042), .IN3(n28041), .IN4(n28040), 
        .QN(s1_addr_o[19]) );
  OA22X1 U32245 ( .IN1(n28103), .IN2(n28808), .IN3(n28057), .IN4(n28805), .Q(
        n28047) );
  OA22X1 U32246 ( .IN1(n28088), .IN2(n28806), .IN3(n28078), .IN4(n28809), .Q(
        n28046) );
  OA22X1 U32247 ( .IN1(n28056), .IN2(n28812), .IN3(n28079), .IN4(n28811), .Q(
        n28045) );
  OA22X1 U32248 ( .IN1(n28097), .IN2(n28807), .IN3(n28090), .IN4(n28810), .Q(
        n28044) );
  NAND4X0 U32249 ( .IN1(n28047), .IN2(n28046), .IN3(n28045), .IN4(n28044), 
        .QN(s1_addr_o[20]) );
  OA22X1 U32250 ( .IN1(n28088), .IN2(n28821), .IN3(n28057), .IN4(n28817), .Q(
        n28051) );
  OA22X1 U32251 ( .IN1(n28091), .IN2(n28824), .IN3(n28090), .IN4(n28819), .Q(
        n28050) );
  OA22X1 U32252 ( .IN1(n28079), .IN2(n28823), .IN3(n28078), .IN4(n28818), .Q(
        n28049) );
  OA22X1 U32253 ( .IN1(n28056), .IN2(n28822), .IN3(n28097), .IN4(n28820), .Q(
        n28048) );
  NAND4X0 U32254 ( .IN1(n28051), .IN2(n28050), .IN3(n28049), .IN4(n28048), 
        .QN(s1_addr_o[21]) );
  OA22X1 U32255 ( .IN1(n28096), .IN2(n28836), .IN3(n28057), .IN4(n28829), .Q(
        n28055) );
  OA22X1 U32256 ( .IN1(n28103), .IN2(n28832), .IN3(n28097), .IN4(n28831), .Q(
        n28054) );
  OA22X1 U32257 ( .IN1(n28090), .IN2(n28838), .IN3(n28079), .IN4(n28834), .Q(
        n28053) );
  OA22X1 U32258 ( .IN1(n28098), .IN2(n28833), .IN3(n28078), .IN4(n28837), .Q(
        n28052) );
  NAND4X0 U32259 ( .IN1(n28055), .IN2(n28054), .IN3(n28053), .IN4(n28052), 
        .QN(s1_addr_o[22]) );
  OA22X1 U32260 ( .IN1(n28056), .IN2(n28848), .IN3(n28096), .IN4(n28852), .Q(
        n28061) );
  OA22X1 U32261 ( .IN1(n28103), .IN2(n28845), .IN3(n28102), .IN4(n28849), .Q(
        n28060) );
  OA22X1 U32262 ( .IN1(n28090), .IN2(n28850), .IN3(n28078), .IN4(n28846), .Q(
        n28059) );
  OA22X1 U32263 ( .IN1(n28097), .IN2(n28843), .IN3(n28057), .IN4(n28851), .Q(
        n28058) );
  NAND4X0 U32264 ( .IN1(n28061), .IN2(n28060), .IN3(n28059), .IN4(n28058), 
        .QN(s1_addr_o[23]) );
  OA22X1 U32265 ( .IN1(n28860), .IN2(n28099), .IN3(n28861), .IN4(n28088), .Q(
        n28065) );
  OA22X1 U32266 ( .IN1(n28864), .IN2(n28103), .IN3(n28857), .IN4(n28100), .Q(
        n28064) );
  OA22X1 U32267 ( .IN1(n28865), .IN2(n28101), .IN3(n28863), .IN4(n28098), .Q(
        n28063) );
  OA22X1 U32268 ( .IN1(n28858), .IN2(n28089), .IN3(n28859), .IN4(n28079), .Q(
        n28062) );
  NAND4X0 U32269 ( .IN1(n28065), .IN2(n28064), .IN3(n28063), .IN4(n28062), 
        .QN(s1_addr_o[24]) );
  OA22X1 U32270 ( .IN1(n28874), .IN2(n28100), .IN3(n28872), .IN4(n28096), .Q(
        n28069) );
  OA22X1 U32271 ( .IN1(n28877), .IN2(n28091), .IN3(n28876), .IN4(n28102), .Q(
        n28068) );
  OA22X1 U32272 ( .IN1(n28873), .IN2(n28097), .IN3(n28871), .IN4(n28078), .Q(
        n28067) );
  OA22X1 U32273 ( .IN1(n28875), .IN2(n28099), .IN3(n28870), .IN4(n28098), .Q(
        n28066) );
  NAND4X0 U32274 ( .IN1(n28069), .IN2(n28068), .IN3(n28067), .IN4(n28066), 
        .QN(s1_addr_o[25]) );
  OA22X1 U32275 ( .IN1(n28885), .IN2(n28089), .IN3(n28889), .IN4(n28099), .Q(
        n28073) );
  OA22X1 U32276 ( .IN1(n28883), .IN2(n28101), .IN3(n28884), .IN4(n28098), .Q(
        n28072) );
  OA22X1 U32277 ( .IN1(n28882), .IN2(n28100), .IN3(n28886), .IN4(n28096), .Q(
        n28071) );
  OA22X1 U32278 ( .IN1(n28887), .IN2(n28103), .IN3(n28888), .IN4(n28102), .Q(
        n28070) );
  NAND4X0 U32279 ( .IN1(n28073), .IN2(n28072), .IN3(n28071), .IN4(n28070), 
        .QN(s1_addr_o[26]) );
  OA22X1 U32280 ( .IN1(n28896), .IN2(n28102), .IN3(n28894), .IN4(n28098), .Q(
        n28077) );
  OA22X1 U32281 ( .IN1(n28899), .IN2(n28089), .IN3(n28897), .IN4(n28078), .Q(
        n28076) );
  OA22X1 U32282 ( .IN1(n28898), .IN2(n28099), .IN3(n28901), .IN4(n28100), .Q(
        n28075) );
  OA22X1 U32283 ( .IN1(n28895), .IN2(n28103), .IN3(n28900), .IN4(n28088), .Q(
        n28074) );
  NAND4X0 U32284 ( .IN1(n28077), .IN2(n28076), .IN3(n28075), .IN4(n28074), 
        .QN(s1_addr_o[27]) );
  OA22X1 U32285 ( .IN1(n28908), .IN2(n28100), .IN3(n28906), .IN4(n28088), .Q(
        n28083) );
  OA22X1 U32286 ( .IN1(n28909), .IN2(n28097), .IN3(n28907), .IN4(n28078), .Q(
        n28082) );
  OA22X1 U32287 ( .IN1(n28911), .IN2(n28091), .IN3(n28913), .IN4(n28099), .Q(
        n28081) );
  OA22X1 U32288 ( .IN1(n28910), .IN2(n28079), .IN3(n28912), .IN4(n28098), .Q(
        n28080) );
  NAND4X0 U32289 ( .IN1(n28083), .IN2(n28082), .IN3(n28081), .IN4(n28080), 
        .QN(s1_addr_o[28]) );
  OA22X1 U32290 ( .IN1(n28920), .IN2(n28102), .IN3(n28919), .IN4(n28100), .Q(
        n28087) );
  OA22X1 U32291 ( .IN1(n28922), .IN2(n28101), .IN3(n28925), .IN4(n28098), .Q(
        n28086) );
  OA22X1 U32292 ( .IN1(n28921), .IN2(n28099), .IN3(n28923), .IN4(n28096), .Q(
        n28085) );
  OA22X1 U32293 ( .IN1(n28926), .IN2(n28097), .IN3(n28924), .IN4(n28091), .Q(
        n28084) );
  NAND4X0 U32294 ( .IN1(n28087), .IN2(n28086), .IN3(n28085), .IN4(n28084), 
        .QN(s1_addr_o[29]) );
  OA22X1 U32295 ( .IN1(n28932), .IN2(n28089), .IN3(n28939), .IN4(n28088), .Q(
        n28095) );
  OA22X1 U32296 ( .IN1(n28933), .IN2(n28099), .IN3(n28936), .IN4(n28102), .Q(
        n28094) );
  OA22X1 U32297 ( .IN1(n28935), .IN2(n28091), .IN3(n28940), .IN4(n28090), .Q(
        n28093) );
  OA22X1 U32298 ( .IN1(n28937), .IN2(n28101), .IN3(n28931), .IN4(n28098), .Q(
        n28092) );
  NAND4X0 U32299 ( .IN1(n28095), .IN2(n28094), .IN3(n28093), .IN4(n28092), 
        .QN(s1_addr_o[30]) );
  OA22X1 U32300 ( .IN1(n28948), .IN2(n28097), .IN3(n28946), .IN4(n28096), .Q(
        n28107) );
  OA22X1 U32301 ( .IN1(n28960), .IN2(n28099), .IN3(n28950), .IN4(n28098), .Q(
        n28106) );
  OA22X1 U32302 ( .IN1(n28956), .IN2(n28101), .IN3(n28958), .IN4(n28100), .Q(
        n28105) );
  OA22X1 U32303 ( .IN1(n28952), .IN2(n28103), .IN3(n28954), .IN4(n28102), .Q(
        n28104) );
  NAND4X0 U32304 ( .IN1(n28107), .IN2(n28106), .IN3(n28105), .IN4(n28104), 
        .QN(s1_addr_o[31]) );
  OA22X1 U32305 ( .IN1(n29273), .IN2(n28109), .IN3(n29330), .IN4(n28108), .Q(
        n28120) );
  OA22X1 U32306 ( .IN1(n29368), .IN2(n28111), .IN3(n29292), .IN4(n28110), .Q(
        n28119) );
  INVX0 U32307 ( .INP(n28112), .ZN(n28113) );
  OA22X1 U32308 ( .IN1(n29349), .IN2(n28114), .IN3(n29235), .IN4(n28113), .Q(
        n28118) );
  OA22X1 U32309 ( .IN1(n29254), .IN2(n28116), .IN3(n29311), .IN4(n28115), .Q(
        n28117) );
  NAND4X0 U32310 ( .IN1(n28120), .IN2(n28119), .IN3(n28118), .IN4(n28117), 
        .QN(s0_stb_o) );
  INVX0 U32311 ( .INP(n28973), .ZN(n28945) );
  INVX0 U32312 ( .INP(n28830), .ZN(n28976) );
  INVX0 U32313 ( .INP(n28976), .ZN(n28959) );
  OA22X1 U32314 ( .IN1(n28945), .IN2(n28122), .IN3(n28959), .IN4(n28121), .Q(
        n28132) );
  INVX0 U32315 ( .INP(n28974), .ZN(n28862) );
  INVX0 U32316 ( .INP(n28975), .ZN(n28844) );
  OA22X1 U32317 ( .IN1(n28862), .IN2(n28124), .IN3(n28844), .IN4(n28123), .Q(
        n28131) );
  INVX0 U32318 ( .INP(n28967), .ZN(n28918) );
  INVX0 U32319 ( .INP(n28965), .ZN(n28835) );
  OA22X1 U32320 ( .IN1(n28918), .IN2(n28126), .IN3(n28835), .IN4(n28125), .Q(
        n28130) );
  INVX0 U32321 ( .INP(n28968), .ZN(n28951) );
  OA22X1 U32322 ( .IN1(n28951), .IN2(n28128), .IN3(n28847), .IN4(n28127), .Q(
        n28129) );
  NAND4X0 U32323 ( .IN1(n28132), .IN2(n28131), .IN3(n28130), .IN4(n28129), 
        .QN(s0_we_o) );
  OA22X1 U32324 ( .IN1(n28949), .IN2(n28134), .IN3(n28844), .IN4(n28133), .Q(
        n28144) );
  OA22X1 U32325 ( .IN1(n28835), .IN2(n28136), .IN3(n28830), .IN4(n28135), .Q(
        n28143) );
  INVX0 U32326 ( .INP(n28973), .ZN(n28938) );
  OA22X1 U32327 ( .IN1(n28938), .IN2(n28138), .IN3(n28847), .IN4(n28137), .Q(
        n28142) );
  INVX0 U32328 ( .INP(n28968), .ZN(n28934) );
  OA22X1 U32329 ( .IN1(n28934), .IN2(n28140), .IN3(n28918), .IN4(n28139), .Q(
        n28141) );
  NAND4X0 U32330 ( .IN1(n28144), .IN2(n28143), .IN3(n28142), .IN4(n28141), 
        .QN(s0_data_o[0]) );
  OA22X1 U32331 ( .IN1(n28934), .IN2(n28146), .IN3(n28918), .IN4(n28145), .Q(
        n28156) );
  INVX0 U32332 ( .INP(n28975), .ZN(n28947) );
  OA22X1 U32333 ( .IN1(n28947), .IN2(n28148), .IN3(n28830), .IN4(n28147), .Q(
        n28155) );
  OA22X1 U32334 ( .IN1(n28862), .IN2(n28150), .IN3(n28945), .IN4(n28149), .Q(
        n28154) );
  OA22X1 U32335 ( .IN1(n28835), .IN2(n28152), .IN3(n28847), .IN4(n28151), .Q(
        n28153) );
  NAND4X0 U32336 ( .IN1(n28156), .IN2(n28155), .IN3(n28154), .IN4(n28153), 
        .QN(s0_data_o[1]) );
  OA22X1 U32337 ( .IN1(n28945), .IN2(n28158), .IN3(n28847), .IN4(n28157), .Q(
        n28168) );
  OA22X1 U32338 ( .IN1(n28949), .IN2(n28160), .IN3(n28918), .IN4(n28159), .Q(
        n28167) );
  INVX0 U32339 ( .INP(n28965), .ZN(n28953) );
  OA22X1 U32340 ( .IN1(n28953), .IN2(n28162), .IN3(n28830), .IN4(n28161), .Q(
        n28166) );
  OA22X1 U32341 ( .IN1(n28934), .IN2(n28164), .IN3(n28844), .IN4(n28163), .Q(
        n28165) );
  NAND4X0 U32342 ( .IN1(n28168), .IN2(n28167), .IN3(n28166), .IN4(n28165), 
        .QN(s0_data_o[2]) );
  OA22X1 U32343 ( .IN1(n28918), .IN2(n28170), .IN3(n28847), .IN4(n28169), .Q(
        n28180) );
  OA22X1 U32344 ( .IN1(n28862), .IN2(n28172), .IN3(n28945), .IN4(n28171), .Q(
        n28179) );
  OA22X1 U32345 ( .IN1(n28934), .IN2(n28174), .IN3(n28830), .IN4(n28173), .Q(
        n28178) );
  OA22X1 U32346 ( .IN1(n28844), .IN2(n28176), .IN3(n28835), .IN4(n28175), .Q(
        n28177) );
  NAND4X0 U32347 ( .IN1(n28180), .IN2(n28179), .IN3(n28178), .IN4(n28177), 
        .QN(s0_data_o[3]) );
  OA22X1 U32348 ( .IN1(n28949), .IN2(n28182), .IN3(n28830), .IN4(n28181), .Q(
        n28192) );
  OA22X1 U32349 ( .IN1(n28934), .IN2(n28184), .IN3(n28835), .IN4(n28183), .Q(
        n28191) );
  OA22X1 U32350 ( .IN1(n28947), .IN2(n28186), .IN3(n28945), .IN4(n28185), .Q(
        n28190) );
  OA22X1 U32351 ( .IN1(n28918), .IN2(n28188), .IN3(n28847), .IN4(n28187), .Q(
        n28189) );
  NAND4X0 U32352 ( .IN1(n28192), .IN2(n28191), .IN3(n28190), .IN4(n28189), 
        .QN(s0_data_o[4]) );
  OA22X1 U32353 ( .IN1(n28844), .IN2(n28194), .IN3(n28918), .IN4(n28193), .Q(
        n28204) );
  OA22X1 U32354 ( .IN1(n28862), .IN2(n28196), .IN3(n28847), .IN4(n28195), .Q(
        n28203) );
  OA22X1 U32355 ( .IN1(n28938), .IN2(n28198), .IN3(n28835), .IN4(n28197), .Q(
        n28202) );
  OA22X1 U32356 ( .IN1(n28934), .IN2(n28200), .IN3(n28830), .IN4(n28199), .Q(
        n28201) );
  NAND4X0 U32357 ( .IN1(n28204), .IN2(n28203), .IN3(n28202), .IN4(n28201), 
        .QN(s0_data_o[5]) );
  OA22X1 U32358 ( .IN1(n28844), .IN2(n28206), .IN3(n28835), .IN4(n28205), .Q(
        n28216) );
  OA22X1 U32359 ( .IN1(n28949), .IN2(n28208), .IN3(n28951), .IN4(n28207), .Q(
        n28215) );
  INVX0 U32360 ( .INP(n28847), .ZN(n28966) );
  INVX0 U32361 ( .INP(n28966), .ZN(n28955) );
  OA22X1 U32362 ( .IN1(n28955), .IN2(n28210), .IN3(n28830), .IN4(n28209), .Q(
        n28214) );
  INVX0 U32363 ( .INP(n28967), .ZN(n28957) );
  OA22X1 U32364 ( .IN1(n28957), .IN2(n28212), .IN3(n28945), .IN4(n28211), .Q(
        n28213) );
  NAND4X0 U32365 ( .IN1(n28216), .IN2(n28215), .IN3(n28214), .IN4(n28213), 
        .QN(s0_data_o[6]) );
  OA22X1 U32366 ( .IN1(n28957), .IN2(n28218), .IN3(n28945), .IN4(n28217), .Q(
        n28228) );
  OA22X1 U32367 ( .IN1(n28862), .IN2(n28220), .IN3(n28951), .IN4(n28219), .Q(
        n28227) );
  OA22X1 U32368 ( .IN1(n28955), .IN2(n28222), .IN3(n28959), .IN4(n28221), .Q(
        n28226) );
  OA22X1 U32369 ( .IN1(n28947), .IN2(n28224), .IN3(n28835), .IN4(n28223), .Q(
        n28225) );
  NAND4X0 U32370 ( .IN1(n28228), .IN2(n28227), .IN3(n28226), .IN4(n28225), 
        .QN(s0_data_o[7]) );
  OA22X1 U32371 ( .IN1(n28862), .IN2(n28230), .IN3(n28835), .IN4(n28229), .Q(
        n28240) );
  OA22X1 U32372 ( .IN1(n28934), .IN2(n28232), .IN3(n28844), .IN4(n28231), .Q(
        n28239) );
  OA22X1 U32373 ( .IN1(n28957), .IN2(n28234), .IN3(n28847), .IN4(n28233), .Q(
        n28238) );
  OA22X1 U32374 ( .IN1(n28945), .IN2(n28236), .IN3(n28959), .IN4(n28235), .Q(
        n28237) );
  NAND4X0 U32375 ( .IN1(n28240), .IN2(n28239), .IN3(n28238), .IN4(n28237), 
        .QN(s0_data_o[8]) );
  OA22X1 U32376 ( .IN1(n28949), .IN2(n28242), .IN3(n28945), .IN4(n28241), .Q(
        n28252) );
  OA22X1 U32377 ( .IN1(n28934), .IN2(n28244), .IN3(n28847), .IN4(n28243), .Q(
        n28251) );
  OA22X1 U32378 ( .IN1(n28947), .IN2(n28246), .IN3(n28835), .IN4(n28245), .Q(
        n28250) );
  OA22X1 U32379 ( .IN1(n28918), .IN2(n28248), .IN3(n28959), .IN4(n28247), .Q(
        n28249) );
  NAND4X0 U32380 ( .IN1(n28252), .IN2(n28251), .IN3(n28250), .IN4(n28249), 
        .QN(s0_data_o[9]) );
  OA22X1 U32381 ( .IN1(n28938), .IN2(n28254), .IN3(n28847), .IN4(n28253), .Q(
        n28264) );
  OA22X1 U32382 ( .IN1(n28957), .IN2(n28256), .IN3(n28835), .IN4(n28255), .Q(
        n28263) );
  OA22X1 U32383 ( .IN1(n28862), .IN2(n28258), .IN3(n28951), .IN4(n28257), .Q(
        n28262) );
  OA22X1 U32384 ( .IN1(n28844), .IN2(n28260), .IN3(n28959), .IN4(n28259), .Q(
        n28261) );
  NAND4X0 U32385 ( .IN1(n28264), .IN2(n28263), .IN3(n28262), .IN4(n28261), 
        .QN(s0_data_o[10]) );
  OA22X1 U32386 ( .IN1(n28949), .IN2(n28266), .IN3(n28844), .IN4(n28265), .Q(
        n28276) );
  OA22X1 U32387 ( .IN1(n28945), .IN2(n28268), .IN3(n28955), .IN4(n28267), .Q(
        n28275) );
  OA22X1 U32388 ( .IN1(n28835), .IN2(n28270), .IN3(n28959), .IN4(n28269), .Q(
        n28274) );
  OA22X1 U32389 ( .IN1(n28934), .IN2(n28272), .IN3(n28918), .IN4(n28271), .Q(
        n28273) );
  NAND4X0 U32390 ( .IN1(n28276), .IN2(n28275), .IN3(n28274), .IN4(n28273), 
        .QN(s0_data_o[11]) );
  OA22X1 U32391 ( .IN1(n28934), .IN2(n28278), .IN3(n28959), .IN4(n28277), .Q(
        n28288) );
  OA22X1 U32392 ( .IN1(n28844), .IN2(n28280), .IN3(n28955), .IN4(n28279), .Q(
        n28287) );
  OA22X1 U32393 ( .IN1(n28918), .IN2(n28282), .IN3(n28835), .IN4(n28281), .Q(
        n28286) );
  OA22X1 U32394 ( .IN1(n28862), .IN2(n28284), .IN3(n28945), .IN4(n28283), .Q(
        n28285) );
  NAND4X0 U32395 ( .IN1(n28288), .IN2(n28287), .IN3(n28286), .IN4(n28285), 
        .QN(s0_data_o[12]) );
  OA22X1 U32396 ( .IN1(n28949), .IN2(n28290), .IN3(n28945), .IN4(n28289), .Q(
        n28300) );
  OA22X1 U32397 ( .IN1(n28957), .IN2(n28292), .IN3(n28955), .IN4(n28291), .Q(
        n28299) );
  OA22X1 U32398 ( .IN1(n28951), .IN2(n28294), .IN3(n28835), .IN4(n28293), .Q(
        n28298) );
  OA22X1 U32399 ( .IN1(n28947), .IN2(n28296), .IN3(n28959), .IN4(n28295), .Q(
        n28297) );
  NAND4X0 U32400 ( .IN1(n28300), .IN2(n28299), .IN3(n28298), .IN4(n28297), 
        .QN(s0_data_o[13]) );
  OA22X1 U32401 ( .IN1(n28953), .IN2(n28302), .IN3(n28955), .IN4(n28301), .Q(
        n28312) );
  OA22X1 U32402 ( .IN1(n28934), .IN2(n28304), .IN3(n28959), .IN4(n28303), .Q(
        n28311) );
  OA22X1 U32403 ( .IN1(n28862), .IN2(n28306), .IN3(n28918), .IN4(n28305), .Q(
        n28310) );
  OA22X1 U32404 ( .IN1(n28844), .IN2(n28308), .IN3(n28945), .IN4(n28307), .Q(
        n28309) );
  NAND4X0 U32405 ( .IN1(n28312), .IN2(n28311), .IN3(n28310), .IN4(n28309), 
        .QN(s0_data_o[14]) );
  OA22X1 U32406 ( .IN1(n28844), .IN2(n28314), .IN3(n28957), .IN4(n28313), .Q(
        n28324) );
  OA22X1 U32407 ( .IN1(n28862), .IN2(n28316), .IN3(n28951), .IN4(n28315), .Q(
        n28323) );
  OA22X1 U32408 ( .IN1(n28835), .IN2(n28318), .IN3(n28955), .IN4(n28317), .Q(
        n28322) );
  OA22X1 U32409 ( .IN1(n28938), .IN2(n28320), .IN3(n28959), .IN4(n28319), .Q(
        n28321) );
  NAND4X0 U32410 ( .IN1(n28324), .IN2(n28323), .IN3(n28322), .IN4(n28321), 
        .QN(s0_data_o[15]) );
  OA22X1 U32411 ( .IN1(n28918), .IN2(n28326), .IN3(n28835), .IN4(n28325), .Q(
        n28336) );
  OA22X1 U32412 ( .IN1(n28847), .IN2(n28328), .IN3(n28959), .IN4(n28327), .Q(
        n28335) );
  OA22X1 U32413 ( .IN1(n28862), .IN2(n28330), .IN3(n28938), .IN4(n28329), .Q(
        n28334) );
  OA22X1 U32414 ( .IN1(n28934), .IN2(n28332), .IN3(n28844), .IN4(n28331), .Q(
        n28333) );
  NAND4X0 U32415 ( .IN1(n28336), .IN2(n28335), .IN3(n28334), .IN4(n28333), 
        .QN(s0_data_o[16]) );
  OA22X1 U32416 ( .IN1(n28957), .IN2(n28338), .IN3(n28945), .IN4(n28337), .Q(
        n28348) );
  OA22X1 U32417 ( .IN1(n28862), .IN2(n28340), .IN3(n28835), .IN4(n28339), .Q(
        n28347) );
  OA22X1 U32418 ( .IN1(n28947), .IN2(n28342), .IN3(n28959), .IN4(n28341), .Q(
        n28346) );
  OA22X1 U32419 ( .IN1(n28934), .IN2(n28344), .IN3(n28955), .IN4(n28343), .Q(
        n28345) );
  NAND4X0 U32420 ( .IN1(n28348), .IN2(n28347), .IN3(n28346), .IN4(n28345), 
        .QN(s0_data_o[17]) );
  OA22X1 U32421 ( .IN1(n28947), .IN2(n28350), .IN3(n28835), .IN4(n28349), .Q(
        n28360) );
  OA22X1 U32422 ( .IN1(n28862), .IN2(n28352), .IN3(n28955), .IN4(n28351), .Q(
        n28359) );
  OA22X1 U32423 ( .IN1(n28945), .IN2(n28354), .IN3(n28959), .IN4(n28353), .Q(
        n28358) );
  OA22X1 U32424 ( .IN1(n28934), .IN2(n28356), .IN3(n28918), .IN4(n28355), .Q(
        n28357) );
  NAND4X0 U32425 ( .IN1(n28360), .IN2(n28359), .IN3(n28358), .IN4(n28357), 
        .QN(s0_data_o[18]) );
  OA22X1 U32426 ( .IN1(n28844), .IN2(n28362), .IN3(n28835), .IN4(n28361), .Q(
        n28372) );
  OA22X1 U32427 ( .IN1(n28951), .IN2(n28364), .IN3(n28957), .IN4(n28363), .Q(
        n28371) );
  OA22X1 U32428 ( .IN1(n28862), .IN2(n28366), .IN3(n28938), .IN4(n28365), .Q(
        n28370) );
  OA22X1 U32429 ( .IN1(n28847), .IN2(n28368), .IN3(n28959), .IN4(n28367), .Q(
        n28369) );
  NAND4X0 U32430 ( .IN1(n28372), .IN2(n28371), .IN3(n28370), .IN4(n28369), 
        .QN(s0_data_o[19]) );
  OA22X1 U32431 ( .IN1(n28947), .IN2(n28374), .IN3(n28918), .IN4(n28373), .Q(
        n28384) );
  OA22X1 U32432 ( .IN1(n28938), .IN2(n28376), .IN3(n28959), .IN4(n28375), .Q(
        n28383) );
  OA22X1 U32433 ( .IN1(n28862), .IN2(n28378), .IN3(n28951), .IN4(n28377), .Q(
        n28382) );
  OA22X1 U32434 ( .IN1(n28953), .IN2(n28380), .IN3(n28955), .IN4(n28379), .Q(
        n28381) );
  NAND4X0 U32435 ( .IN1(n28384), .IN2(n28383), .IN3(n28382), .IN4(n28381), 
        .QN(s0_data_o[20]) );
  OA22X1 U32436 ( .IN1(n28934), .IN2(n28386), .IN3(n28835), .IN4(n28385), .Q(
        n28396) );
  OA22X1 U32437 ( .IN1(n28957), .IN2(n28388), .IN3(n28938), .IN4(n28387), .Q(
        n28395) );
  OA22X1 U32438 ( .IN1(n28844), .IN2(n28390), .IN3(n28955), .IN4(n28389), .Q(
        n28394) );
  OA22X1 U32439 ( .IN1(n28862), .IN2(n28392), .IN3(n28959), .IN4(n28391), .Q(
        n28393) );
  NAND4X0 U32440 ( .IN1(n28396), .IN2(n28395), .IN3(n28394), .IN4(n28393), 
        .QN(s0_data_o[21]) );
  OA22X1 U32441 ( .IN1(n28938), .IN2(n28398), .IN3(n28959), .IN4(n28397), .Q(
        n28408) );
  OA22X1 U32442 ( .IN1(n28862), .IN2(n28400), .IN3(n28835), .IN4(n28399), .Q(
        n28407) );
  OA22X1 U32443 ( .IN1(n28951), .IN2(n28402), .IN3(n28955), .IN4(n28401), .Q(
        n28406) );
  OA22X1 U32444 ( .IN1(n28844), .IN2(n28404), .IN3(n28918), .IN4(n28403), .Q(
        n28405) );
  NAND4X0 U32445 ( .IN1(n28408), .IN2(n28407), .IN3(n28406), .IN4(n28405), 
        .QN(s0_data_o[22]) );
  OA22X1 U32446 ( .IN1(n28938), .IN2(n28410), .IN3(n28955), .IN4(n28409), .Q(
        n28420) );
  OA22X1 U32447 ( .IN1(n28953), .IN2(n28412), .IN3(n28830), .IN4(n28411), .Q(
        n28419) );
  OA22X1 U32448 ( .IN1(n28947), .IN2(n28414), .IN3(n28957), .IN4(n28413), .Q(
        n28418) );
  OA22X1 U32449 ( .IN1(n28862), .IN2(n28416), .IN3(n28951), .IN4(n28415), .Q(
        n28417) );
  NAND4X0 U32450 ( .IN1(n28420), .IN2(n28419), .IN3(n28418), .IN4(n28417), 
        .QN(s0_data_o[23]) );
  OA22X1 U32451 ( .IN1(n28844), .IN2(n28422), .IN3(n28918), .IN4(n28421), .Q(
        n28432) );
  OA22X1 U32452 ( .IN1(n28934), .IN2(n28424), .IN3(n28830), .IN4(n28423), .Q(
        n28431) );
  OA22X1 U32453 ( .IN1(n28862), .IN2(n28426), .IN3(n28945), .IN4(n28425), .Q(
        n28430) );
  OA22X1 U32454 ( .IN1(n28953), .IN2(n28428), .IN3(n28955), .IN4(n28427), .Q(
        n28429) );
  NAND4X0 U32455 ( .IN1(n28432), .IN2(n28431), .IN3(n28430), .IN4(n28429), 
        .QN(s0_data_o[24]) );
  OA22X1 U32456 ( .IN1(n28947), .IN2(n28434), .IN3(n28945), .IN4(n28433), .Q(
        n28444) );
  OA22X1 U32457 ( .IN1(n28847), .IN2(n28436), .IN3(n28830), .IN4(n28435), .Q(
        n28443) );
  OA22X1 U32458 ( .IN1(n28862), .IN2(n28438), .IN3(n28953), .IN4(n28437), .Q(
        n28442) );
  OA22X1 U32459 ( .IN1(n28934), .IN2(n28440), .IN3(n28957), .IN4(n28439), .Q(
        n28441) );
  NAND4X0 U32460 ( .IN1(n28444), .IN2(n28443), .IN3(n28442), .IN4(n28441), 
        .QN(s0_data_o[25]) );
  OA22X1 U32461 ( .IN1(n28957), .IN2(n28446), .IN3(n28830), .IN4(n28445), .Q(
        n28456) );
  OA22X1 U32462 ( .IN1(n28835), .IN2(n28448), .IN3(n28955), .IN4(n28447), .Q(
        n28455) );
  OA22X1 U32463 ( .IN1(n28844), .IN2(n28450), .IN3(n28938), .IN4(n28449), .Q(
        n28454) );
  OA22X1 U32464 ( .IN1(n28862), .IN2(n28452), .IN3(n28951), .IN4(n28451), .Q(
        n28453) );
  NAND4X0 U32465 ( .IN1(n28456), .IN2(n28455), .IN3(n28454), .IN4(n28453), 
        .QN(s0_data_o[26]) );
  OA22X1 U32466 ( .IN1(n28957), .IN2(n28458), .IN3(n28945), .IN4(n28457), .Q(
        n28468) );
  OA22X1 U32467 ( .IN1(n28847), .IN2(n28460), .IN3(n28830), .IN4(n28459), .Q(
        n28467) );
  OA22X1 U32468 ( .IN1(n28862), .IN2(n28462), .IN3(n28951), .IN4(n28461), .Q(
        n28466) );
  OA22X1 U32469 ( .IN1(n28947), .IN2(n28464), .IN3(n28835), .IN4(n28463), .Q(
        n28465) );
  NAND4X0 U32470 ( .IN1(n28468), .IN2(n28467), .IN3(n28466), .IN4(n28465), 
        .QN(s0_data_o[27]) );
  OA22X1 U32471 ( .IN1(n28957), .IN2(n28470), .IN3(n28955), .IN4(n28469), .Q(
        n28480) );
  OA22X1 U32472 ( .IN1(n28947), .IN2(n28472), .IN3(n28945), .IN4(n28471), .Q(
        n28479) );
  OA22X1 U32473 ( .IN1(n28949), .IN2(n28474), .IN3(n28830), .IN4(n28473), .Q(
        n28478) );
  OA22X1 U32474 ( .IN1(n28951), .IN2(n28476), .IN3(n28953), .IN4(n28475), .Q(
        n28477) );
  NAND4X0 U32475 ( .IN1(n28480), .IN2(n28479), .IN3(n28478), .IN4(n28477), 
        .QN(s0_data_o[28]) );
  OA22X1 U32476 ( .IN1(n28934), .IN2(n28482), .IN3(n28830), .IN4(n28481), .Q(
        n28492) );
  OA22X1 U32477 ( .IN1(n28949), .IN2(n28484), .IN3(n28835), .IN4(n28483), .Q(
        n28491) );
  OA22X1 U32478 ( .IN1(n28957), .IN2(n28486), .IN3(n28955), .IN4(n28485), .Q(
        n28490) );
  OA22X1 U32479 ( .IN1(n28844), .IN2(n28488), .IN3(n28945), .IN4(n28487), .Q(
        n28489) );
  NAND4X0 U32480 ( .IN1(n28492), .IN2(n28491), .IN3(n28490), .IN4(n28489), 
        .QN(s0_data_o[29]) );
  OA22X1 U32481 ( .IN1(n28949), .IN2(n28494), .IN3(n28938), .IN4(n28493), .Q(
        n28504) );
  OA22X1 U32482 ( .IN1(n28957), .IN2(n28496), .IN3(n28953), .IN4(n28495), .Q(
        n28503) );
  OA22X1 U32483 ( .IN1(n28951), .IN2(n28498), .IN3(n28844), .IN4(n28497), .Q(
        n28502) );
  OA22X1 U32484 ( .IN1(n28847), .IN2(n28500), .IN3(n28830), .IN4(n28499), .Q(
        n28501) );
  NAND4X0 U32485 ( .IN1(n28504), .IN2(n28503), .IN3(n28502), .IN4(n28501), 
        .QN(s0_data_o[30]) );
  OA22X1 U32486 ( .IN1(n28844), .IN2(n28506), .IN3(n28918), .IN4(n28505), .Q(
        n28516) );
  OA22X1 U32487 ( .IN1(n28953), .IN2(n28508), .IN3(n28830), .IN4(n28507), .Q(
        n28515) );
  OA22X1 U32488 ( .IN1(n28949), .IN2(n28510), .IN3(n28951), .IN4(n28509), .Q(
        n28514) );
  OA22X1 U32489 ( .IN1(n28938), .IN2(n28512), .IN3(n28955), .IN4(n28511), .Q(
        n28513) );
  NAND4X0 U32490 ( .IN1(n28516), .IN2(n28515), .IN3(n28514), .IN4(n28513), 
        .QN(s0_data_o[31]) );
  OA22X1 U32491 ( .IN1(n28949), .IN2(n28518), .IN3(n28951), .IN4(n28517), .Q(
        n28528) );
  OA22X1 U32492 ( .IN1(n28953), .IN2(n28520), .IN3(n28830), .IN4(n28519), .Q(
        n28527) );
  OA22X1 U32493 ( .IN1(n28844), .IN2(n28522), .IN3(n28847), .IN4(n28521), .Q(
        n28526) );
  OA22X1 U32494 ( .IN1(n28957), .IN2(n28524), .IN3(n28938), .IN4(n28523), .Q(
        n28525) );
  NAND4X0 U32495 ( .IN1(n28528), .IN2(n28527), .IN3(n28526), .IN4(n28525), 
        .QN(s0_sel_o[0]) );
  OA22X1 U32496 ( .IN1(n28947), .IN2(n28530), .IN3(n28830), .IN4(n28529), .Q(
        n28540) );
  OA22X1 U32497 ( .IN1(n28951), .IN2(n28532), .IN3(n28847), .IN4(n28531), .Q(
        n28539) );
  OA22X1 U32498 ( .IN1(n28949), .IN2(n28534), .IN3(n28835), .IN4(n28533), .Q(
        n28538) );
  OA22X1 U32499 ( .IN1(n28957), .IN2(n28536), .IN3(n28945), .IN4(n28535), .Q(
        n28537) );
  NAND4X0 U32500 ( .IN1(n28540), .IN2(n28539), .IN3(n28538), .IN4(n28537), 
        .QN(s0_sel_o[1]) );
  OA22X1 U32501 ( .IN1(n28953), .IN2(n28542), .IN3(n28830), .IN4(n28541), .Q(
        n28552) );
  OA22X1 U32502 ( .IN1(n28949), .IN2(n28544), .IN3(n28844), .IN4(n28543), .Q(
        n28551) );
  OA22X1 U32503 ( .IN1(n28934), .IN2(n28546), .IN3(n28847), .IN4(n28545), .Q(
        n28550) );
  OA22X1 U32504 ( .IN1(n28957), .IN2(n28548), .IN3(n28945), .IN4(n28547), .Q(
        n28549) );
  NAND4X0 U32505 ( .IN1(n28552), .IN2(n28551), .IN3(n28550), .IN4(n28549), 
        .QN(s0_sel_o[2]) );
  OA22X1 U32506 ( .IN1(n28934), .IN2(n28554), .IN3(n28844), .IN4(n28553), .Q(
        n28564) );
  OA22X1 U32507 ( .IN1(n28938), .IN2(n28556), .IN3(n28830), .IN4(n28555), .Q(
        n28563) );
  OA22X1 U32508 ( .IN1(n28862), .IN2(n28558), .IN3(n28918), .IN4(n28557), .Q(
        n28562) );
  OA22X1 U32509 ( .IN1(n28953), .IN2(n28560), .IN3(n28847), .IN4(n28559), .Q(
        n28561) );
  NAND4X0 U32510 ( .IN1(n28564), .IN2(n28563), .IN3(n28562), .IN4(n28561), 
        .QN(s0_sel_o[3]) );
  OA22X1 U32511 ( .IN1(n28957), .IN2(n28566), .IN3(n28847), .IN4(n28565), .Q(
        n28576) );
  OA22X1 U32512 ( .IN1(n28938), .IN2(n28568), .IN3(n28835), .IN4(n28567), .Q(
        n28575) );
  OA22X1 U32513 ( .IN1(n28951), .IN2(n28570), .IN3(n28830), .IN4(n28569), .Q(
        n28574) );
  OA22X1 U32514 ( .IN1(n28862), .IN2(n28572), .IN3(n28844), .IN4(n28571), .Q(
        n28573) );
  NAND4X0 U32515 ( .IN1(n28576), .IN2(n28575), .IN3(n28574), .IN4(n28573), 
        .QN(s0_addr_o[0]) );
  OA22X1 U32516 ( .IN1(n28951), .IN2(n28578), .IN3(n28847), .IN4(n28577), .Q(
        n28588) );
  OA22X1 U32517 ( .IN1(n28949), .IN2(n28580), .IN3(n28938), .IN4(n28579), .Q(
        n28587) );
  OA22X1 U32518 ( .IN1(n28844), .IN2(n28582), .IN3(n28918), .IN4(n28581), .Q(
        n28586) );
  OA22X1 U32519 ( .IN1(n28953), .IN2(n28584), .IN3(n28830), .IN4(n28583), .Q(
        n28585) );
  NAND4X0 U32520 ( .IN1(n28588), .IN2(n28587), .IN3(n28586), .IN4(n28585), 
        .QN(s0_addr_o[1]) );
  OA22X1 U32521 ( .IN1(n28590), .IN2(n28945), .IN3(n28589), .IN4(n28934), .Q(
        n28600) );
  OA22X1 U32522 ( .IN1(n28592), .IN2(n28957), .IN3(n28591), .IN4(n28949), .Q(
        n28599) );
  OA22X1 U32523 ( .IN1(n28594), .IN2(n28947), .IN3(n28593), .IN4(n28953), .Q(
        n28598) );
  OA22X1 U32524 ( .IN1(n28596), .IN2(n28959), .IN3(n28595), .IN4(n28847), .Q(
        n28597) );
  NAND4X0 U32525 ( .IN1(n28600), .IN2(n28599), .IN3(n28598), .IN4(n28597), 
        .QN(s0_addr_o[2]) );
  OA22X1 U32526 ( .IN1(n28602), .IN2(n28953), .IN3(n28601), .IN4(n28949), .Q(
        n28612) );
  OA22X1 U32527 ( .IN1(n28604), .IN2(n28947), .IN3(n28603), .IN4(n28847), .Q(
        n28611) );
  OA22X1 U32528 ( .IN1(n28606), .IN2(n28938), .IN3(n28605), .IN4(n28934), .Q(
        n28610) );
  OA22X1 U32529 ( .IN1(n28608), .IN2(n28959), .IN3(n28607), .IN4(n28957), .Q(
        n28609) );
  NAND4X0 U32530 ( .IN1(n28612), .IN2(n28611), .IN3(n28610), .IN4(n28609), 
        .QN(s0_addr_o[3]) );
  OA22X1 U32531 ( .IN1(n28614), .IN2(n28835), .IN3(n28613), .IN4(n28844), .Q(
        n28624) );
  OA22X1 U32532 ( .IN1(n28616), .IN2(n28951), .IN3(n28615), .IN4(n28945), .Q(
        n28623) );
  OA22X1 U32533 ( .IN1(n28618), .IN2(n28918), .IN3(n28617), .IN4(n28949), .Q(
        n28622) );
  OA22X1 U32534 ( .IN1(n28620), .IN2(n28955), .IN3(n28619), .IN4(n28959), .Q(
        n28621) );
  NAND4X0 U32535 ( .IN1(n28624), .IN2(n28623), .IN3(n28622), .IN4(n28621), 
        .QN(s0_addr_o[4]) );
  OA22X1 U32536 ( .IN1(n28626), .IN2(n28957), .IN3(n28625), .IN4(n28959), .Q(
        n28636) );
  OA22X1 U32537 ( .IN1(n28628), .IN2(n28955), .IN3(n28627), .IN4(n28953), .Q(
        n28635) );
  OA22X1 U32538 ( .IN1(n28630), .IN2(n28934), .IN3(n28629), .IN4(n28949), .Q(
        n28634) );
  OA22X1 U32539 ( .IN1(n28632), .IN2(n28947), .IN3(n28631), .IN4(n28945), .Q(
        n28633) );
  NAND4X0 U32540 ( .IN1(n28636), .IN2(n28635), .IN3(n28634), .IN4(n28633), 
        .QN(s0_addr_o[5]) );
  OA22X1 U32541 ( .IN1(n28938), .IN2(n28638), .IN3(n28953), .IN4(n28637), .Q(
        n28648) );
  OA22X1 U32542 ( .IN1(n28934), .IN2(n28640), .IN3(n28830), .IN4(n28639), .Q(
        n28647) );
  OA22X1 U32543 ( .IN1(n28949), .IN2(n28642), .IN3(n28847), .IN4(n28641), .Q(
        n28646) );
  OA22X1 U32544 ( .IN1(n28947), .IN2(n28644), .IN3(n28918), .IN4(n28643), .Q(
        n28645) );
  NAND4X0 U32545 ( .IN1(n28648), .IN2(n28647), .IN3(n28646), .IN4(n28645), 
        .QN(s0_addr_o[6]) );
  OA22X1 U32546 ( .IN1(n28938), .IN2(n28650), .IN3(n28953), .IN4(n28649), .Q(
        n28660) );
  OA22X1 U32547 ( .IN1(n28934), .IN2(n28652), .IN3(n28847), .IN4(n28651), .Q(
        n28659) );
  OA22X1 U32548 ( .IN1(n28949), .IN2(n28654), .IN3(n28918), .IN4(n28653), .Q(
        n28658) );
  OA22X1 U32549 ( .IN1(n28844), .IN2(n28656), .IN3(n28830), .IN4(n28655), .Q(
        n28657) );
  NAND4X0 U32550 ( .IN1(n28660), .IN2(n28659), .IN3(n28658), .IN4(n28657), 
        .QN(s0_addr_o[7]) );
  OA22X1 U32551 ( .IN1(n28835), .IN2(n28662), .IN3(n28847), .IN4(n28661), .Q(
        n28672) );
  OA22X1 U32552 ( .IN1(n28862), .IN2(n28664), .IN3(n28951), .IN4(n28663), .Q(
        n28671) );
  OA22X1 U32553 ( .IN1(n28947), .IN2(n28666), .IN3(n28918), .IN4(n28665), .Q(
        n28670) );
  OA22X1 U32554 ( .IN1(n28938), .IN2(n28668), .IN3(n28830), .IN4(n28667), .Q(
        n28669) );
  NAND4X0 U32555 ( .IN1(n28672), .IN2(n28671), .IN3(n28670), .IN4(n28669), 
        .QN(s0_addr_o[8]) );
  OA22X1 U32556 ( .IN1(n28844), .IN2(n28674), .IN3(n28938), .IN4(n28673), .Q(
        n28684) );
  OA22X1 U32557 ( .IN1(n28957), .IN2(n28676), .IN3(n28847), .IN4(n28675), .Q(
        n28683) );
  OA22X1 U32558 ( .IN1(n28953), .IN2(n28678), .IN3(n28830), .IN4(n28677), .Q(
        n28682) );
  OA22X1 U32559 ( .IN1(n28862), .IN2(n28680), .IN3(n28951), .IN4(n28679), .Q(
        n28681) );
  NAND4X0 U32560 ( .IN1(n28684), .IN2(n28683), .IN3(n28682), .IN4(n28681), 
        .QN(s0_addr_o[9]) );
  OA22X1 U32561 ( .IN1(n28934), .IN2(n28686), .IN3(n28945), .IN4(n28685), .Q(
        n28696) );
  OA22X1 U32562 ( .IN1(n28947), .IN2(n28688), .IN3(n28957), .IN4(n28687), .Q(
        n28695) );
  OA22X1 U32563 ( .IN1(n28847), .IN2(n28690), .IN3(n28830), .IN4(n28689), .Q(
        n28694) );
  OA22X1 U32564 ( .IN1(n28949), .IN2(n28692), .IN3(n28835), .IN4(n28691), .Q(
        n28693) );
  NAND4X0 U32565 ( .IN1(n28696), .IN2(n28695), .IN3(n28694), .IN4(n28693), 
        .QN(s0_addr_o[10]) );
  OA22X1 U32566 ( .IN1(n28951), .IN2(n28698), .IN3(n28844), .IN4(n28697), .Q(
        n28708) );
  OA22X1 U32567 ( .IN1(n28847), .IN2(n28700), .IN3(n28830), .IN4(n28699), .Q(
        n28707) );
  OA22X1 U32568 ( .IN1(n28949), .IN2(n28702), .IN3(n28938), .IN4(n28701), .Q(
        n28706) );
  OA22X1 U32569 ( .IN1(n28957), .IN2(n28704), .IN3(n28953), .IN4(n28703), .Q(
        n28705) );
  NAND4X0 U32570 ( .IN1(n28708), .IN2(n28707), .IN3(n28706), .IN4(n28705), 
        .QN(s0_addr_o[11]) );
  OA22X1 U32571 ( .IN1(n28934), .IN2(n28710), .IN3(n28938), .IN4(n28709), .Q(
        n28720) );
  OA22X1 U32572 ( .IN1(n28844), .IN2(n28712), .IN3(n28847), .IN4(n28711), .Q(
        n28719) );
  OA22X1 U32573 ( .IN1(n28949), .IN2(n28714), .IN3(n28830), .IN4(n28713), .Q(
        n28718) );
  OA22X1 U32574 ( .IN1(n28918), .IN2(n28716), .IN3(n28953), .IN4(n28715), .Q(
        n28717) );
  NAND4X0 U32575 ( .IN1(n28720), .IN2(n28719), .IN3(n28718), .IN4(n28717), 
        .QN(s0_addr_o[12]) );
  OA22X1 U32576 ( .IN1(n28862), .IN2(n28722), .IN3(n28835), .IN4(n28721), .Q(
        n28732) );
  OA22X1 U32577 ( .IN1(n28957), .IN2(n28724), .IN3(n28945), .IN4(n28723), .Q(
        n28731) );
  OA22X1 U32578 ( .IN1(n28947), .IN2(n28726), .IN3(n28847), .IN4(n28725), .Q(
        n28730) );
  OA22X1 U32579 ( .IN1(n28951), .IN2(n28728), .IN3(n28830), .IN4(n28727), .Q(
        n28729) );
  NAND4X0 U32580 ( .IN1(n28732), .IN2(n28731), .IN3(n28730), .IN4(n28729), 
        .QN(s0_addr_o[13]) );
  OA22X1 U32581 ( .IN1(n28949), .IN2(n28734), .IN3(n28847), .IN4(n28733), .Q(
        n28744) );
  OA22X1 U32582 ( .IN1(n28844), .IN2(n28736), .IN3(n28918), .IN4(n28735), .Q(
        n28743) );
  OA22X1 U32583 ( .IN1(n28934), .IN2(n28738), .IN3(n28835), .IN4(n28737), .Q(
        n28742) );
  OA22X1 U32584 ( .IN1(n28938), .IN2(n28740), .IN3(n28830), .IN4(n28739), .Q(
        n28741) );
  NAND4X0 U32585 ( .IN1(n28744), .IN2(n28743), .IN3(n28742), .IN4(n28741), 
        .QN(s0_addr_o[14]) );
  OA22X1 U32586 ( .IN1(n28862), .IN2(n28746), .IN3(n28830), .IN4(n28745), .Q(
        n28756) );
  OA22X1 U32587 ( .IN1(n28951), .IN2(n28748), .IN3(n28945), .IN4(n28747), .Q(
        n28755) );
  OA22X1 U32588 ( .IN1(n28947), .IN2(n28750), .IN3(n28847), .IN4(n28749), .Q(
        n28754) );
  OA22X1 U32589 ( .IN1(n28957), .IN2(n28752), .IN3(n28953), .IN4(n28751), .Q(
        n28753) );
  NAND4X0 U32590 ( .IN1(n28756), .IN2(n28755), .IN3(n28754), .IN4(n28753), 
        .QN(s0_addr_o[15]) );
  OA22X1 U32591 ( .IN1(n28862), .IN2(n28758), .IN3(n28835), .IN4(n28757), .Q(
        n28768) );
  OA22X1 U32592 ( .IN1(n28947), .IN2(n28760), .IN3(n28938), .IN4(n28759), .Q(
        n28767) );
  OA22X1 U32593 ( .IN1(n28934), .IN2(n28762), .IN3(n28918), .IN4(n28761), .Q(
        n28766) );
  OA22X1 U32594 ( .IN1(n28847), .IN2(n28764), .IN3(n28830), .IN4(n28763), .Q(
        n28765) );
  NAND4X0 U32595 ( .IN1(n28768), .IN2(n28767), .IN3(n28766), .IN4(n28765), 
        .QN(s0_addr_o[16]) );
  OA22X1 U32596 ( .IN1(n28847), .IN2(n28770), .IN3(n28830), .IN4(n28769), .Q(
        n28780) );
  OA22X1 U32597 ( .IN1(n28862), .IN2(n28772), .IN3(n28953), .IN4(n28771), .Q(
        n28779) );
  OA22X1 U32598 ( .IN1(n28844), .IN2(n28774), .IN3(n28918), .IN4(n28773), .Q(
        n28778) );
  OA22X1 U32599 ( .IN1(n28951), .IN2(n28776), .IN3(n28945), .IN4(n28775), .Q(
        n28777) );
  NAND4X0 U32600 ( .IN1(n28780), .IN2(n28779), .IN3(n28778), .IN4(n28777), 
        .QN(s0_addr_o[17]) );
  OA22X1 U32601 ( .IN1(n28918), .IN2(n28782), .IN3(n28830), .IN4(n28781), .Q(
        n28792) );
  OA22X1 U32602 ( .IN1(n28938), .IN2(n28784), .IN3(n28953), .IN4(n28783), .Q(
        n28791) );
  OA22X1 U32603 ( .IN1(n28949), .IN2(n28786), .IN3(n28847), .IN4(n28785), .Q(
        n28790) );
  OA22X1 U32604 ( .IN1(n28951), .IN2(n28788), .IN3(n28844), .IN4(n28787), .Q(
        n28789) );
  NAND4X0 U32605 ( .IN1(n28792), .IN2(n28791), .IN3(n28790), .IN4(n28789), 
        .QN(s0_addr_o[18]) );
  OA22X1 U32606 ( .IN1(n28957), .IN2(n28794), .IN3(n28847), .IN4(n28793), .Q(
        n28804) );
  OA22X1 U32607 ( .IN1(n28949), .IN2(n28796), .IN3(n28835), .IN4(n28795), .Q(
        n28803) );
  OA22X1 U32608 ( .IN1(n28947), .IN2(n28798), .IN3(n28938), .IN4(n28797), .Q(
        n28802) );
  OA22X1 U32609 ( .IN1(n28934), .IN2(n28800), .IN3(n28830), .IN4(n28799), .Q(
        n28801) );
  NAND4X0 U32610 ( .IN1(n28804), .IN2(n28803), .IN3(n28802), .IN4(n28801), 
        .QN(s0_addr_o[19]) );
  OA22X1 U32611 ( .IN1(n28938), .IN2(n28806), .IN3(n28830), .IN4(n28805), .Q(
        n28816) );
  OA22X1 U32612 ( .IN1(n28951), .IN2(n28808), .IN3(n28844), .IN4(n28807), .Q(
        n28815) );
  OA22X1 U32613 ( .IN1(n28918), .IN2(n28810), .IN3(n28847), .IN4(n28809), .Q(
        n28814) );
  OA22X1 U32614 ( .IN1(n28862), .IN2(n28812), .IN3(n28835), .IN4(n28811), .Q(
        n28813) );
  NAND4X0 U32615 ( .IN1(n28816), .IN2(n28815), .IN3(n28814), .IN4(n28813), 
        .QN(s0_addr_o[20]) );
  OA22X1 U32616 ( .IN1(n28955), .IN2(n28818), .IN3(n28830), .IN4(n28817), .Q(
        n28828) );
  OA22X1 U32617 ( .IN1(n28947), .IN2(n28820), .IN3(n28918), .IN4(n28819), .Q(
        n28827) );
  OA22X1 U32618 ( .IN1(n28949), .IN2(n28822), .IN3(n28938), .IN4(n28821), .Q(
        n28826) );
  OA22X1 U32619 ( .IN1(n28951), .IN2(n28824), .IN3(n28953), .IN4(n28823), .Q(
        n28825) );
  NAND4X0 U32620 ( .IN1(n28828), .IN2(n28827), .IN3(n28826), .IN4(n28825), 
        .QN(s0_addr_o[21]) );
  OA22X1 U32621 ( .IN1(n28947), .IN2(n28831), .IN3(n28830), .IN4(n28829), .Q(
        n28842) );
  OA22X1 U32622 ( .IN1(n28862), .IN2(n28833), .IN3(n28951), .IN4(n28832), .Q(
        n28841) );
  OA22X1 U32623 ( .IN1(n28945), .IN2(n28836), .IN3(n28835), .IN4(n28834), .Q(
        n28840) );
  OA22X1 U32624 ( .IN1(n28957), .IN2(n28838), .IN3(n28847), .IN4(n28837), .Q(
        n28839) );
  NAND4X0 U32625 ( .IN1(n28842), .IN2(n28841), .IN3(n28840), .IN4(n28839), 
        .QN(s0_addr_o[22]) );
  OA22X1 U32626 ( .IN1(n28934), .IN2(n28845), .IN3(n28844), .IN4(n28843), .Q(
        n28856) );
  OA22X1 U32627 ( .IN1(n28862), .IN2(n28848), .IN3(n28847), .IN4(n28846), .Q(
        n28855) );
  OA22X1 U32628 ( .IN1(n28957), .IN2(n28850), .IN3(n28953), .IN4(n28849), .Q(
        n28854) );
  OA22X1 U32629 ( .IN1(n28938), .IN2(n28852), .IN3(n28959), .IN4(n28851), .Q(
        n28853) );
  NAND4X0 U32630 ( .IN1(n28856), .IN2(n28855), .IN3(n28854), .IN4(n28853), 
        .QN(s0_addr_o[23]) );
  OA22X1 U32631 ( .IN1(n28858), .IN2(n28947), .IN3(n28857), .IN4(n28918), .Q(
        n28869) );
  OA22X1 U32632 ( .IN1(n28860), .IN2(n28959), .IN3(n28859), .IN4(n28953), .Q(
        n28868) );
  OA22X1 U32633 ( .IN1(n28863), .IN2(n28862), .IN3(n28861), .IN4(n28945), .Q(
        n28867) );
  OA22X1 U32634 ( .IN1(n28865), .IN2(n28955), .IN3(n28864), .IN4(n28951), .Q(
        n28866) );
  NAND4X0 U32635 ( .IN1(n28869), .IN2(n28868), .IN3(n28867), .IN4(n28866), 
        .QN(s0_addr_o[24]) );
  OA22X1 U32636 ( .IN1(n28871), .IN2(n28955), .IN3(n28870), .IN4(n28949), .Q(
        n28881) );
  OA22X1 U32637 ( .IN1(n28873), .IN2(n28947), .IN3(n28872), .IN4(n28945), .Q(
        n28880) );
  OA22X1 U32638 ( .IN1(n28875), .IN2(n28959), .IN3(n28874), .IN4(n28918), .Q(
        n28879) );
  OA22X1 U32639 ( .IN1(n28877), .IN2(n28951), .IN3(n28876), .IN4(n28953), .Q(
        n28878) );
  NAND4X0 U32640 ( .IN1(n28881), .IN2(n28880), .IN3(n28879), .IN4(n28878), 
        .QN(s0_addr_o[25]) );
  OA22X1 U32641 ( .IN1(n28883), .IN2(n28955), .IN3(n28882), .IN4(n28918), .Q(
        n28893) );
  OA22X1 U32642 ( .IN1(n28885), .IN2(n28947), .IN3(n28884), .IN4(n28949), .Q(
        n28892) );
  OA22X1 U32643 ( .IN1(n28887), .IN2(n28934), .IN3(n28886), .IN4(n28938), .Q(
        n28891) );
  OA22X1 U32644 ( .IN1(n28889), .IN2(n28959), .IN3(n28888), .IN4(n28953), .Q(
        n28890) );
  NAND4X0 U32645 ( .IN1(n28893), .IN2(n28892), .IN3(n28891), .IN4(n28890), 
        .QN(s0_addr_o[26]) );
  OA22X1 U32646 ( .IN1(n28895), .IN2(n28951), .IN3(n28894), .IN4(n28949), .Q(
        n28905) );
  OA22X1 U32647 ( .IN1(n28897), .IN2(n28955), .IN3(n28896), .IN4(n28953), .Q(
        n28904) );
  OA22X1 U32648 ( .IN1(n28899), .IN2(n28947), .IN3(n28898), .IN4(n28959), .Q(
        n28903) );
  OA22X1 U32649 ( .IN1(n28901), .IN2(n28918), .IN3(n28900), .IN4(n28945), .Q(
        n28902) );
  NAND4X0 U32650 ( .IN1(n28905), .IN2(n28904), .IN3(n28903), .IN4(n28902), 
        .QN(s0_addr_o[27]) );
  OA22X1 U32651 ( .IN1(n28907), .IN2(n28955), .IN3(n28906), .IN4(n28945), .Q(
        n28917) );
  OA22X1 U32652 ( .IN1(n28909), .IN2(n28947), .IN3(n28908), .IN4(n28918), .Q(
        n28916) );
  OA22X1 U32653 ( .IN1(n28911), .IN2(n28934), .IN3(n28910), .IN4(n28953), .Q(
        n28915) );
  OA22X1 U32654 ( .IN1(n28913), .IN2(n28959), .IN3(n28912), .IN4(n28949), .Q(
        n28914) );
  NAND4X0 U32655 ( .IN1(n28917), .IN2(n28916), .IN3(n28915), .IN4(n28914), 
        .QN(s0_addr_o[28]) );
  OA22X1 U32656 ( .IN1(n28920), .IN2(n28953), .IN3(n28919), .IN4(n28918), .Q(
        n28930) );
  OA22X1 U32657 ( .IN1(n28922), .IN2(n28955), .IN3(n28921), .IN4(n28959), .Q(
        n28929) );
  OA22X1 U32658 ( .IN1(n28924), .IN2(n28951), .IN3(n28923), .IN4(n28938), .Q(
        n28928) );
  OA22X1 U32659 ( .IN1(n28926), .IN2(n28947), .IN3(n28925), .IN4(n28949), .Q(
        n28927) );
  NAND4X0 U32660 ( .IN1(n28930), .IN2(n28929), .IN3(n28928), .IN4(n28927), 
        .QN(s0_addr_o[29]) );
  OA22X1 U32661 ( .IN1(n28932), .IN2(n28947), .IN3(n28931), .IN4(n28949), .Q(
        n28944) );
  OA22X1 U32662 ( .IN1(n28935), .IN2(n28934), .IN3(n28933), .IN4(n28959), .Q(
        n28943) );
  OA22X1 U32663 ( .IN1(n28937), .IN2(n28955), .IN3(n28936), .IN4(n28953), .Q(
        n28942) );
  OA22X1 U32664 ( .IN1(n28940), .IN2(n28957), .IN3(n28939), .IN4(n28938), .Q(
        n28941) );
  NAND4X0 U32665 ( .IN1(n28944), .IN2(n28943), .IN3(n28942), .IN4(n28941), 
        .QN(s0_addr_o[30]) );
  OA22X1 U32666 ( .IN1(n28948), .IN2(n28947), .IN3(n28946), .IN4(n28945), .Q(
        n28964) );
  OA22X1 U32667 ( .IN1(n28952), .IN2(n28951), .IN3(n28950), .IN4(n28949), .Q(
        n28963) );
  OA22X1 U32668 ( .IN1(n28956), .IN2(n28955), .IN3(n28954), .IN4(n28953), .Q(
        n28962) );
  OA22X1 U32669 ( .IN1(n28960), .IN2(n28959), .IN3(n28958), .IN4(n28957), .Q(
        n28961) );
  NAND4X0 U32670 ( .IN1(n28964), .IN2(n28963), .IN3(n28962), .IN4(n28961), 
        .QN(s0_addr_o[31]) );
  NAND3X0 U32671 ( .IN1(m5s0_cyc), .IN2(n28965), .IN3(\s0/m5_cyc_r ), .QN(
        n28972) );
  NAND3X0 U32672 ( .IN1(m6s0_cyc), .IN2(n28966), .IN3(\s0/m6_cyc_r ), .QN(
        n28971) );
  NAND3X0 U32673 ( .IN1(m3s0_cyc), .IN2(n28967), .IN3(\s0/m3_cyc_r ), .QN(
        n28970) );
  NAND3X0 U32674 ( .IN1(m1s0_cyc), .IN2(n28968), .IN3(\s0/m1_cyc_r ), .QN(
        n28969) );
  NAND4X0 U32675 ( .IN1(n28972), .IN2(n28971), .IN3(n28970), .IN4(n28969), 
        .QN(n28982) );
  NAND3X0 U32676 ( .IN1(m4s0_cyc), .IN2(n28973), .IN3(\s0/m4_cyc_r ), .QN(
        n28980) );
  NAND3X0 U32677 ( .IN1(m0s0_cyc), .IN2(n28974), .IN3(\s0/m0_cyc_r ), .QN(
        n28979) );
  NAND3X0 U32678 ( .IN1(m2s0_cyc), .IN2(n28975), .IN3(\s0/m2_cyc_r ), .QN(
        n28978) );
  NAND3X0 U32679 ( .IN1(m7s0_cyc), .IN2(n28976), .IN3(\s0/m7_cyc_r ), .QN(
        n28977) );
  NAND4X0 U32680 ( .IN1(n28980), .IN2(n28979), .IN3(n28978), .IN4(n28977), 
        .QN(n28981) );
  NOR2X0 U32681 ( .IN1(n28982), .IN2(n28981), .QN(n18193) );
  INVX0 U32682 ( .INP(n18193), .ZN(s0_cyc_o) );
  NAND3X0 U32683 ( .IN1(m6s1_cyc), .IN2(n28983), .IN3(\s1/m6_cyc_r ), .QN(
        n28990) );
  NAND3X0 U32684 ( .IN1(m0s1_cyc), .IN2(n28984), .IN3(\s1/m0_cyc_r ), .QN(
        n28989) );
  NAND3X0 U32685 ( .IN1(m2s1_cyc), .IN2(n28985), .IN3(\s1/m2_cyc_r ), .QN(
        n28988) );
  NAND3X0 U32686 ( .IN1(m3s1_cyc), .IN2(n28986), .IN3(\s1/m3_cyc_r ), .QN(
        n28987) );
  NAND4X0 U32687 ( .IN1(n28990), .IN2(n28989), .IN3(n28988), .IN4(n28987), 
        .QN(n29000) );
  NAND3X0 U32688 ( .IN1(m5s1_cyc), .IN2(n28991), .IN3(\s1/m5_cyc_r ), .QN(
        n28998) );
  NAND3X0 U32689 ( .IN1(m4s1_cyc), .IN2(n28992), .IN3(\s1/m4_cyc_r ), .QN(
        n28997) );
  NAND3X0 U32690 ( .IN1(m1s1_cyc), .IN2(n28993), .IN3(\s1/m1_cyc_r ), .QN(
        n28996) );
  NAND3X0 U32691 ( .IN1(m7s1_cyc), .IN2(n28994), .IN3(\s1/m7_cyc_r ), .QN(
        n28995) );
  NAND4X0 U32692 ( .IN1(n28998), .IN2(n28997), .IN3(n28996), .IN4(n28995), 
        .QN(n28999) );
  NOR2X0 U32693 ( .IN1(n29000), .IN2(n28999), .QN(n18192) );
  INVX0 U32694 ( .INP(n18192), .ZN(s1_cyc_o) );
  NAND3X0 U32695 ( .IN1(n29001), .IN2(m6s2_cyc), .IN3(\s2/m6_cyc_r ), .QN(
        n29008) );
  NAND3X0 U32696 ( .IN1(n29002), .IN2(m0s2_cyc), .IN3(\s2/m0_cyc_r ), .QN(
        n29007) );
  NAND3X0 U32697 ( .IN1(n29003), .IN2(m2s2_cyc), .IN3(\s2/m2_cyc_r ), .QN(
        n29006) );
  NAND3X0 U32698 ( .IN1(n29004), .IN2(m7s2_cyc), .IN3(\s2/m7_cyc_r ), .QN(
        n29005) );
  NAND4X0 U32699 ( .IN1(n29008), .IN2(n29007), .IN3(n29006), .IN4(n29005), 
        .QN(n29018) );
  NAND3X0 U32700 ( .IN1(n29009), .IN2(m1s2_cyc), .IN3(\s2/m1_cyc_r ), .QN(
        n29016) );
  NAND3X0 U32701 ( .IN1(n29010), .IN2(m5s2_cyc), .IN3(\s2/m5_cyc_r ), .QN(
        n29015) );
  NAND3X0 U32702 ( .IN1(n29011), .IN2(m3s2_cyc), .IN3(\s2/m3_cyc_r ), .QN(
        n29014) );
  NAND3X0 U32703 ( .IN1(n29012), .IN2(m4s2_cyc), .IN3(\s2/m4_cyc_r ), .QN(
        n29013) );
  NAND4X0 U32704 ( .IN1(n29016), .IN2(n29015), .IN3(n29014), .IN4(n29013), 
        .QN(n29017) );
  NOR2X0 U32705 ( .IN1(n29018), .IN2(n29017), .QN(n18191) );
  INVX0 U32706 ( .INP(n18191), .ZN(s2_cyc_o) );
  NAND3X0 U32707 ( .IN1(m5s3_cyc), .IN2(n29019), .IN3(\s3/m5_cyc_r ), .QN(
        n29026) );
  NAND3X0 U32708 ( .IN1(m7s3_cyc), .IN2(n29020), .IN3(\s3/m7_cyc_r ), .QN(
        n29025) );
  NAND3X0 U32709 ( .IN1(m2s3_cyc), .IN2(n29021), .IN3(\s3/m2_cyc_r ), .QN(
        n29024) );
  NAND3X0 U32710 ( .IN1(m4s3_cyc), .IN2(n29022), .IN3(\s3/m4_cyc_r ), .QN(
        n29023) );
  NAND4X0 U32711 ( .IN1(n29026), .IN2(n29025), .IN3(n29024), .IN4(n29023), 
        .QN(n29036) );
  NAND3X0 U32712 ( .IN1(m1s3_cyc), .IN2(n29027), .IN3(\s3/m1_cyc_r ), .QN(
        n29034) );
  NAND3X0 U32713 ( .IN1(m3s3_cyc), .IN2(n29028), .IN3(\s3/m3_cyc_r ), .QN(
        n29033) );
  NAND3X0 U32714 ( .IN1(m6s3_cyc), .IN2(n29029), .IN3(\s3/m6_cyc_r ), .QN(
        n29032) );
  NAND3X0 U32715 ( .IN1(m0s3_cyc), .IN2(n29030), .IN3(\s3/m0_cyc_r ), .QN(
        n29031) );
  NAND4X0 U32716 ( .IN1(n29034), .IN2(n29033), .IN3(n29032), .IN4(n29031), 
        .QN(n29035) );
  NOR2X0 U32717 ( .IN1(n29036), .IN2(n29035), .QN(n18190) );
  INVX0 U32718 ( .INP(n18190), .ZN(s3_cyc_o) );
  NAND3X0 U32719 ( .IN1(m2s4_cyc), .IN2(n29037), .IN3(\s4/m2_cyc_r ), .QN(
        n29044) );
  NAND3X0 U32720 ( .IN1(m0s4_cyc), .IN2(n29038), .IN3(\s4/m0_cyc_r ), .QN(
        n29043) );
  NAND3X0 U32721 ( .IN1(m6s4_cyc), .IN2(n29039), .IN3(\s4/m6_cyc_r ), .QN(
        n29042) );
  NAND3X0 U32722 ( .IN1(m1s4_cyc), .IN2(n29040), .IN3(\s4/m1_cyc_r ), .QN(
        n29041) );
  NAND4X0 U32723 ( .IN1(n29044), .IN2(n29043), .IN3(n29042), .IN4(n29041), 
        .QN(n29054) );
  NAND3X0 U32724 ( .IN1(m5s4_cyc), .IN2(n29045), .IN3(\s4/m5_cyc_r ), .QN(
        n29052) );
  NAND3X0 U32725 ( .IN1(m3s4_cyc), .IN2(n29046), .IN3(\s4/m3_cyc_r ), .QN(
        n29051) );
  NAND3X0 U32726 ( .IN1(m7s4_cyc), .IN2(n29047), .IN3(\s4/m7_cyc_r ), .QN(
        n29050) );
  NAND3X0 U32727 ( .IN1(m4s4_cyc), .IN2(n29048), .IN3(\s4/m4_cyc_r ), .QN(
        n29049) );
  NAND4X0 U32728 ( .IN1(n29052), .IN2(n29051), .IN3(n29050), .IN4(n29049), 
        .QN(n29053) );
  NOR2X0 U32729 ( .IN1(n29054), .IN2(n29053), .QN(n18189) );
  INVX0 U32730 ( .INP(n18189), .ZN(s4_cyc_o) );
  NAND3X0 U32731 ( .IN1(n29055), .IN2(m2s5_cyc), .IN3(\s5/m2_cyc_r ), .QN(
        n29062) );
  NAND3X0 U32732 ( .IN1(n29056), .IN2(m5s5_cyc), .IN3(\s5/m5_cyc_r ), .QN(
        n29061) );
  NAND3X0 U32733 ( .IN1(n29057), .IN2(m6s5_cyc), .IN3(\s5/m6_cyc_r ), .QN(
        n29060) );
  NAND3X0 U32734 ( .IN1(n29058), .IN2(m1s5_cyc), .IN3(\s5/m1_cyc_r ), .QN(
        n29059) );
  NAND4X0 U32735 ( .IN1(n29062), .IN2(n29061), .IN3(n29060), .IN4(n29059), 
        .QN(n29072) );
  NAND3X0 U32736 ( .IN1(n29063), .IN2(m4s5_cyc), .IN3(\s5/m4_cyc_r ), .QN(
        n29070) );
  NAND3X0 U32737 ( .IN1(n29064), .IN2(m3s5_cyc), .IN3(\s5/m3_cyc_r ), .QN(
        n29069) );
  NAND3X0 U32738 ( .IN1(n29065), .IN2(m7s5_cyc), .IN3(\s5/m7_cyc_r ), .QN(
        n29068) );
  NAND3X0 U32739 ( .IN1(n29066), .IN2(m0s5_cyc), .IN3(\s5/m0_cyc_r ), .QN(
        n29067) );
  NAND4X0 U32740 ( .IN1(n29070), .IN2(n29069), .IN3(n29068), .IN4(n29067), 
        .QN(n29071) );
  NOR2X0 U32741 ( .IN1(n29072), .IN2(n29071), .QN(n18188) );
  INVX0 U32742 ( .INP(n18188), .ZN(s5_cyc_o) );
  NAND3X0 U32743 ( .IN1(m3s6_cyc), .IN2(n29073), .IN3(\s6/m3_cyc_r ), .QN(
        n29080) );
  NAND3X0 U32744 ( .IN1(m6s6_cyc), .IN2(n29074), .IN3(\s6/m6_cyc_r ), .QN(
        n29079) );
  NAND3X0 U32745 ( .IN1(m7s6_cyc), .IN2(n29075), .IN3(\s6/m7_cyc_r ), .QN(
        n29078) );
  NAND3X0 U32746 ( .IN1(m1s6_cyc), .IN2(n29076), .IN3(\s6/m1_cyc_r ), .QN(
        n29077) );
  NAND4X0 U32747 ( .IN1(n29080), .IN2(n29079), .IN3(n29078), .IN4(n29077), 
        .QN(n29090) );
  NAND3X0 U32748 ( .IN1(m0s6_cyc), .IN2(n29081), .IN3(\s6/m0_cyc_r ), .QN(
        n29088) );
  NAND3X0 U32749 ( .IN1(m2s6_cyc), .IN2(n29082), .IN3(\s6/m2_cyc_r ), .QN(
        n29087) );
  NAND3X0 U32750 ( .IN1(m4s6_cyc), .IN2(n29083), .IN3(\s6/m4_cyc_r ), .QN(
        n29086) );
  NAND3X0 U32751 ( .IN1(m5s6_cyc), .IN2(n29084), .IN3(\s6/m5_cyc_r ), .QN(
        n29085) );
  NAND4X0 U32752 ( .IN1(n29088), .IN2(n29087), .IN3(n29086), .IN4(n29085), 
        .QN(n29089) );
  NOR2X0 U32753 ( .IN1(n29090), .IN2(n29089), .QN(n18187) );
  INVX0 U32754 ( .INP(n18187), .ZN(s6_cyc_o) );
  NAND3X0 U32755 ( .IN1(n29091), .IN2(m2s7_cyc), .IN3(\s7/m2_cyc_r ), .QN(
        n29098) );
  NAND3X0 U32756 ( .IN1(n29092), .IN2(m3s7_cyc), .IN3(\s7/m3_cyc_r ), .QN(
        n29097) );
  NAND3X0 U32757 ( .IN1(n29093), .IN2(m1s7_cyc), .IN3(\s7/m1_cyc_r ), .QN(
        n29096) );
  NAND3X0 U32758 ( .IN1(n29094), .IN2(m5s7_cyc), .IN3(\s7/m5_cyc_r ), .QN(
        n29095) );
  NAND4X0 U32759 ( .IN1(n29098), .IN2(n29097), .IN3(n29096), .IN4(n29095), 
        .QN(n29108) );
  NAND3X0 U32760 ( .IN1(n29099), .IN2(m0s7_cyc), .IN3(\s7/m0_cyc_r ), .QN(
        n29106) );
  NAND3X0 U32761 ( .IN1(n29100), .IN2(m6s7_cyc), .IN3(\s7/m6_cyc_r ), .QN(
        n29105) );
  NAND3X0 U32762 ( .IN1(n29101), .IN2(m4s7_cyc), .IN3(\s7/m4_cyc_r ), .QN(
        n29104) );
  NAND3X0 U32763 ( .IN1(n29102), .IN2(m7s7_cyc), .IN3(\s7/m7_cyc_r ), .QN(
        n29103) );
  NAND4X0 U32764 ( .IN1(n29106), .IN2(n29105), .IN3(n29104), .IN4(n29103), 
        .QN(n29107) );
  NOR2X0 U32765 ( .IN1(n29108), .IN2(n29107), .QN(n18186) );
  INVX0 U32766 ( .INP(n18186), .ZN(s7_cyc_o) );
  NAND3X0 U32767 ( .IN1(m6s8_cyc), .IN2(n29109), .IN3(\s8/m6_cyc_r ), .QN(
        n29116) );
  NAND3X0 U32768 ( .IN1(m4s8_cyc), .IN2(n29110), .IN3(\s8/m4_cyc_r ), .QN(
        n29115) );
  NAND3X0 U32769 ( .IN1(m7s8_cyc), .IN2(n29111), .IN3(\s8/m7_cyc_r ), .QN(
        n29114) );
  NAND3X0 U32770 ( .IN1(m2s8_cyc), .IN2(n29112), .IN3(\s8/m2_cyc_r ), .QN(
        n29113) );
  NAND4X0 U32771 ( .IN1(n29116), .IN2(n29115), .IN3(n29114), .IN4(n29113), 
        .QN(n29126) );
  NAND3X0 U32772 ( .IN1(m1s8_cyc), .IN2(n29117), .IN3(\s8/m1_cyc_r ), .QN(
        n29124) );
  NAND3X0 U32773 ( .IN1(m5s8_cyc), .IN2(n29118), .IN3(\s8/m5_cyc_r ), .QN(
        n29123) );
  NAND3X0 U32774 ( .IN1(m3s8_cyc), .IN2(n29119), .IN3(\s8/m3_cyc_r ), .QN(
        n29122) );
  NAND3X0 U32775 ( .IN1(m0s8_cyc), .IN2(n29120), .IN3(\s8/m0_cyc_r ), .QN(
        n29121) );
  NAND4X0 U32776 ( .IN1(n29124), .IN2(n29123), .IN3(n29122), .IN4(n29121), 
        .QN(n29125) );
  NOR2X0 U32777 ( .IN1(n29126), .IN2(n29125), .QN(n18185) );
  INVX0 U32778 ( .INP(n18185), .ZN(s8_cyc_o) );
  NAND3X0 U32779 ( .IN1(n29127), .IN2(m3s9_cyc), .IN3(\s9/m3_cyc_r ), .QN(
        n29134) );
  NAND3X0 U32780 ( .IN1(n29128), .IN2(m4s9_cyc), .IN3(\s9/m4_cyc_r ), .QN(
        n29133) );
  NAND3X0 U32781 ( .IN1(n29129), .IN2(m7s9_cyc), .IN3(\s9/m7_cyc_r ), .QN(
        n29132) );
  NAND3X0 U32782 ( .IN1(n29130), .IN2(m0s9_cyc), .IN3(\s9/m0_cyc_r ), .QN(
        n29131) );
  NAND4X0 U32783 ( .IN1(n29134), .IN2(n29133), .IN3(n29132), .IN4(n29131), 
        .QN(n29144) );
  NAND3X0 U32784 ( .IN1(n29135), .IN2(m2s9_cyc), .IN3(\s9/m2_cyc_r ), .QN(
        n29142) );
  NAND3X0 U32785 ( .IN1(n29136), .IN2(m5s9_cyc), .IN3(\s9/m5_cyc_r ), .QN(
        n29141) );
  NAND3X0 U32786 ( .IN1(n29137), .IN2(m1s9_cyc), .IN3(\s9/m1_cyc_r ), .QN(
        n29140) );
  NAND3X0 U32787 ( .IN1(n29138), .IN2(m6s9_cyc), .IN3(\s9/m6_cyc_r ), .QN(
        n29139) );
  NAND4X0 U32788 ( .IN1(n29142), .IN2(n29141), .IN3(n29140), .IN4(n29139), 
        .QN(n29143) );
  NOR2X0 U32789 ( .IN1(n29144), .IN2(n29143), .QN(n18184) );
  INVX0 U32790 ( .INP(n18184), .ZN(s9_cyc_o) );
  NAND3X0 U32791 ( .IN1(n29145), .IN2(m6s10_cyc), .IN3(\s10/m6_cyc_r ), .QN(
        n29152) );
  NAND3X0 U32792 ( .IN1(n29146), .IN2(m7s10_cyc), .IN3(\s10/m7_cyc_r ), .QN(
        n29151) );
  NAND3X0 U32793 ( .IN1(n29147), .IN2(m3s10_cyc), .IN3(\s10/m3_cyc_r ), .QN(
        n29150) );
  NAND3X0 U32794 ( .IN1(n29148), .IN2(m2s10_cyc), .IN3(\s10/m2_cyc_r ), .QN(
        n29149) );
  NAND4X0 U32795 ( .IN1(n29152), .IN2(n29151), .IN3(n29150), .IN4(n29149), 
        .QN(n29162) );
  NAND3X0 U32796 ( .IN1(n29153), .IN2(m1s10_cyc), .IN3(\s10/m1_cyc_r ), .QN(
        n29160) );
  NAND3X0 U32797 ( .IN1(n29154), .IN2(m4s10_cyc), .IN3(\s10/m4_cyc_r ), .QN(
        n29159) );
  NAND3X0 U32798 ( .IN1(n29155), .IN2(m0s10_cyc), .IN3(\s10/m0_cyc_r ), .QN(
        n29158) );
  NAND3X0 U32799 ( .IN1(n29156), .IN2(m5s10_cyc), .IN3(\s10/m5_cyc_r ), .QN(
        n29157) );
  NAND4X0 U32800 ( .IN1(n29160), .IN2(n29159), .IN3(n29158), .IN4(n29157), 
        .QN(n29161) );
  NOR2X0 U32801 ( .IN1(n29162), .IN2(n29161), .QN(n18183) );
  INVX0 U32802 ( .INP(n18183), .ZN(s10_cyc_o) );
  NAND3X0 U32803 ( .IN1(m1s11_cyc), .IN2(n29163), .IN3(\s11/m1_cyc_r ), .QN(
        n29170) );
  NAND3X0 U32804 ( .IN1(m2s11_cyc), .IN2(n29164), .IN3(\s11/m2_cyc_r ), .QN(
        n29169) );
  NAND3X0 U32805 ( .IN1(m0s11_cyc), .IN2(n29165), .IN3(\s11/m0_cyc_r ), .QN(
        n29168) );
  NAND3X0 U32806 ( .IN1(m3s11_cyc), .IN2(n29166), .IN3(\s11/m3_cyc_r ), .QN(
        n29167) );
  NAND4X0 U32807 ( .IN1(n29170), .IN2(n29169), .IN3(n29168), .IN4(n29167), 
        .QN(n29180) );
  NAND3X0 U32808 ( .IN1(m6s11_cyc), .IN2(n29171), .IN3(\s11/m6_cyc_r ), .QN(
        n29178) );
  NAND3X0 U32809 ( .IN1(m4s11_cyc), .IN2(n29172), .IN3(\s11/m4_cyc_r ), .QN(
        n29177) );
  NAND3X0 U32810 ( .IN1(m5s11_cyc), .IN2(n29173), .IN3(\s11/m5_cyc_r ), .QN(
        n29176) );
  NAND3X0 U32811 ( .IN1(m7s11_cyc), .IN2(n29174), .IN3(\s11/m7_cyc_r ), .QN(
        n29175) );
  NAND4X0 U32812 ( .IN1(n29178), .IN2(n29177), .IN3(n29176), .IN4(n29175), 
        .QN(n29179) );
  NOR2X0 U32813 ( .IN1(n29180), .IN2(n29179), .QN(n18182) );
  INVX0 U32814 ( .INP(n18182), .ZN(s11_cyc_o) );
  NAND3X0 U32815 ( .IN1(n29181), .IN2(m1s12_cyc), .IN3(\s12/m1_cyc_r ), .QN(
        n29188) );
  NAND3X0 U32816 ( .IN1(n29182), .IN2(m4s12_cyc), .IN3(\s12/m4_cyc_r ), .QN(
        n29187) );
  NAND3X0 U32817 ( .IN1(n29183), .IN2(m6s12_cyc), .IN3(\s12/m6_cyc_r ), .QN(
        n29186) );
  NAND3X0 U32818 ( .IN1(n29184), .IN2(m3s12_cyc), .IN3(\s12/m3_cyc_r ), .QN(
        n29185) );
  NAND4X0 U32819 ( .IN1(n29188), .IN2(n29187), .IN3(n29186), .IN4(n29185), 
        .QN(n29198) );
  NAND3X0 U32820 ( .IN1(n29189), .IN2(m5s12_cyc), .IN3(\s12/m5_cyc_r ), .QN(
        n29196) );
  NAND3X0 U32821 ( .IN1(n29190), .IN2(m7s12_cyc), .IN3(\s12/m7_cyc_r ), .QN(
        n29195) );
  NAND3X0 U32822 ( .IN1(n29191), .IN2(m0s12_cyc), .IN3(\s12/m0_cyc_r ), .QN(
        n29194) );
  NAND3X0 U32823 ( .IN1(n29192), .IN2(m2s12_cyc), .IN3(\s12/m2_cyc_r ), .QN(
        n29193) );
  NAND4X0 U32824 ( .IN1(n29196), .IN2(n29195), .IN3(n29194), .IN4(n29193), 
        .QN(n29197) );
  NOR2X0 U32825 ( .IN1(n29198), .IN2(n29197), .QN(n18181) );
  INVX0 U32826 ( .INP(n18181), .ZN(s12_cyc_o) );
  NAND3X0 U32827 ( .IN1(n29199), .IN2(m5s13_cyc), .IN3(\s13/m5_cyc_r ), .QN(
        n29206) );
  NAND3X0 U32828 ( .IN1(n29200), .IN2(m1s13_cyc), .IN3(\s13/m1_cyc_r ), .QN(
        n29205) );
  NAND3X0 U32829 ( .IN1(n29201), .IN2(m7s13_cyc), .IN3(\s13/m7_cyc_r ), .QN(
        n29204) );
  NAND3X0 U32830 ( .IN1(n29202), .IN2(m0s13_cyc), .IN3(\s13/m0_cyc_r ), .QN(
        n29203) );
  NAND4X0 U32831 ( .IN1(n29206), .IN2(n29205), .IN3(n29204), .IN4(n29203), 
        .QN(n29216) );
  NAND3X0 U32832 ( .IN1(n29207), .IN2(m2s13_cyc), .IN3(\s13/m2_cyc_r ), .QN(
        n29214) );
  NAND3X0 U32833 ( .IN1(n29208), .IN2(m6s13_cyc), .IN3(\s13/m6_cyc_r ), .QN(
        n29213) );
  NAND3X0 U32834 ( .IN1(n29209), .IN2(m4s13_cyc), .IN3(\s13/m4_cyc_r ), .QN(
        n29212) );
  NAND3X0 U32835 ( .IN1(n29210), .IN2(m3s13_cyc), .IN3(\s13/m3_cyc_r ), .QN(
        n29211) );
  NAND4X0 U32836 ( .IN1(n29214), .IN2(n29213), .IN3(n29212), .IN4(n29211), 
        .QN(n29215) );
  NOR2X0 U32837 ( .IN1(n29216), .IN2(n29215), .QN(n18180) );
  INVX0 U32838 ( .INP(n18180), .ZN(s13_cyc_o) );
  NAND3X0 U32839 ( .IN1(n29217), .IN2(m2s14_cyc), .IN3(\s14/m2_cyc_r ), .QN(
        n29224) );
  NAND3X0 U32840 ( .IN1(n29218), .IN2(m0s14_cyc), .IN3(\s14/m0_cyc_r ), .QN(
        n29223) );
  NAND3X0 U32841 ( .IN1(n29219), .IN2(m4s14_cyc), .IN3(\s14/m4_cyc_r ), .QN(
        n29222) );
  NAND3X0 U32842 ( .IN1(n29220), .IN2(m6s14_cyc), .IN3(\s14/m6_cyc_r ), .QN(
        n29221) );
  NAND4X0 U32843 ( .IN1(n29224), .IN2(n29223), .IN3(n29222), .IN4(n29221), 
        .QN(n29234) );
  NAND3X0 U32844 ( .IN1(n29225), .IN2(m3s14_cyc), .IN3(\s14/m3_cyc_r ), .QN(
        n29232) );
  NAND3X0 U32845 ( .IN1(n29226), .IN2(m5s14_cyc), .IN3(\s14/m5_cyc_r ), .QN(
        n29231) );
  NAND3X0 U32846 ( .IN1(n29227), .IN2(m1s14_cyc), .IN3(\s14/m1_cyc_r ), .QN(
        n29230) );
  NAND3X0 U32847 ( .IN1(n29228), .IN2(m7s14_cyc), .IN3(\s14/m7_cyc_r ), .QN(
        n29229) );
  NAND4X0 U32848 ( .IN1(n29232), .IN2(n29231), .IN3(n29230), .IN4(n29229), 
        .QN(n29233) );
  NOR2X0 U32849 ( .IN1(n29234), .IN2(n29233), .QN(n18179) );
  INVX0 U32850 ( .INP(n18179), .ZN(s14_cyc_o) );
  AND2X1 U32851 ( .IN1(m0_cyc_i), .IN2(n29235), .Q(n29253) );
  AND2X1 U32852 ( .IN1(m0_stb_i), .IN2(m0_cyc_i), .Q(n29251) );
  AO22X1 U32853 ( .IN1(m0s15_cyc), .IN2(n29253), .IN3(n29236), .IN4(n29251), 
        .Q(n18177) );
  AO22X1 U32854 ( .IN1(n29237), .IN2(n29251), .IN3(m0s14_cyc), .IN4(n29253), 
        .Q(n18176) );
  AO22X1 U32855 ( .IN1(n29238), .IN2(n29251), .IN3(m0s13_cyc), .IN4(n29253), 
        .Q(n18175) );
  AO22X1 U32856 ( .IN1(n29239), .IN2(n29251), .IN3(m0s12_cyc), .IN4(n29253), 
        .Q(n18174) );
  AO22X1 U32857 ( .IN1(m0s11_cyc), .IN2(n29253), .IN3(n29240), .IN4(n29251), 
        .Q(n18173) );
  AO22X1 U32858 ( .IN1(n29241), .IN2(n29251), .IN3(m0s10_cyc), .IN4(n29253), 
        .Q(n18172) );
  AO22X1 U32859 ( .IN1(n29242), .IN2(n29251), .IN3(m0s9_cyc), .IN4(n29253), 
        .Q(n18171) );
  AO22X1 U32860 ( .IN1(m0s8_cyc), .IN2(n29253), .IN3(n29243), .IN4(n29251), 
        .Q(n18170) );
  AO22X1 U32861 ( .IN1(n29244), .IN2(n29251), .IN3(m0s7_cyc), .IN4(n29253), 
        .Q(n18169) );
  AO22X1 U32862 ( .IN1(m0s6_cyc), .IN2(n29253), .IN3(n29245), .IN4(n29251), 
        .Q(n18168) );
  AO22X1 U32863 ( .IN1(n29246), .IN2(n29251), .IN3(m0s5_cyc), .IN4(n29253), 
        .Q(n18167) );
  AO22X1 U32864 ( .IN1(m0s4_cyc), .IN2(n29253), .IN3(n29247), .IN4(n29251), 
        .Q(n18166) );
  AO22X1 U32865 ( .IN1(m0s3_cyc), .IN2(n29253), .IN3(n29248), .IN4(n29251), 
        .Q(n18165) );
  AO22X1 U32866 ( .IN1(n29249), .IN2(n29251), .IN3(m0s2_cyc), .IN4(n29253), 
        .Q(n18164) );
  AO22X1 U32867 ( .IN1(m0s1_cyc), .IN2(n29253), .IN3(n29250), .IN4(n29251), 
        .Q(n18163) );
  AO22X1 U32868 ( .IN1(m0s0_cyc), .IN2(n29253), .IN3(n29252), .IN4(n29251), 
        .Q(n18162) );
  AND2X1 U32869 ( .IN1(m1_cyc_i), .IN2(n29254), .Q(n29272) );
  AND2X1 U32870 ( .IN1(m1_stb_i), .IN2(m1_cyc_i), .Q(n29270) );
  AO22X1 U32871 ( .IN1(m1s15_cyc), .IN2(n29272), .IN3(n29255), .IN4(n29270), 
        .Q(n18161) );
  AO22X1 U32872 ( .IN1(n29256), .IN2(n29270), .IN3(m1s14_cyc), .IN4(n29272), 
        .Q(n18160) );
  AO22X1 U32873 ( .IN1(n29257), .IN2(n29270), .IN3(m1s13_cyc), .IN4(n29272), 
        .Q(n18159) );
  AO22X1 U32874 ( .IN1(n29258), .IN2(n29270), .IN3(m1s12_cyc), .IN4(n29272), 
        .Q(n18158) );
  AO22X1 U32875 ( .IN1(m1s11_cyc), .IN2(n29272), .IN3(n29259), .IN4(n29270), 
        .Q(n18157) );
  AO22X1 U32876 ( .IN1(n29260), .IN2(n29270), .IN3(m1s10_cyc), .IN4(n29272), 
        .Q(n18156) );
  AO22X1 U32877 ( .IN1(n29261), .IN2(n29270), .IN3(m1s9_cyc), .IN4(n29272), 
        .Q(n18155) );
  AO22X1 U32878 ( .IN1(m1s8_cyc), .IN2(n29272), .IN3(n29262), .IN4(n29270), 
        .Q(n18154) );
  AO22X1 U32879 ( .IN1(n29263), .IN2(n29270), .IN3(m1s7_cyc), .IN4(n29272), 
        .Q(n18153) );
  AO22X1 U32880 ( .IN1(m1s6_cyc), .IN2(n29272), .IN3(n29264), .IN4(n29270), 
        .Q(n18152) );
  AO22X1 U32881 ( .IN1(n29265), .IN2(n29270), .IN3(m1s5_cyc), .IN4(n29272), 
        .Q(n18151) );
  AO22X1 U32882 ( .IN1(m1s4_cyc), .IN2(n29272), .IN3(n29266), .IN4(n29270), 
        .Q(n18150) );
  AO22X1 U32883 ( .IN1(m1s3_cyc), .IN2(n29272), .IN3(n29267), .IN4(n29270), 
        .Q(n18149) );
  AO22X1 U32884 ( .IN1(n29268), .IN2(n29270), .IN3(m1s2_cyc), .IN4(n29272), 
        .Q(n18148) );
  AO22X1 U32885 ( .IN1(m1s1_cyc), .IN2(n29272), .IN3(n29269), .IN4(n29270), 
        .Q(n18147) );
  AO22X1 U32886 ( .IN1(m1s0_cyc), .IN2(n29272), .IN3(n29271), .IN4(n29270), 
        .Q(n18146) );
  AND2X1 U32887 ( .IN1(m2_cyc_i), .IN2(n29273), .Q(n29291) );
  AND2X1 U32888 ( .IN1(m2_stb_i), .IN2(m2_cyc_i), .Q(n29289) );
  AO22X1 U32889 ( .IN1(m2s15_cyc), .IN2(n29291), .IN3(n29274), .IN4(n29289), 
        .Q(n18145) );
  AO22X1 U32890 ( .IN1(n29275), .IN2(n29289), .IN3(m2s14_cyc), .IN4(n29291), 
        .Q(n18144) );
  AO22X1 U32891 ( .IN1(n29276), .IN2(n29289), .IN3(m2s13_cyc), .IN4(n29291), 
        .Q(n18143) );
  AO22X1 U32892 ( .IN1(n29277), .IN2(n29289), .IN3(m2s12_cyc), .IN4(n29291), 
        .Q(n18142) );
  AO22X1 U32893 ( .IN1(m2s11_cyc), .IN2(n29291), .IN3(n29278), .IN4(n29289), 
        .Q(n18141) );
  AO22X1 U32894 ( .IN1(n29279), .IN2(n29289), .IN3(m2s10_cyc), .IN4(n29291), 
        .Q(n18140) );
  AO22X1 U32895 ( .IN1(n29280), .IN2(n29289), .IN3(m2s9_cyc), .IN4(n29291), 
        .Q(n18139) );
  AO22X1 U32896 ( .IN1(m2s8_cyc), .IN2(n29291), .IN3(n29281), .IN4(n29289), 
        .Q(n18138) );
  AO22X1 U32897 ( .IN1(n29282), .IN2(n29289), .IN3(m2s7_cyc), .IN4(n29291), 
        .Q(n18137) );
  AO22X1 U32898 ( .IN1(m2s6_cyc), .IN2(n29291), .IN3(n29283), .IN4(n29289), 
        .Q(n18136) );
  AO22X1 U32899 ( .IN1(n29284), .IN2(n29289), .IN3(m2s5_cyc), .IN4(n29291), 
        .Q(n18135) );
  AO22X1 U32900 ( .IN1(m2s4_cyc), .IN2(n29291), .IN3(n29285), .IN4(n29289), 
        .Q(n18134) );
  AO22X1 U32901 ( .IN1(m2s3_cyc), .IN2(n29291), .IN3(n29286), .IN4(n29289), 
        .Q(n18133) );
  AO22X1 U32902 ( .IN1(n29287), .IN2(n29289), .IN3(m2s2_cyc), .IN4(n29291), 
        .Q(n18132) );
  AO22X1 U32903 ( .IN1(m2s1_cyc), .IN2(n29291), .IN3(n29288), .IN4(n29289), 
        .Q(n18131) );
  AO22X1 U32904 ( .IN1(m2s0_cyc), .IN2(n29291), .IN3(n29290), .IN4(n29289), 
        .Q(n18130) );
  AND2X1 U32905 ( .IN1(m3_cyc_i), .IN2(n29292), .Q(n29310) );
  AND2X1 U32906 ( .IN1(m3_stb_i), .IN2(m3_cyc_i), .Q(n29308) );
  AO22X1 U32907 ( .IN1(m3s15_cyc), .IN2(n29310), .IN3(n29293), .IN4(n29308), 
        .Q(n18129) );
  AO22X1 U32908 ( .IN1(n29294), .IN2(n29308), .IN3(m3s14_cyc), .IN4(n29310), 
        .Q(n18128) );
  AO22X1 U32909 ( .IN1(n29295), .IN2(n29308), .IN3(m3s13_cyc), .IN4(n29310), 
        .Q(n18127) );
  AO22X1 U32910 ( .IN1(n29296), .IN2(n29308), .IN3(m3s12_cyc), .IN4(n29310), 
        .Q(n18126) );
  AO22X1 U32911 ( .IN1(m3s11_cyc), .IN2(n29310), .IN3(n29297), .IN4(n29308), 
        .Q(n18125) );
  AO22X1 U32912 ( .IN1(n29298), .IN2(n29308), .IN3(m3s10_cyc), .IN4(n29310), 
        .Q(n18124) );
  AO22X1 U32913 ( .IN1(n29299), .IN2(n29308), .IN3(m3s9_cyc), .IN4(n29310), 
        .Q(n18123) );
  AO22X1 U32914 ( .IN1(m3s8_cyc), .IN2(n29310), .IN3(n29300), .IN4(n29308), 
        .Q(n18122) );
  AO22X1 U32915 ( .IN1(n29301), .IN2(n29308), .IN3(m3s7_cyc), .IN4(n29310), 
        .Q(n18121) );
  AO22X1 U32916 ( .IN1(m3s6_cyc), .IN2(n29310), .IN3(n29302), .IN4(n29308), 
        .Q(n18120) );
  AO22X1 U32917 ( .IN1(n29303), .IN2(n29308), .IN3(m3s5_cyc), .IN4(n29310), 
        .Q(n18119) );
  AO22X1 U32918 ( .IN1(m3s4_cyc), .IN2(n29310), .IN3(n29304), .IN4(n29308), 
        .Q(n18118) );
  AO22X1 U32919 ( .IN1(m3s3_cyc), .IN2(n29310), .IN3(n29305), .IN4(n29308), 
        .Q(n18117) );
  AO22X1 U32920 ( .IN1(n29306), .IN2(n29308), .IN3(m3s2_cyc), .IN4(n29310), 
        .Q(n18116) );
  AO22X1 U32921 ( .IN1(m3s1_cyc), .IN2(n29310), .IN3(n29307), .IN4(n29308), 
        .Q(n18115) );
  AO22X1 U32922 ( .IN1(m3s0_cyc), .IN2(n29310), .IN3(n29309), .IN4(n29308), 
        .Q(n18114) );
  AND2X1 U32923 ( .IN1(m4_cyc_i), .IN2(n29311), .Q(n29329) );
  AND2X1 U32924 ( .IN1(m4_stb_i), .IN2(m4_cyc_i), .Q(n29327) );
  AO22X1 U32925 ( .IN1(m4s15_cyc), .IN2(n29329), .IN3(n29312), .IN4(n29327), 
        .Q(n18113) );
  AO22X1 U32926 ( .IN1(n29313), .IN2(n29327), .IN3(m4s14_cyc), .IN4(n29329), 
        .Q(n18112) );
  AO22X1 U32927 ( .IN1(n29314), .IN2(n29327), .IN3(m4s13_cyc), .IN4(n29329), 
        .Q(n18111) );
  AO22X1 U32928 ( .IN1(n29315), .IN2(n29327), .IN3(m4s12_cyc), .IN4(n29329), 
        .Q(n18110) );
  AO22X1 U32929 ( .IN1(m4s11_cyc), .IN2(n29329), .IN3(n29316), .IN4(n29327), 
        .Q(n18109) );
  AO22X1 U32930 ( .IN1(n29317), .IN2(n29327), .IN3(m4s10_cyc), .IN4(n29329), 
        .Q(n18108) );
  AO22X1 U32931 ( .IN1(n29318), .IN2(n29327), .IN3(m4s9_cyc), .IN4(n29329), 
        .Q(n18107) );
  AO22X1 U32932 ( .IN1(m4s8_cyc), .IN2(n29329), .IN3(n29319), .IN4(n29327), 
        .Q(n18106) );
  AO22X1 U32933 ( .IN1(n29320), .IN2(n29327), .IN3(m4s7_cyc), .IN4(n29329), 
        .Q(n18105) );
  AO22X1 U32934 ( .IN1(m4s6_cyc), .IN2(n29329), .IN3(n29321), .IN4(n29327), 
        .Q(n18104) );
  AO22X1 U32935 ( .IN1(n29322), .IN2(n29327), .IN3(m4s5_cyc), .IN4(n29329), 
        .Q(n18103) );
  AO22X1 U32936 ( .IN1(m4s4_cyc), .IN2(n29329), .IN3(n29323), .IN4(n29327), 
        .Q(n18102) );
  AO22X1 U32937 ( .IN1(m4s3_cyc), .IN2(n29329), .IN3(n29324), .IN4(n29327), 
        .Q(n18101) );
  AO22X1 U32938 ( .IN1(n29325), .IN2(n29327), .IN3(m4s2_cyc), .IN4(n29329), 
        .Q(n18100) );
  AO22X1 U32939 ( .IN1(m4s1_cyc), .IN2(n29329), .IN3(n29326), .IN4(n29327), 
        .Q(n18099) );
  AO22X1 U32940 ( .IN1(m4s0_cyc), .IN2(n29329), .IN3(n29328), .IN4(n29327), 
        .Q(n18098) );
  AND2X1 U32941 ( .IN1(m5_cyc_i), .IN2(n29330), .Q(n29348) );
  AND2X1 U32942 ( .IN1(m5_stb_i), .IN2(m5_cyc_i), .Q(n29346) );
  AO22X1 U32943 ( .IN1(m5s15_cyc), .IN2(n29348), .IN3(n29331), .IN4(n29346), 
        .Q(n18097) );
  AO22X1 U32944 ( .IN1(n29332), .IN2(n29346), .IN3(m5s14_cyc), .IN4(n29348), 
        .Q(n18096) );
  AO22X1 U32945 ( .IN1(n29333), .IN2(n29346), .IN3(m5s13_cyc), .IN4(n29348), 
        .Q(n18095) );
  AO22X1 U32946 ( .IN1(n29334), .IN2(n29346), .IN3(m5s12_cyc), .IN4(n29348), 
        .Q(n18094) );
  AO22X1 U32947 ( .IN1(m5s11_cyc), .IN2(n29348), .IN3(n29335), .IN4(n29346), 
        .Q(n18093) );
  AO22X1 U32948 ( .IN1(n29336), .IN2(n29346), .IN3(m5s10_cyc), .IN4(n29348), 
        .Q(n18092) );
  AO22X1 U32949 ( .IN1(n29337), .IN2(n29346), .IN3(m5s9_cyc), .IN4(n29348), 
        .Q(n18091) );
  AO22X1 U32950 ( .IN1(m5s8_cyc), .IN2(n29348), .IN3(n29338), .IN4(n29346), 
        .Q(n18090) );
  AO22X1 U32951 ( .IN1(n29339), .IN2(n29346), .IN3(m5s7_cyc), .IN4(n29348), 
        .Q(n18089) );
  AO22X1 U32952 ( .IN1(m5s6_cyc), .IN2(n29348), .IN3(n29340), .IN4(n29346), 
        .Q(n18088) );
  AO22X1 U32953 ( .IN1(n29341), .IN2(n29346), .IN3(m5s5_cyc), .IN4(n29348), 
        .Q(n18087) );
  AO22X1 U32954 ( .IN1(m5s4_cyc), .IN2(n29348), .IN3(n29342), .IN4(n29346), 
        .Q(n18086) );
  AO22X1 U32955 ( .IN1(m5s3_cyc), .IN2(n29348), .IN3(n29343), .IN4(n29346), 
        .Q(n18085) );
  AO22X1 U32956 ( .IN1(n29344), .IN2(n29346), .IN3(m5s2_cyc), .IN4(n29348), 
        .Q(n18084) );
  AO22X1 U32957 ( .IN1(m5s1_cyc), .IN2(n29348), .IN3(n29345), .IN4(n29346), 
        .Q(n18083) );
  AO22X1 U32958 ( .IN1(m5s0_cyc), .IN2(n29348), .IN3(n29347), .IN4(n29346), 
        .Q(n18082) );
  AND2X1 U32959 ( .IN1(m6_cyc_i), .IN2(n29349), .Q(n29367) );
  AND2X1 U32960 ( .IN1(m6_stb_i), .IN2(m6_cyc_i), .Q(n29365) );
  AO22X1 U32961 ( .IN1(m6s15_cyc), .IN2(n29367), .IN3(n29350), .IN4(n29365), 
        .Q(n18081) );
  AO22X1 U32962 ( .IN1(n29351), .IN2(n29365), .IN3(m6s14_cyc), .IN4(n29367), 
        .Q(n18080) );
  AO22X1 U32963 ( .IN1(n29352), .IN2(n29365), .IN3(m6s13_cyc), .IN4(n29367), 
        .Q(n18079) );
  AO22X1 U32964 ( .IN1(n29353), .IN2(n29365), .IN3(m6s12_cyc), .IN4(n29367), 
        .Q(n18078) );
  AO22X1 U32965 ( .IN1(m6s11_cyc), .IN2(n29367), .IN3(n29354), .IN4(n29365), 
        .Q(n18077) );
  AO22X1 U32966 ( .IN1(n29355), .IN2(n29365), .IN3(m6s10_cyc), .IN4(n29367), 
        .Q(n18076) );
  AO22X1 U32967 ( .IN1(n29356), .IN2(n29365), .IN3(m6s9_cyc), .IN4(n29367), 
        .Q(n18075) );
  AO22X1 U32968 ( .IN1(m6s8_cyc), .IN2(n29367), .IN3(n29357), .IN4(n29365), 
        .Q(n18074) );
  AO22X1 U32969 ( .IN1(n29358), .IN2(n29365), .IN3(m6s7_cyc), .IN4(n29367), 
        .Q(n18073) );
  AO22X1 U32970 ( .IN1(m6s6_cyc), .IN2(n29367), .IN3(n29359), .IN4(n29365), 
        .Q(n18072) );
  AO22X1 U32971 ( .IN1(n29360), .IN2(n29365), .IN3(m6s5_cyc), .IN4(n29367), 
        .Q(n18071) );
  AO22X1 U32972 ( .IN1(m6s4_cyc), .IN2(n29367), .IN3(n29361), .IN4(n29365), 
        .Q(n18070) );
  AO22X1 U32973 ( .IN1(m6s3_cyc), .IN2(n29367), .IN3(n29362), .IN4(n29365), 
        .Q(n18069) );
  AO22X1 U32974 ( .IN1(n29363), .IN2(n29365), .IN3(m6s2_cyc), .IN4(n29367), 
        .Q(n18068) );
  AO22X1 U32975 ( .IN1(m6s1_cyc), .IN2(n29367), .IN3(n29364), .IN4(n29365), 
        .Q(n18067) );
  AO22X1 U32976 ( .IN1(m6s0_cyc), .IN2(n29367), .IN3(n29366), .IN4(n29365), 
        .Q(n18066) );
  AND2X1 U32977 ( .IN1(m7_cyc_i), .IN2(n29368), .Q(n29386) );
  AND2X1 U32978 ( .IN1(m7_stb_i), .IN2(m7_cyc_i), .Q(n29384) );
  AO22X1 U32979 ( .IN1(m7s15_cyc), .IN2(n29386), .IN3(n29369), .IN4(n29384), 
        .Q(n18065) );
  AO22X1 U32980 ( .IN1(n29370), .IN2(n29384), .IN3(m7s14_cyc), .IN4(n29386), 
        .Q(n18064) );
  AO22X1 U32981 ( .IN1(n29371), .IN2(n29384), .IN3(m7s13_cyc), .IN4(n29386), 
        .Q(n18063) );
  AO22X1 U32982 ( .IN1(n29372), .IN2(n29384), .IN3(m7s12_cyc), .IN4(n29386), 
        .Q(n18062) );
  AO22X1 U32983 ( .IN1(m7s11_cyc), .IN2(n29386), .IN3(n29373), .IN4(n29384), 
        .Q(n18061) );
  AO22X1 U32984 ( .IN1(n29374), .IN2(n29384), .IN3(m7s10_cyc), .IN4(n29386), 
        .Q(n18060) );
  AO22X1 U32985 ( .IN1(n29375), .IN2(n29384), .IN3(m7s9_cyc), .IN4(n29386), 
        .Q(n18059) );
  AO22X1 U32986 ( .IN1(m7s8_cyc), .IN2(n29386), .IN3(n29376), .IN4(n29384), 
        .Q(n18058) );
  AO22X1 U32987 ( .IN1(n29377), .IN2(n29384), .IN3(m7s7_cyc), .IN4(n29386), 
        .Q(n18057) );
  AO22X1 U32988 ( .IN1(m7s6_cyc), .IN2(n29386), .IN3(n29378), .IN4(n29384), 
        .Q(n18056) );
  AO22X1 U32989 ( .IN1(n29379), .IN2(n29384), .IN3(m7s5_cyc), .IN4(n29386), 
        .Q(n18055) );
  AO22X1 U32990 ( .IN1(m7s4_cyc), .IN2(n29386), .IN3(n29380), .IN4(n29384), 
        .Q(n18054) );
  AO22X1 U32991 ( .IN1(m7s3_cyc), .IN2(n29386), .IN3(n29381), .IN4(n29384), 
        .Q(n18053) );
  AO22X1 U32992 ( .IN1(n29382), .IN2(n29384), .IN3(m7s2_cyc), .IN4(n29386), 
        .Q(n18052) );
  AO22X1 U32993 ( .IN1(m7s1_cyc), .IN2(n29386), .IN3(n29383), .IN4(n29384), 
        .Q(n18051) );
  AO22X1 U32994 ( .IN1(m7s0_cyc), .IN2(n29386), .IN3(n29385), .IN4(n29384), 
        .Q(n18050) );
  NOR2X0 U32995 ( .IN1(n29387), .IN2(n34379), .QN(n29388) );
  MUX21X1 U32996 ( .IN1(n34623), .IN2(s15_data_o[0]), .S(n29388), .Q(n18049)
         );
  MUX21X1 U32997 ( .IN1(n34572), .IN2(s15_data_o[1]), .S(n29388), .Q(n18048)
         );
  MUX21X1 U32998 ( .IN1(n34624), .IN2(s15_data_o[2]), .S(n29388), .Q(n18047)
         );
  MUX21X1 U32999 ( .IN1(n34573), .IN2(s15_data_o[3]), .S(n29388), .Q(n18046)
         );
  MUX21X1 U33000 ( .IN1(n34612), .IN2(s15_data_o[4]), .S(n29388), .Q(n18045)
         );
  MUX21X1 U33001 ( .IN1(n34574), .IN2(s15_data_o[5]), .S(n29388), .Q(n18044)
         );
  MUX21X1 U33002 ( .IN1(n34613), .IN2(s15_data_o[6]), .S(n29388), .Q(n18043)
         );
  MUX21X1 U33003 ( .IN1(n34561), .IN2(s15_data_o[7]), .S(n29388), .Q(n18042)
         );
  MUX21X1 U33004 ( .IN1(n34304), .IN2(s15_data_o[8]), .S(n29388), .Q(n18041)
         );
  MUX21X1 U33005 ( .IN1(n34519), .IN2(s15_data_o[9]), .S(n29388), .Q(n18040)
         );
  MUX21X1 U33006 ( .IN1(n34305), .IN2(s15_data_o[10]), .S(n29388), .Q(n18039)
         );
  MUX21X1 U33007 ( .IN1(n34520), .IN2(s15_data_o[11]), .S(n29388), .Q(n18038)
         );
  MUX21X1 U33008 ( .IN1(n34614), .IN2(s15_data_o[12]), .S(n29388), .Q(n18037)
         );
  MUX21X1 U33009 ( .IN1(n34575), .IN2(s15_data_o[13]), .S(n29388), .Q(n18036)
         );
  MUX21X1 U33010 ( .IN1(n34625), .IN2(s15_data_o[14]), .S(n29388), .Q(n18035)
         );
  MUX21X1 U33011 ( .IN1(n34562), .IN2(s15_data_o[15]), .S(n29388), .Q(n18034)
         );
  NAND2X0 U33012 ( .IN1(\s0/msel/gnt_p3 [1]), .IN2(n29445), .QN(n29413) );
  OA21X1 U33013 ( .IN1(\s0/msel/gnt_p3 [1]), .IN2(n29431), .IN3(n29413), .Q(
        n29465) );
  NAND2X0 U33014 ( .IN1(\s0/msel/gnt_p3 [1]), .IN2(n29436), .QN(n29412) );
  OA21X1 U33015 ( .IN1(\s0/msel/gnt_p3 [1]), .IN2(n29422), .IN3(n29412), .Q(
        n29468) );
  NOR2X0 U33016 ( .IN1(\s0/msel/gnt_p3 [0]), .IN2(n29468), .QN(n29389) );
  NOR2X0 U33017 ( .IN1(\s0/msel/gnt_p3 [1]), .IN2(n29398), .QN(n29403) );
  NOR2X0 U33018 ( .IN1(n29389), .IN2(n29403), .QN(n29391) );
  NAND2X0 U33019 ( .IN1(n29397), .IN2(n29400), .QN(n29390) );
  NAND3X0 U33020 ( .IN1(n29465), .IN2(n29391), .IN3(n29390), .QN(n29396) );
  NOR2X0 U33021 ( .IN1(n34259), .IN2(n34423), .QN(n29392) );
  OA21X1 U33022 ( .IN1(n29392), .IN2(n29400), .IN3(n34549), .Q(n29410) );
  INVX0 U33023 ( .INP(n29392), .ZN(n29447) );
  AO21X1 U33024 ( .IN1(n29459), .IN2(n34259), .IN3(n29461), .Q(n29411) );
  OA222X1 U33025 ( .IN1(n29447), .IN2(n29433), .IN3(n34423), .IN4(
        \s0/msel/gnt_p3 [0]), .IN5(n29411), .IN6(\s0/msel/gnt_p3 [1]), .Q(
        n29393) );
  NOR2X0 U33026 ( .IN1(n29394), .IN2(n29393), .QN(n29395) );
  AO22X1 U33027 ( .IN1(\s0/msel/gnt_p3 [2]), .IN2(n29396), .IN3(n29410), .IN4(
        n29395), .Q(n18033) );
  NOR2X0 U33028 ( .IN1(\s0/msel/gnt_p3 [1]), .IN2(n29460), .QN(n29443) );
  INVX0 U33029 ( .INP(n29397), .ZN(n29399) );
  OA21X1 U33030 ( .IN1(n29443), .IN2(n29399), .IN3(n29398), .Q(n29409) );
  INVX0 U33031 ( .INP(n29445), .ZN(n29424) );
  NAND2X0 U33032 ( .IN1(\s0/msel/gnt_p3 [1]), .IN2(n34259), .QN(n29439) );
  AO221X1 U33033 ( .IN1(n29424), .IN2(n29408), .IN3(n29424), .IN4(n29399), 
        .IN5(n29439), .Q(n29406) );
  AO221X1 U33034 ( .IN1(n29400), .IN2(n29408), .IN3(n29400), .IN4(n29447), 
        .IN5(n29399), .Q(n29402) );
  NAND2X0 U33035 ( .IN1(n34259), .IN2(n34423), .QN(n29450) );
  INVX0 U33036 ( .INP(n29450), .ZN(n29401) );
  INVX0 U33037 ( .INP(n29431), .ZN(n29414) );
  AO222X1 U33038 ( .IN1(n29402), .IN2(n29409), .IN3(n29402), .IN4(n29450), 
        .IN5(n29401), .IN6(n29414), .Q(n29405) );
  NAND2X0 U33039 ( .IN1(\s0/msel/gnt_p3 [0]), .IN2(n29403), .QN(n29404) );
  AND4X1 U33040 ( .IN1(\s0/msel/gnt_p3 [2]), .IN2(n29406), .IN3(n29405), .IN4(
        n29404), .Q(n29407) );
  AO221X1 U33041 ( .IN1(n29410), .IN2(n29409), .IN3(n29410), .IN4(n29408), 
        .IN5(n29407), .Q(n29417) );
  INVX0 U33042 ( .INP(n29433), .ZN(n29420) );
  OA21X1 U33043 ( .IN1(n29420), .IN2(n29447), .IN3(n34549), .Q(n29464) );
  OA21X1 U33044 ( .IN1(n29411), .IN2(n29417), .IN3(n29464), .Q(n29419) );
  INVX0 U33045 ( .INP(n29422), .ZN(n29449) );
  OA21X1 U33046 ( .IN1(n29449), .IN2(n29417), .IN3(n29412), .Q(n29416) );
  OA21X1 U33047 ( .IN1(n29414), .IN2(n29417), .IN3(n29413), .Q(n29415) );
  OA221X1 U33048 ( .IN1(\s0/msel/gnt_p3 [0]), .IN2(n29416), .IN3(n34259), 
        .IN4(n29415), .IN5(\s0/msel/gnt_p3 [2]), .Q(n29418) );
  OAI22X1 U33049 ( .IN1(n29419), .IN2(n29418), .IN3(n34423), .IN4(n29417), 
        .QN(n18032) );
  NOR2X0 U33050 ( .IN1(n29459), .IN2(n29460), .QN(n29428) );
  INVX0 U33051 ( .INP(n29428), .ZN(n29421) );
  NOR2X0 U33052 ( .IN1(n29421), .IN2(n29420), .QN(n29427) );
  NAND2X0 U33053 ( .IN1(n29431), .IN2(n34259), .QN(n29423) );
  NAND3X0 U33054 ( .IN1(n29423), .IN2(n29422), .IN3(n29428), .QN(n29425) );
  INVX0 U33055 ( .INP(n29461), .ZN(n29434) );
  OA21X1 U33056 ( .IN1(n29459), .IN2(n29434), .IN3(n29424), .Q(n29441) );
  NAND2X0 U33057 ( .IN1(n29425), .IN2(n29441), .QN(n29426) );
  NOR2X0 U33058 ( .IN1(n29427), .IN2(n29426), .QN(n29430) );
  NAND2X0 U33059 ( .IN1(\s0/msel/gnt_p3 [0]), .IN2(n29428), .QN(n29429) );
  OA221X1 U33060 ( .IN1(n29436), .IN2(n29441), .IN3(n29436), .IN4(n29429), 
        .IN5(n29431), .Q(n29448) );
  OA22X1 U33061 ( .IN1(n29436), .IN2(n29430), .IN3(n29448), .IN4(n29450), .Q(
        n29458) );
  NOR2X0 U33062 ( .IN1(n29449), .IN2(n29431), .QN(n29432) );
  NOR2X0 U33063 ( .IN1(n29433), .IN2(n29432), .QN(n29437) );
  OA21X1 U33064 ( .IN1(n29460), .IN2(n29437), .IN3(n29434), .Q(n29451) );
  NOR3X0 U33065 ( .IN1(n29451), .IN2(n29459), .IN3(n29447), .QN(n29435) );
  NOR2X0 U33066 ( .IN1(n29435), .IN2(n34549), .QN(n29457) );
  NOR2X0 U33067 ( .IN1(n29449), .IN2(n29436), .QN(n29444) );
  INVX0 U33068 ( .INP(n29444), .ZN(n29440) );
  OR3X1 U33069 ( .IN1(n29459), .IN2(n29440), .IN3(n34259), .Q(n29438) );
  NAND2X0 U33070 ( .IN1(n29438), .IN2(n29437), .QN(n29446) );
  INVX0 U33071 ( .INP(n29446), .ZN(n29442) );
  AO221X1 U33072 ( .IN1(n29442), .IN2(n29441), .IN3(n29442), .IN4(n29440), 
        .IN5(n29439), .Q(n29456) );
  OA221X1 U33073 ( .IN1(n29446), .IN2(n29445), .IN3(n29446), .IN4(n29444), 
        .IN5(n29443), .Q(n29454) );
  NOR3X0 U33074 ( .IN1(n29449), .IN2(n29448), .IN3(n29447), .QN(n29453) );
  NOR2X0 U33075 ( .IN1(n29451), .IN2(n29450), .QN(n29452) );
  NOR4X0 U33076 ( .IN1(\s0/msel/gnt_p3 [2]), .IN2(n29454), .IN3(n29453), .IN4(
        n29452), .QN(n29455) );
  AO22X1 U33077 ( .IN1(n29458), .IN2(n29457), .IN3(n29456), .IN4(n29455), .Q(
        n29466) );
  AO221X1 U33078 ( .IN1(\s0/msel/gnt_p3 [1]), .IN2(n29460), .IN3(n34423), 
        .IN4(n29459), .IN5(n29466), .Q(n29463) );
  NAND3X0 U33079 ( .IN1(\s0/msel/gnt_p3 [0]), .IN2(n29461), .IN3(n34423), .QN(
        n29462) );
  NAND3X0 U33080 ( .IN1(n29464), .IN2(n29463), .IN3(n29462), .QN(n29471) );
  NOR2X0 U33081 ( .IN1(n29465), .IN2(n34259), .QN(n29470) );
  INVX0 U33082 ( .INP(n29466), .ZN(n29467) );
  OA221X1 U33083 ( .IN1(\s0/msel/gnt_p3 [0]), .IN2(\s0/msel/gnt_p3 [2]), .IN3(
        \s0/msel/gnt_p3 [0]), .IN4(n29468), .IN5(n29467), .Q(n29469) );
  AO221X1 U33084 ( .IN1(n29471), .IN2(n29470), .IN3(n29471), .IN4(n34549), 
        .IN5(n29469), .Q(n18031) );
  INVX0 U33085 ( .INP(n29506), .ZN(n29529) );
  INVX0 U33086 ( .INP(n29519), .ZN(n29516) );
  MUX21X1 U33087 ( .IN1(n29529), .IN2(n29516), .S(\s0/msel/gnt_p1 [1]), .Q(
        n29545) );
  NAND3X0 U33088 ( .IN1(\s0/msel/gnt_p1 [2]), .IN2(n29545), .IN3(n34250), .QN(
        n29479) );
  NAND2X0 U33089 ( .IN1(\s0/msel/gnt_p1 [1]), .IN2(n29508), .QN(n29543) );
  NAND2X0 U33090 ( .IN1(n34669), .IN2(n29515), .QN(n29542) );
  INVX0 U33091 ( .INP(n29472), .ZN(n29473) );
  AO221X1 U33092 ( .IN1(n29543), .IN2(n29490), .IN3(n29543), .IN4(n29542), 
        .IN5(n29473), .Q(n29474) );
  NAND2X0 U33093 ( .IN1(\s0/msel/gnt_p1 [2]), .IN2(n29474), .QN(n29478) );
  NAND2X0 U33094 ( .IN1(\s0/msel/gnt_p1 [1]), .IN2(n34250), .QN(n29532) );
  OA22X1 U33095 ( .IN1(n29526), .IN2(n29532), .IN3(n29507), .IN4(n34669), .Q(
        n29496) );
  OA21X1 U33096 ( .IN1(\s0/msel/gnt_p1 [0]), .IN2(n29527), .IN3(n29509), .Q(
        n29498) );
  OA22X1 U33097 ( .IN1(\s0/msel/gnt_p1 [1]), .IN2(n29498), .IN3(
        \s0/msel/gnt_p1 [1]), .IN4(n29485), .Q(n29476) );
  NAND4X0 U33098 ( .IN1(n29496), .IN2(n29476), .IN3(n34432), .IN4(n29475), 
        .QN(n29477) );
  NAND3X0 U33099 ( .IN1(n29479), .IN2(n29478), .IN3(n29477), .QN(n18030) );
  OA21X1 U33100 ( .IN1(n29481), .IN2(n29490), .IN3(n29480), .Q(n29484) );
  OAI21X1 U33101 ( .IN1(n29486), .IN2(n29482), .IN3(n29485), .QN(n29483) );
  AO221X1 U33102 ( .IN1(\s0/msel/gnt_p1 [1]), .IN2(n29484), .IN3(n34669), 
        .IN4(n29483), .IN5(n29520), .Q(n29495) );
  NOR2X0 U33103 ( .IN1(n29485), .IN2(n29487), .QN(n29493) );
  INVX0 U33104 ( .INP(n29508), .ZN(n29489) );
  NAND3X0 U33105 ( .IN1(\s0/msel/gnt_p1 [0]), .IN2(n34669), .IN3(n29519), .QN(
        n29531) );
  NOR2X0 U33106 ( .IN1(n29487), .IN2(n29486), .QN(n29488) );
  OA22X1 U33107 ( .IN1(n29489), .IN2(n29531), .IN3(n29488), .IN4(n29543), .Q(
        n29492) );
  OA21X1 U33108 ( .IN1(n29493), .IN2(n29490), .IN3(n29515), .Q(n29491) );
  NAND2X0 U33109 ( .IN1(n34250), .IN2(n34669), .QN(n29521) );
  OA22X1 U33110 ( .IN1(n29493), .IN2(n29492), .IN3(n29491), .IN4(n29521), .Q(
        n29494) );
  MUX21X1 U33111 ( .IN1(n29495), .IN2(n29494), .S(\s0/msel/gnt_p1 [2]), .Q(
        n29505) );
  NAND2X0 U33112 ( .IN1(n29496), .IN2(n34432), .QN(n29497) );
  AO21X1 U33113 ( .IN1(n29498), .IN2(n29505), .IN3(n29497), .Q(n29504) );
  NOR2X0 U33114 ( .IN1(n29532), .IN2(n29519), .QN(n29502) );
  NOR2X0 U33115 ( .IN1(n29506), .IN2(\s0/msel/gnt_p1 [0]), .QN(n29500) );
  NAND2X0 U33116 ( .IN1(n29505), .IN2(n29515), .QN(n29499) );
  NOR2X0 U33117 ( .IN1(n29500), .IN2(n29499), .QN(n29501) );
  OR3X1 U33118 ( .IN1(n29502), .IN2(n29501), .IN3(n34432), .Q(n29503) );
  AO22X1 U33119 ( .IN1(\s0/msel/gnt_p1 [1]), .IN2(n29505), .IN3(n29504), .IN4(
        n29503), .Q(n18029) );
  AO221X1 U33120 ( .IN1(\s0/msel/gnt_p1 [1]), .IN2(n29507), .IN3(n34669), 
        .IN4(n29509), .IN5(n34250), .Q(n29541) );
  NOR2X0 U33121 ( .IN1(\s0/msel/gnt_p1 [1]), .IN2(n29527), .QN(n29540) );
  NAND2X0 U33122 ( .IN1(n29519), .IN2(n29506), .QN(n29510) );
  OA21X1 U33123 ( .IN1(n29529), .IN2(n29515), .IN3(n29507), .Q(n29530) );
  OA21X1 U33124 ( .IN1(n34250), .IN2(n29510), .IN3(n29530), .Q(n29512) );
  OA21X1 U33125 ( .IN1(n29514), .IN2(n29512), .IN3(n29509), .Q(n29524) );
  INVX0 U33126 ( .INP(n29527), .ZN(n29525) );
  AND2X1 U33127 ( .IN1(n29525), .IN2(n29530), .Q(n29511) );
  OA21X1 U33128 ( .IN1(n29509), .IN2(n29525), .IN3(n29508), .Q(n29534) );
  OA22X1 U33129 ( .IN1(n29512), .IN2(n29511), .IN3(n29534), .IN4(n29510), .Q(
        n29513) );
  OA22X1 U33130 ( .IN1(n29524), .IN2(n29521), .IN3(n29514), .IN4(n29513), .Q(
        n29518) );
  OA21X1 U33131 ( .IN1(n29516), .IN2(n29534), .IN3(n29515), .Q(n29523) );
  OR4X1 U33132 ( .IN1(n34669), .IN2(n34250), .IN3(n29529), .IN4(n29523), .Q(
        n29517) );
  NAND3X0 U33133 ( .IN1(n34432), .IN2(n29518), .IN3(n29517), .QN(n29539) );
  NAND4X0 U33134 ( .IN1(n29520), .IN2(n29527), .IN3(n29526), .IN4(n29519), 
        .QN(n29522) );
  AO21X1 U33135 ( .IN1(n29523), .IN2(n29522), .IN3(n29521), .Q(n29537) );
  OR3X1 U33136 ( .IN1(n34669), .IN2(n29525), .IN3(n29524), .Q(n29536) );
  NAND2X0 U33137 ( .IN1(n29527), .IN2(n29526), .QN(n29528) );
  AO22X1 U33138 ( .IN1(n29534), .IN2(n29533), .IN3(n29532), .IN4(n29531), .Q(
        n29535) );
  NAND4X0 U33139 ( .IN1(\s0/msel/gnt_p1 [2]), .IN2(n29537), .IN3(n29536), 
        .IN4(n29535), .QN(n29538) );
  NAND2X0 U33140 ( .IN1(n29539), .IN2(n29538), .QN(n29544) );
  AO221X1 U33141 ( .IN1(n29541), .IN2(n29540), .IN3(n29541), .IN4(n29544), 
        .IN5(\s0/msel/gnt_p1 [2]), .Q(n29548) );
  NAND4X0 U33142 ( .IN1(\s0/msel/gnt_p1 [2]), .IN2(\s0/msel/gnt_p1 [0]), .IN3(
        n29543), .IN4(n29542), .QN(n29547) );
  AO221X1 U33143 ( .IN1(n34250), .IN2(n29545), .IN3(n34250), .IN4(n34432), 
        .IN5(n29544), .Q(n29546) );
  NAND3X0 U33144 ( .IN1(n29548), .IN2(n29547), .IN3(n29546), .QN(n18028) );
  NAND2X0 U33145 ( .IN1(\s0/msel/gnt_p0 [1]), .IN2(n34240), .QN(n29551) );
  INVX0 U33146 ( .INP(n29551), .ZN(n29574) );
  NAND3X0 U33147 ( .IN1(n13787), .IN2(n13761), .IN3(m2s0_cyc), .QN(n29594) );
  INVX0 U33148 ( .INP(n29594), .ZN(n29609) );
  NAND2X0 U33149 ( .IN1(n29574), .IN2(n29609), .QN(n29549) );
  NAND3X0 U33150 ( .IN1(n13735), .IN2(n13709), .IN3(m3s0_cyc), .QN(n29591) );
  NAND2X0 U33151 ( .IN1(\s0/msel/gnt_p0 [0]), .IN2(\s0/msel/gnt_p0 [1]), .QN(
        n29552) );
  OR2X1 U33152 ( .IN1(n29591), .IN2(n29552), .Q(n29622) );
  NAND3X0 U33153 ( .IN1(n29549), .IN2(n29622), .IN3(n34440), .QN(n29582) );
  NAND3X0 U33154 ( .IN1(n13896), .IN2(n13865), .IN3(m0s0_cyc), .QN(n29595) );
  NAND3X0 U33155 ( .IN1(n13839), .IN2(n13813), .IN3(m1s0_cyc), .QN(n29625) );
  MUX21X1 U33156 ( .IN1(n29595), .IN2(n29625), .S(\s0/msel/gnt_p0 [0]), .Q(
        n29584) );
  NAND3X0 U33157 ( .IN1(n13631), .IN2(n13605), .IN3(m5s0_cyc), .QN(n29597) );
  NAND3X0 U33158 ( .IN1(n13683), .IN2(n13657), .IN3(m4s0_cyc), .QN(n29605) );
  NAND2X0 U33159 ( .IN1(n29597), .IN2(n29605), .QN(n29565) );
  NAND3X0 U33160 ( .IN1(n13527), .IN2(n13471), .IN3(m7s0_cyc), .QN(n29596) );
  NAND3X0 U33161 ( .IN1(n13579), .IN2(n13553), .IN3(m6s0_cyc), .QN(n29606) );
  NAND2X0 U33162 ( .IN1(n29596), .IN2(n29606), .QN(n29572) );
  OAI22X1 U33163 ( .IN1(\s0/msel/gnt_p0 [1]), .IN2(n29584), .IN3(n29565), 
        .IN4(n29572), .QN(n29550) );
  NOR2X0 U33164 ( .IN1(n29582), .IN2(n29550), .QN(n29555) );
  INVX0 U33165 ( .INP(n29591), .ZN(n29575) );
  INVX0 U33166 ( .INP(n29625), .ZN(n29592) );
  NAND2X0 U33167 ( .IN1(n34240), .IN2(n34453), .QN(n29612) );
  NOR2X0 U33168 ( .IN1(\s0/msel/gnt_p0 [1]), .IN2(n34240), .QN(n29566) );
  INVX0 U33169 ( .INP(n29566), .ZN(n29624) );
  OA21X1 U33170 ( .IN1(n29592), .IN2(n29612), .IN3(n29624), .Q(n29569) );
  NAND2X0 U33171 ( .IN1(n29594), .IN2(n29591), .QN(n29579) );
  OA22X1 U33172 ( .IN1(n29575), .IN2(n29551), .IN3(n29569), .IN4(n29579), .Q(
        n29553) );
  NAND2X0 U33173 ( .IN1(n29553), .IN2(n29552), .QN(n29554) );
  NAND2X0 U33174 ( .IN1(n29555), .IN2(n29554), .QN(n29564) );
  INVX0 U33175 ( .INP(n29595), .ZN(n29623) );
  NOR2X0 U33176 ( .IN1(n29623), .IN2(n29609), .QN(n29598) );
  AND3X1 U33177 ( .IN1(n29598), .IN2(n29625), .IN3(n29591), .Q(n29559) );
  NAND2X0 U33178 ( .IN1(n34453), .IN2(n29597), .QN(n29627) );
  NOR2X0 U33179 ( .IN1(n29572), .IN2(n29627), .QN(n29557) );
  NAND2X0 U33180 ( .IN1(\s0/msel/gnt_p0 [1]), .IN2(n29596), .QN(n29628) );
  INVX0 U33181 ( .INP(n29628), .ZN(n29556) );
  NOR2X0 U33182 ( .IN1(n29557), .IN2(n29556), .QN(n29558) );
  NOR2X0 U33183 ( .IN1(n29559), .IN2(n29558), .QN(n29561) );
  INVX0 U33184 ( .INP(n29605), .ZN(n29615) );
  INVX0 U33185 ( .INP(n29606), .ZN(n29600) );
  MUX21X1 U33186 ( .IN1(n29615), .IN2(n29600), .S(\s0/msel/gnt_p0 [1]), .Q(
        n29630) );
  NAND2X0 U33187 ( .IN1(n34240), .IN2(n29630), .QN(n29560) );
  NAND2X0 U33188 ( .IN1(n29561), .IN2(n29560), .QN(n29562) );
  NAND2X0 U33189 ( .IN1(\s0/msel/gnt_p0 [2]), .IN2(n29562), .QN(n29563) );
  NAND2X0 U33190 ( .IN1(n29564), .IN2(n29563), .QN(n18027) );
  INVX0 U33191 ( .INP(n29565), .ZN(n29571) );
  NOR2X0 U33192 ( .IN1(n29623), .IN2(n29592), .QN(n29580) );
  NAND3X0 U33193 ( .IN1(n29566), .IN2(n29596), .IN3(n29606), .QN(n29567) );
  OA221X1 U33194 ( .IN1(n29628), .IN2(n29571), .IN3(n29628), .IN4(n29580), 
        .IN5(n29567), .Q(n29568) );
  AO221X1 U33195 ( .IN1(n29568), .IN2(n29572), .IN3(n29568), .IN4(n29612), 
        .IN5(n34440), .Q(n29581) );
  INVX0 U33196 ( .INP(n29569), .ZN(n29570) );
  OAI221X1 U33197 ( .IN1(n29579), .IN2(n29572), .IN3(n29579), .IN4(n29571), 
        .IN5(n29570), .QN(n29578) );
  OR2X1 U33198 ( .IN1(n29572), .IN2(n29580), .Q(n29573) );
  NAND4X0 U33199 ( .IN1(\s0/msel/gnt_p0 [1]), .IN2(n29605), .IN3(n29597), 
        .IN4(n29573), .QN(n29577) );
  NAND2X0 U33200 ( .IN1(n29575), .IN2(n29574), .QN(n29576) );
  NAND4X0 U33201 ( .IN1(n34440), .IN2(n29578), .IN3(n29577), .IN4(n29576), 
        .QN(n29583) );
  OA221X1 U33202 ( .IN1(n29581), .IN2(n29580), .IN3(n29581), .IN4(n29579), 
        .IN5(n29583), .Q(n29590) );
  AO21X1 U33203 ( .IN1(n29584), .IN2(n29583), .IN3(n29582), .Q(n29589) );
  NAND2X0 U33204 ( .IN1(n29615), .IN2(n34240), .QN(n29585) );
  NAND3X0 U33205 ( .IN1(n29585), .IN2(n29597), .IN3(n29590), .QN(n29587) );
  NAND3X0 U33206 ( .IN1(\s0/msel/gnt_p0 [1]), .IN2(n29600), .IN3(n34240), .QN(
        n29586) );
  NAND3X0 U33207 ( .IN1(\s0/msel/gnt_p0 [2]), .IN2(n29587), .IN3(n29586), .QN(
        n29588) );
  AO22X1 U33208 ( .IN1(\s0/msel/gnt_p0 [1]), .IN2(n29590), .IN3(n29589), .IN4(
        n29588), .Q(n18026) );
  OA21X1 U33209 ( .IN1(n29597), .IN2(n29615), .IN3(n29591), .Q(n29611) );
  INVX0 U33210 ( .INP(n29611), .ZN(n29593) );
  AO21X1 U33211 ( .IN1(n29594), .IN2(n29593), .IN3(n29592), .Q(n29613) );
  NAND3X0 U33212 ( .IN1(\s0/msel/gnt_p0 [1]), .IN2(n29613), .IN3(n29595), .QN(
        n29604) );
  OA21X1 U33213 ( .IN1(n29623), .IN2(n29625), .IN3(n29596), .Q(n29608) );
  OA21X1 U33214 ( .IN1(n29608), .IN2(n29600), .IN3(n29597), .Q(n29616) );
  OR2X1 U33215 ( .IN1(n29612), .IN2(n29616), .Q(n29603) );
  INVX0 U33216 ( .INP(n29598), .ZN(n29599) );
  AO221X1 U33217 ( .IN1(n29611), .IN2(n29615), .IN3(n29611), .IN4(n34240), 
        .IN5(n29599), .Q(n29601) );
  AO21X1 U33218 ( .IN1(n29608), .IN2(n29601), .IN3(n29600), .Q(n29602) );
  NAND4X0 U33219 ( .IN1(\s0/msel/gnt_p0 [2]), .IN2(n29604), .IN3(n29603), 
        .IN4(n29602), .QN(n29621) );
  NAND2X0 U33220 ( .IN1(n29606), .IN2(n29605), .QN(n29607) );
  AO221X1 U33221 ( .IN1(n29608), .IN2(n29623), .IN3(n29608), .IN4(n34240), 
        .IN5(n29607), .Q(n29610) );
  AO21X1 U33222 ( .IN1(n29611), .IN2(n29610), .IN3(n29609), .Q(n29619) );
  INVX0 U33223 ( .INP(n29612), .ZN(n29614) );
  NAND2X0 U33224 ( .IN1(n29614), .IN2(n29613), .QN(n29618) );
  OR4X1 U33225 ( .IN1(n34453), .IN2(n34240), .IN3(n29616), .IN4(n29615), .Q(
        n29617) );
  NAND4X0 U33226 ( .IN1(n34440), .IN2(n29619), .IN3(n29618), .IN4(n29617), 
        .QN(n29620) );
  NAND2X0 U33227 ( .IN1(n29621), .IN2(n29620), .QN(n29629) );
  OA221X1 U33228 ( .IN1(n29629), .IN2(n29623), .IN3(n29629), .IN4(n34453), 
        .IN5(n29622), .Q(n29626) );
  AO221X1 U33229 ( .IN1(n29626), .IN2(n29625), .IN3(n29626), .IN4(n29624), 
        .IN5(\s0/msel/gnt_p0 [2]), .Q(n29633) );
  NAND4X0 U33230 ( .IN1(\s0/msel/gnt_p0 [2]), .IN2(\s0/msel/gnt_p0 [0]), .IN3(
        n29628), .IN4(n29627), .QN(n29632) );
  AO221X1 U33231 ( .IN1(n34240), .IN2(n34440), .IN3(n34240), .IN4(n29630), 
        .IN5(n29629), .Q(n29631) );
  NAND3X0 U33232 ( .IN1(n29633), .IN2(n29632), .IN3(n29631), .QN(n18025) );
  INVX0 U33233 ( .INP(n29685), .ZN(n29679) );
  MUX21X1 U33234 ( .IN1(n29664), .IN2(n29679), .S(\s0/msel/gnt_p2 [1]), .Q(
        n29728) );
  MUX21X1 U33235 ( .IN1(n29647), .IN2(n29654), .S(\s0/msel/gnt_p2 [1]), .Q(
        n29678) );
  OA22X1 U33236 ( .IN1(\s0/msel/gnt_p2 [0]), .IN2(n29678), .IN3(
        \s0/msel/gnt_p2 [1]), .IN4(n29634), .Q(n29636) );
  NAND2X0 U33237 ( .IN1(n29636), .IN2(n29635), .QN(n29643) );
  NAND2X0 U33238 ( .IN1(\s0/msel/gnt_p2 [0]), .IN2(\s0/msel/gnt_p2 [1]), .QN(
        n29672) );
  INVX0 U33239 ( .INP(n29672), .ZN(n29656) );
  NAND2X0 U33240 ( .IN1(n29637), .IN2(n29656), .QN(n29723) );
  NOR2X0 U33241 ( .IN1(\s0/msel/gnt_p2 [0]), .IN2(n34286), .QN(n29655) );
  NAND2X0 U33242 ( .IN1(n29688), .IN2(n29655), .QN(n29638) );
  AND3X1 U33243 ( .IN1(n34473), .IN2(n29723), .IN3(n29638), .Q(n29652) );
  INVX0 U33244 ( .INP(n29695), .ZN(n29719) );
  INVX0 U33245 ( .INP(n29686), .ZN(n29717) );
  MUX21X1 U33246 ( .IN1(n29719), .IN2(n29717), .S(\s0/msel/gnt_p2 [0]), .Q(
        n29653) );
  NAND2X0 U33247 ( .IN1(n34286), .IN2(n29653), .QN(n29641) );
  AND2X1 U33248 ( .IN1(n34286), .IN2(n29686), .Q(n29651) );
  AO22X1 U33249 ( .IN1(n29660), .IN2(n29651), .IN3(\s0/msel/gnt_p2 [1]), .IN4(
        n29680), .Q(n29639) );
  AND4X1 U33250 ( .IN1(n29652), .IN2(n29641), .IN3(n29640), .IN4(n29639), .Q(
        n29642) );
  AO221X1 U33251 ( .IN1(\s0/msel/gnt_p2 [2]), .IN2(n29728), .IN3(
        \s0/msel/gnt_p2 [2]), .IN4(n29643), .IN5(n29642), .Q(n18024) );
  NAND2X0 U33252 ( .IN1(n29644), .IN2(n29646), .QN(n29648) );
  NAND2X0 U33253 ( .IN1(n29660), .IN2(n29648), .QN(n29650) );
  NOR2X0 U33254 ( .IN1(n29704), .IN2(n29672), .QN(n29714) );
  OA21X1 U33255 ( .IN1(n29646), .IN2(n29645), .IN3(n29697), .Q(n29662) );
  NAND4X0 U33256 ( .IN1(n29697), .IN2(n29695), .IN3(n29686), .IN4(n29647), 
        .QN(n29658) );
  NAND3X0 U33257 ( .IN1(n29680), .IN2(n29658), .IN3(n29648), .QN(n29649) );
  AOI222X1 U33258 ( .IN1(n29651), .IN2(n29650), .IN3(n29714), .IN4(n29662), 
        .IN5(n29649), .IN6(n29655), .QN(n29668) );
  OA21X1 U33259 ( .IN1(n29668), .IN2(n29653), .IN3(n29652), .Q(n29677) );
  NOR2X0 U33260 ( .IN1(n34473), .IN2(n34290), .QN(n29727) );
  INVX0 U33261 ( .INP(n29654), .ZN(n29699) );
  NOR2X0 U33262 ( .IN1(n29699), .IN2(\s0/msel/gnt_p2 [1]), .QN(n29657) );
  NOR2X0 U33263 ( .IN1(n29655), .IN2(n29657), .QN(n29706) );
  NOR2X0 U33264 ( .IN1(n29679), .IN2(n29706), .QN(n29659) );
  AO222X1 U33265 ( .IN1(n29659), .IN2(n29658), .IN3(n29659), .IN4(n29657), 
        .IN5(n29658), .IN6(n29656), .Q(n29666) );
  OR2X1 U33266 ( .IN1(n29661), .IN2(n29660), .Q(n29665) );
  NOR2X0 U33267 ( .IN1(\s0/msel/gnt_p2 [0]), .IN2(\s0/msel/gnt_p2 [1]), .QN(
        n29694) );
  INVX0 U33268 ( .INP(n29694), .ZN(n29702) );
  NOR2X0 U33269 ( .IN1(n29662), .IN2(n29702), .QN(n29663) );
  AO22X1 U33270 ( .IN1(n29666), .IN2(n29665), .IN3(n29664), .IN4(n29663), .Q(
        n29667) );
  MUX21X1 U33271 ( .IN1(n29668), .IN2(n29667), .S(\s0/msel/gnt_p2 [2]), .Q(
        n29675) );
  NOR2X0 U33272 ( .IN1(n29675), .IN2(n29704), .QN(n29671) );
  NAND2X0 U33273 ( .IN1(\s0/msel/gnt_p2 [1]), .IN2(n29699), .QN(n29669) );
  NAND2X0 U33274 ( .IN1(n29669), .IN2(\s0/msel/gnt_p2 [2]), .QN(n29670) );
  NOR2X0 U33275 ( .IN1(n29671), .IN2(n29670), .QN(n29673) );
  OA22X1 U33276 ( .IN1(n29727), .IN2(n29673), .IN3(n29672), .IN4(n29685), .Q(
        n29676) );
  AOI21X1 U33277 ( .IN1(n29697), .IN2(n29727), .IN3(\s0/msel/gnt_p2 [1]), .QN(
        n29674) );
  OAI22X1 U33278 ( .IN1(n29677), .IN2(n29676), .IN3(n29675), .IN4(n29674), 
        .QN(n18023) );
  AO21X1 U33279 ( .IN1(\s0/msel/gnt_p2 [2]), .IN2(n29678), .IN3(
        \s0/msel/gnt_p2 [0]), .Q(n29726) );
  NOR2X0 U33280 ( .IN1(n29699), .IN2(n29704), .QN(n29683) );
  NAND3X0 U33281 ( .IN1(n29716), .IN2(n29679), .IN3(n29683), .QN(n29682) );
  INVX0 U33282 ( .INP(n29683), .ZN(n29687) );
  OA21X1 U33283 ( .IN1(n29704), .IN2(n29697), .IN3(n29680), .Q(n29705) );
  OA21X1 U33284 ( .IN1(n34290), .IN2(n29687), .IN3(n29705), .Q(n29681) );
  OA21X1 U33285 ( .IN1(n29688), .IN2(n29681), .IN3(n29686), .Q(n29700) );
  NAND2X0 U33286 ( .IN1(n29682), .IN2(n29700), .QN(n29693) );
  NAND3X0 U33287 ( .IN1(n29683), .IN2(\s0/msel/gnt_p2 [0]), .IN3(n29695), .QN(
        n29684) );
  NAND2X0 U33288 ( .IN1(n29684), .IN2(n29705), .QN(n29691) );
  OA21X1 U33289 ( .IN1(n29719), .IN2(n29686), .IN3(n29685), .Q(n29707) );
  NOR2X0 U33290 ( .IN1(n29707), .IN2(n29687), .QN(n29690) );
  NOR2X0 U33291 ( .IN1(\s0/msel/gnt_p2 [1]), .IN2(n29688), .QN(n29689) );
  OA22X1 U33292 ( .IN1(n29691), .IN2(n29690), .IN3(n29689), .IN4(n34290), .Q(
        n29692) );
  AO221X1 U33293 ( .IN1(n29694), .IN2(n29693), .IN3(n29702), .IN4(n29692), 
        .IN5(\s0/msel/gnt_p2 [2]), .Q(n29715) );
  NAND2X0 U33294 ( .IN1(n29716), .IN2(n29695), .QN(n29703) );
  INVX0 U33295 ( .INP(n29703), .ZN(n29696) );
  NAND2X0 U33296 ( .IN1(\s0/msel/gnt_p2 [0]), .IN2(n29696), .QN(n29698) );
  OA221X1 U33297 ( .IN1(n29699), .IN2(n29698), .IN3(n29699), .IN4(n29707), 
        .IN5(n29697), .Q(n29701) );
  INVX0 U33298 ( .INP(n29701), .ZN(n29713) );
  OR3X1 U33299 ( .IN1(n34286), .IN2(n29719), .IN3(n29700), .Q(n29711) );
  OR2X1 U33300 ( .IN1(n29702), .IN2(n29701), .Q(n29710) );
  AO221X1 U33301 ( .IN1(n29705), .IN2(n29704), .IN3(n29705), .IN4(n34290), 
        .IN5(n29703), .Q(n29708) );
  AO21X1 U33302 ( .IN1(n29708), .IN2(n29707), .IN3(n29706), .Q(n29709) );
  NAND4X0 U33303 ( .IN1(\s0/msel/gnt_p2 [2]), .IN2(n29711), .IN3(n29710), 
        .IN4(n29709), .QN(n29712) );
  OA221X1 U33304 ( .IN1(n29715), .IN2(n29714), .IN3(n29715), .IN4(n29713), 
        .IN5(n29712), .Q(n29725) );
  NAND3X0 U33305 ( .IN1(\s0/msel/gnt_p2 [1]), .IN2(n29725), .IN3(n29716), .QN(
        n29722) );
  NAND2X0 U33306 ( .IN1(\s0/msel/gnt_p2 [0]), .IN2(n29717), .QN(n29720) );
  INVX0 U33307 ( .INP(n29725), .ZN(n29718) );
  AO221X1 U33308 ( .IN1(n29720), .IN2(n29719), .IN3(n29720), .IN4(n29718), 
        .IN5(\s0/msel/gnt_p2 [1]), .Q(n29721) );
  NAND3X0 U33309 ( .IN1(n29723), .IN2(n29722), .IN3(n29721), .QN(n29724) );
  AO222X1 U33310 ( .IN1(n29728), .IN2(n29727), .IN3(n29726), .IN4(n29725), 
        .IN5(n29724), .IN6(n34473), .Q(n18022) );
  NOR2X0 U33311 ( .IN1(n29729), .IN2(n34379), .QN(n29730) );
  MUX21X1 U33312 ( .IN1(n34294), .IN2(s15_data_o[0]), .S(n29730), .Q(n18021)
         );
  MUX21X1 U33313 ( .IN1(n34557), .IN2(s15_data_o[1]), .S(n29730), .Q(n18020)
         );
  MUX21X1 U33314 ( .IN1(n34293), .IN2(s15_data_o[2]), .S(n29730), .Q(n18019)
         );
  MUX21X1 U33315 ( .IN1(n34555), .IN2(s15_data_o[3]), .S(n29730), .Q(n18018)
         );
  MUX21X1 U33316 ( .IN1(n34297), .IN2(s15_data_o[4]), .S(n29730), .Q(n18017)
         );
  MUX21X1 U33317 ( .IN1(n34558), .IN2(s15_data_o[5]), .S(n29730), .Q(n18016)
         );
  MUX21X1 U33318 ( .IN1(n34335), .IN2(s15_data_o[6]), .S(n29730), .Q(n18015)
         );
  MUX21X1 U33319 ( .IN1(n34521), .IN2(s15_data_o[7]), .S(n29730), .Q(n18014)
         );
  MUX21X1 U33320 ( .IN1(n34336), .IN2(s15_data_o[8]), .S(n29730), .Q(n18013)
         );
  MUX21X1 U33321 ( .IN1(n34483), .IN2(s15_data_o[9]), .S(n29730), .Q(n18012)
         );
  MUX21X1 U33322 ( .IN1(n34295), .IN2(s15_data_o[10]), .S(n29730), .Q(n18011)
         );
  MUX21X1 U33323 ( .IN1(n34556), .IN2(s15_data_o[11]), .S(n29730), .Q(n18010)
         );
  MUX21X1 U33324 ( .IN1(n34306), .IN2(s15_data_o[12]), .S(n29730), .Q(n18009)
         );
  MUX21X1 U33325 ( .IN1(n34522), .IN2(s15_data_o[13]), .S(n29730), .Q(n18008)
         );
  MUX21X1 U33326 ( .IN1(n34296), .IN2(s15_data_o[14]), .S(n29730), .Q(n18007)
         );
  MUX21X1 U33327 ( .IN1(n34559), .IN2(s15_data_o[15]), .S(n29730), .Q(n18006)
         );
  NOR2X0 U33328 ( .IN1(n29732), .IN2(n29731), .QN(n34072) );
  NAND2X0 U33329 ( .IN1(n29733), .IN2(n29789), .QN(n29779) );
  OA221X1 U33330 ( .IN1(n29791), .IN2(n29734), .IN3(n29791), .IN4(n29779), 
        .IN5(n29752), .Q(n29735) );
  OA21X1 U33331 ( .IN1(n29741), .IN2(n29736), .IN3(n29735), .Q(n29740) );
  NAND2X0 U33332 ( .IN1(\s1/msel/gnt_p3 [1]), .IN2(n29789), .QN(n29738) );
  OA222X1 U33333 ( .IN1(n29752), .IN2(n29791), .IN3(n29738), .IN4(
        \s1/msel/gnt_p3 [0]), .IN5(n29737), .IN6(\s1/msel/gnt_p3 [1]), .Q(
        n29739) );
  NOR3X0 U33334 ( .IN1(n34072), .IN2(n29740), .IN3(n29739), .QN(n29748) );
  NOR2X0 U33335 ( .IN1(\s1/msel/gnt_p3 [1]), .IN2(n29750), .QN(n29799) );
  NOR2X0 U33336 ( .IN1(n29742), .IN2(n29741), .QN(n34071) );
  NOR2X0 U33337 ( .IN1(n29799), .IN2(n34071), .QN(n29745) );
  NAND2X0 U33338 ( .IN1(n29765), .IN2(n29763), .QN(n29795) );
  NAND2X0 U33339 ( .IN1(n29756), .IN2(n29795), .QN(n29743) );
  NAND2X0 U33340 ( .IN1(n29752), .IN2(n29743), .QN(n29744) );
  NAND2X0 U33341 ( .IN1(n29745), .IN2(n29744), .QN(n29747) );
  NAND2X0 U33342 ( .IN1(\s1/msel/gnt_p3 [2]), .IN2(n29758), .QN(n29746) );
  OA22X1 U33343 ( .IN1(\s1/msel/gnt_p3 [2]), .IN2(n29748), .IN3(n29747), .IN4(
        n29746), .Q(n18005) );
  OA21X1 U33344 ( .IN1(n29765), .IN2(n29750), .IN3(n29749), .Q(n29766) );
  OA21X1 U33345 ( .IN1(n29773), .IN2(n29766), .IN3(n29751), .Q(n29774) );
  NOR3X0 U33346 ( .IN1(n29753), .IN2(n29774), .IN3(n29752), .QN(n29788) );
  NAND2X0 U33347 ( .IN1(n29790), .IN2(n29789), .QN(n29757) );
  NOR2X0 U33348 ( .IN1(n34280), .IN2(n29757), .QN(n29755) );
  NAND2X0 U33349 ( .IN1(n29792), .IN2(n29790), .QN(n29759) );
  NAND2X0 U33350 ( .IN1(n29758), .IN2(n29759), .QN(n29769) );
  AO221X1 U33351 ( .IN1(n29756), .IN2(n29755), .IN3(n29756), .IN4(n29769), 
        .IN5(n29754), .Q(n29775) );
  INVX0 U33352 ( .INP(n29756), .ZN(n29764) );
  NAND2X0 U33353 ( .IN1(\s1/msel/gnt_p3 [2]), .IN2(n29764), .QN(n29762) );
  AO221X1 U33354 ( .IN1(n29766), .IN2(n29765), .IN3(n29766), .IN4(n34280), 
        .IN5(n29757), .Q(n29760) );
  NAND4X0 U33355 ( .IN1(\s1/msel/gnt_p3 [2]), .IN2(n29760), .IN3(n29759), 
        .IN4(n29758), .QN(n29761) );
  AO22X1 U33356 ( .IN1(n29763), .IN2(n29775), .IN3(n29762), .IN4(n29761), .Q(
        n29787) );
  NOR2X0 U33357 ( .IN1(n29765), .IN2(n29764), .QN(n29770) );
  NAND3X0 U33358 ( .IN1(n29790), .IN2(\s1/msel/gnt_p3 [0]), .IN3(n29770), .QN(
        n29767) );
  NAND2X0 U33359 ( .IN1(n29767), .IN2(n29766), .QN(n29778) );
  OA221X1 U33360 ( .IN1(n29778), .IN2(n29770), .IN3(n29778), .IN4(n29769), 
        .IN5(n29768), .Q(n29786) );
  NAND2X0 U33361 ( .IN1(n29771), .IN2(n29770), .QN(n29780) );
  AO221X1 U33362 ( .IN1(n29774), .IN2(n29773), .IN3(n29774), .IN4(n29780), 
        .IN5(n29772), .Q(n29784) );
  NAND3X0 U33363 ( .IN1(n29777), .IN2(n29776), .IN3(n29775), .QN(n29783) );
  INVX0 U33364 ( .INP(n29778), .ZN(n29781) );
  AO21X1 U33365 ( .IN1(n29781), .IN2(n29780), .IN3(n29779), .Q(n29782) );
  NAND4X0 U33366 ( .IN1(n34428), .IN2(n29784), .IN3(n29783), .IN4(n29782), 
        .QN(n29785) );
  OA22X1 U33367 ( .IN1(n29788), .IN2(n29787), .IN3(n29786), .IN4(n29785), .Q(
        n29794) );
  OA221X1 U33368 ( .IN1(\s1/msel/gnt_p3 [1]), .IN2(n29790), .IN3(n34427), 
        .IN4(n29789), .IN5(n29794), .Q(n29804) );
  OA221X1 U33369 ( .IN1(\s1/msel/gnt_p3 [1]), .IN2(n29792), .IN3(n34427), 
        .IN4(n29791), .IN5(\s1/msel/gnt_p3 [0]), .Q(n29803) );
  NOR2X0 U33370 ( .IN1(n29793), .IN2(\s1/msel/gnt_p3 [0]), .QN(n29797) );
  NAND2X0 U33371 ( .IN1(n29795), .IN2(n29794), .QN(n29796) );
  NOR2X0 U33372 ( .IN1(n29797), .IN2(n29796), .QN(n29798) );
  AO221X1 U33373 ( .IN1(n29801), .IN2(n29800), .IN3(n29801), .IN4(n29799), 
        .IN5(n29798), .Q(n29802) );
  AO221X1 U33374 ( .IN1(n34428), .IN2(n29804), .IN3(n34428), .IN4(n29803), 
        .IN5(n29802), .Q(n18003) );
  NAND2X0 U33375 ( .IN1(n13472), .IN2(m7s1_cyc), .QN(n29887) );
  OR2X1 U33376 ( .IN1(n13528), .IN2(n29887), .Q(n29844) );
  NAND2X0 U33377 ( .IN1(n13606), .IN2(m5s1_cyc), .QN(n29888) );
  NOR2X0 U33378 ( .IN1(n13632), .IN2(n29888), .QN(n29850) );
  INVX0 U33379 ( .INP(n29850), .ZN(n29842) );
  NAND2X0 U33380 ( .IN1(\s1/msel/gnt_p1 [0]), .IN2(\s1/msel/gnt_p1 [2]), .QN(
        n29805) );
  AO221X1 U33381 ( .IN1(\s1/msel/gnt_p1 [1]), .IN2(n29844), .IN3(n34392), 
        .IN4(n29842), .IN5(n29805), .Q(n29885) );
  NAND2X0 U33382 ( .IN1(n13866), .IN2(m0s1_cyc), .QN(n29891) );
  NOR2X0 U33383 ( .IN1(n13898), .IN2(n29891), .QN(n29879) );
  NAND2X0 U33384 ( .IN1(n13814), .IN2(m1s1_cyc), .QN(n29890) );
  NOR2X0 U33385 ( .IN1(n13840), .IN2(n29890), .QN(n29877) );
  NOR2X0 U33386 ( .IN1(n29879), .IN2(n29877), .QN(n34074) );
  NAND2X0 U33387 ( .IN1(n13762), .IN2(m2s1_cyc), .QN(n29889) );
  NOR2X0 U33388 ( .IN1(n13788), .IN2(n29889), .QN(n29854) );
  NAND3X0 U33389 ( .IN1(n13710), .IN2(m3s1_cyc), .IN3(n34335), .QN(n29841) );
  INVX0 U33390 ( .INP(n29841), .ZN(n29866) );
  NOR2X0 U33391 ( .IN1(n29854), .IN2(n29866), .QN(n34076) );
  NAND3X0 U33392 ( .IN1(n13658), .IN2(m4s1_cyc), .IN3(n34336), .QN(n29857) );
  INVX0 U33393 ( .INP(n29857), .ZN(n29843) );
  NAND3X0 U33394 ( .IN1(n13554), .IN2(m6s1_cyc), .IN3(n34306), .QN(n29865) );
  INVX0 U33395 ( .INP(n29865), .ZN(n29834) );
  MUX21X1 U33396 ( .IN1(n29843), .IN2(n29834), .S(\s1/msel/gnt_p1 [1]), .Q(
        n29883) );
  AOI22X1 U33397 ( .IN1(n34074), .IN2(n34076), .IN3(n34673), .IN4(n29883), 
        .QN(n29807) );
  NOR2X0 U33398 ( .IN1(n29834), .IN2(n34673), .QN(n29862) );
  OA21X1 U33399 ( .IN1(\s1/msel/gnt_p1 [1]), .IN2(n29862), .IN3(n29844), .Q(
        n29820) );
  NAND2X0 U33400 ( .IN1(n29865), .IN2(n29844), .QN(n29818) );
  INVX0 U33401 ( .INP(n29818), .ZN(n34075) );
  AND2X1 U33402 ( .IN1(n29842), .IN2(n34075), .Q(n29806) );
  AO221X1 U33403 ( .IN1(n29807), .IN2(n29820), .IN3(n29807), .IN4(n29806), 
        .IN5(n34446), .Q(n29815) );
  NOR2X0 U33404 ( .IN1(n34673), .IN2(n34392), .QN(n29811) );
  NAND2X0 U33405 ( .IN1(n29866), .IN2(n29811), .QN(n29880) );
  NOR2X0 U33406 ( .IN1(\s1/msel/gnt_p1 [0]), .IN2(n34392), .QN(n29863) );
  NAND2X0 U33407 ( .IN1(n29854), .IN2(n29863), .QN(n29808) );
  AND3X1 U33408 ( .IN1(n34446), .IN2(n29880), .IN3(n29808), .Q(n29831) );
  INVX0 U33409 ( .INP(n29877), .ZN(n29847) );
  AND2X1 U33410 ( .IN1(n34392), .IN2(n29847), .Q(n29825) );
  AO22X1 U33411 ( .IN1(n34076), .IN2(n29825), .IN3(n29863), .IN4(n29841), .Q(
        n29810) );
  MUX21X1 U33412 ( .IN1(n29879), .IN2(n29877), .S(\s1/msel/gnt_p1 [0]), .Q(
        n29832) );
  INVX0 U33413 ( .INP(n29832), .ZN(n29809) );
  OA22X1 U33414 ( .IN1(n29811), .IN2(n29810), .IN3(\s1/msel/gnt_p1 [1]), .IN4(
        n29809), .Q(n29813) );
  NOR2X0 U33415 ( .IN1(n29850), .IN2(n29843), .QN(n34073) );
  NAND2X0 U33416 ( .IN1(n34075), .IN2(n34073), .QN(n29812) );
  NAND3X0 U33417 ( .IN1(n29831), .IN2(n29813), .IN3(n29812), .QN(n29814) );
  NAND3X0 U33418 ( .IN1(n29885), .IN2(n29815), .IN3(n29814), .QN(n18002) );
  NAND2X0 U33419 ( .IN1(n34673), .IN2(n34392), .QN(n29868) );
  INVX0 U33420 ( .INP(n29868), .ZN(n29822) );
  NAND2X0 U33421 ( .IN1(n34076), .IN2(n34075), .QN(n29816) );
  OR2X1 U33422 ( .IN1(n29818), .IN2(n34074), .Q(n29824) );
  NAND3X0 U33423 ( .IN1(n29842), .IN2(n29816), .IN3(n29824), .QN(n29821) );
  INVX0 U33424 ( .INP(n34076), .ZN(n29817) );
  AO221X1 U33425 ( .IN1(n34073), .IN2(\s1/msel/gnt_p1 [1]), .IN3(n34073), 
        .IN4(n29818), .IN5(n29817), .Q(n29826) );
  NAND2X0 U33426 ( .IN1(n34074), .IN2(n29826), .QN(n29819) );
  AO22X1 U33427 ( .IN1(n29822), .IN2(n29821), .IN3(n29820), .IN4(n29819), .Q(
        n29823) );
  NAND2X0 U33428 ( .IN1(\s1/msel/gnt_p1 [2]), .IN2(n29823), .QN(n29833) );
  NAND4X0 U33429 ( .IN1(\s1/msel/gnt_p1 [1]), .IN2(n29857), .IN3(n29842), 
        .IN4(n29824), .QN(n29829) );
  NAND2X0 U33430 ( .IN1(n29866), .IN2(n29863), .QN(n29828) );
  NAND2X0 U33431 ( .IN1(n29826), .IN2(n29825), .QN(n29827) );
  NAND4X0 U33432 ( .IN1(n34446), .IN2(n29829), .IN3(n29828), .IN4(n29827), 
        .QN(n29830) );
  NAND2X0 U33433 ( .IN1(n29833), .IN2(n29830), .QN(n29838) );
  OA21X1 U33434 ( .IN1(n29838), .IN2(n29832), .IN3(n29831), .Q(n29840) );
  INVX0 U33435 ( .INP(n29833), .ZN(n29837) );
  OA221X1 U33436 ( .IN1(\s1/msel/gnt_p1 [0]), .IN2(n29843), .IN3(n34673), 
        .IN4(n29850), .IN5(\s1/msel/gnt_p1 [2]), .Q(n29836) );
  NAND2X0 U33437 ( .IN1(\s1/msel/gnt_p1 [1]), .IN2(n29834), .QN(n29835) );
  OA22X1 U33438 ( .IN1(n29837), .IN2(n29836), .IN3(\s1/msel/gnt_p1 [0]), .IN4(
        n29835), .Q(n29839) );
  OAI22X1 U33439 ( .IN1(n29840), .IN2(n29839), .IN3(n34392), .IN4(n29838), 
        .QN(n18001) );
  NAND2X0 U33440 ( .IN1(n29865), .IN2(n29857), .QN(n29845) );
  OA21X1 U33441 ( .IN1(n29843), .IN2(n29842), .IN3(n29841), .Q(n29856) );
  OA21X1 U33442 ( .IN1(n34673), .IN2(n29845), .IN3(n29856), .Q(n29848) );
  AND2X1 U33443 ( .IN1(n29879), .IN2(n29856), .Q(n29846) );
  OA21X1 U33444 ( .IN1(n29847), .IN2(n29879), .IN3(n29844), .Q(n29858) );
  OA22X1 U33445 ( .IN1(n29848), .IN2(n29846), .IN3(n29858), .IN4(n29845), .Q(
        n29849) );
  OA21X1 U33446 ( .IN1(n29854), .IN2(n29848), .IN3(n29847), .Q(n29871) );
  OA22X1 U33447 ( .IN1(n29854), .IN2(n29849), .IN3(n29871), .IN4(n29868), .Q(
        n29853) );
  INVX0 U33448 ( .INP(n29858), .ZN(n29851) );
  AO21X1 U33449 ( .IN1(n29865), .IN2(n29851), .IN3(n29850), .Q(n29864) );
  NAND4X0 U33450 ( .IN1(\s1/msel/gnt_p1 [1]), .IN2(\s1/msel/gnt_p1 [0]), .IN3(
        n29864), .IN4(n29857), .QN(n29852) );
  NAND3X0 U33451 ( .IN1(n34446), .IN2(n29853), .IN3(n29852), .QN(n29876) );
  NOR2X0 U33452 ( .IN1(n29879), .IN2(n29854), .QN(n29867) );
  INVX0 U33453 ( .INP(n29867), .ZN(n29855) );
  NOR2X0 U33454 ( .IN1(n29856), .IN2(n29855), .QN(n29861) );
  NAND3X0 U33455 ( .IN1(\s1/msel/gnt_p1 [0]), .IN2(n29867), .IN3(n29857), .QN(
        n29859) );
  NAND2X0 U33456 ( .IN1(n29859), .IN2(n29858), .QN(n29860) );
  OAI22X1 U33457 ( .IN1(n29863), .IN2(n29862), .IN3(n29861), .IN4(n29860), 
        .QN(n29874) );
  INVX0 U33458 ( .INP(n29864), .ZN(n29870) );
  NAND3X0 U33459 ( .IN1(n29867), .IN2(n29866), .IN3(n29865), .QN(n29869) );
  AO21X1 U33460 ( .IN1(n29870), .IN2(n29869), .IN3(n29868), .Q(n29873) );
  OR3X1 U33461 ( .IN1(n34392), .IN2(n29879), .IN3(n29871), .Q(n29872) );
  NAND4X0 U33462 ( .IN1(\s1/msel/gnt_p1 [2]), .IN2(n29874), .IN3(n29873), 
        .IN4(n29872), .QN(n29875) );
  NAND2X0 U33463 ( .IN1(n29876), .IN2(n29875), .QN(n29882) );
  NAND2X0 U33464 ( .IN1(\s1/msel/gnt_p1 [0]), .IN2(n29877), .QN(n29878) );
  OA222X1 U33465 ( .IN1(n29882), .IN2(n29879), .IN3(n29882), .IN4(n34392), 
        .IN5(\s1/msel/gnt_p1 [1]), .IN6(n29878), .Q(n29881) );
  AO21X1 U33466 ( .IN1(n29881), .IN2(n29880), .IN3(\s1/msel/gnt_p1 [2]), .Q(
        n29886) );
  AO221X1 U33467 ( .IN1(n34673), .IN2(n34446), .IN3(n34673), .IN4(n29883), 
        .IN5(n29882), .Q(n29884) );
  NAND3X0 U33468 ( .IN1(n29886), .IN2(n29885), .IN3(n29884), .QN(n18000) );
  NAND3X0 U33469 ( .IN1(n13684), .IN2(n13658), .IN3(m4s1_cyc), .QN(n29934) );
  INVX0 U33470 ( .INP(n29934), .ZN(n29945) );
  NAND3X0 U33471 ( .IN1(n13580), .IN2(n13554), .IN3(m6s1_cyc), .QN(n29933) );
  INVX0 U33472 ( .INP(n29933), .ZN(n29947) );
  MUX21X1 U33473 ( .IN1(n29945), .IN2(n29947), .S(\s1/msel/gnt_p0 [1]), .Q(
        n29957) );
  NOR2X0 U33474 ( .IN1(n34296), .IN2(n29887), .QN(n29931) );
  INVX0 U33475 ( .INP(n29931), .ZN(n29940) );
  NAND2X0 U33476 ( .IN1(\s1/msel/gnt_p0 [1]), .IN2(n29940), .QN(n29958) );
  OR2X1 U33477 ( .IN1(n34295), .IN2(n29888), .Q(n29942) );
  NOR2X0 U33478 ( .IN1(n29947), .IN2(n29931), .QN(n29905) );
  NAND2X0 U33479 ( .IN1(n29942), .IN2(n29905), .QN(n29892) );
  NAND3X0 U33480 ( .IN1(n13736), .IN2(n13710), .IN3(m3s1_cyc), .QN(n29929) );
  INVX0 U33481 ( .INP(n29929), .ZN(n29895) );
  NOR2X0 U33482 ( .IN1(n34297), .IN2(n29889), .QN(n29944) );
  NOR2X0 U33483 ( .IN1(n29895), .IN2(n29944), .QN(n29902) );
  NOR2X0 U33484 ( .IN1(n34293), .IN2(n29890), .QN(n29930) );
  NOR2X0 U33485 ( .IN1(n34294), .IN2(n29891), .QN(n29949) );
  NOR2X0 U33486 ( .IN1(n29930), .IN2(n29949), .QN(n29909) );
  AO222X1 U33487 ( .IN1(n34233), .IN2(n29957), .IN3(n29958), .IN4(n29892), 
        .IN5(n29902), .IN6(n29909), .Q(n29901) );
  NAND3X0 U33488 ( .IN1(\s1/msel/gnt_p0 [0]), .IN2(\s1/msel/gnt_p0 [1]), .IN3(
        n29895), .QN(n29962) );
  NAND2X0 U33489 ( .IN1(\s1/msel/gnt_p0 [1]), .IN2(n34233), .QN(n29919) );
  INVX0 U33490 ( .INP(n29919), .ZN(n29893) );
  NAND2X0 U33491 ( .IN1(n29944), .IN2(n29893), .QN(n29894) );
  AND3X1 U33492 ( .IN1(n34454), .IN2(n29962), .IN3(n29894), .Q(n29917) );
  INVX0 U33493 ( .INP(n29905), .ZN(n29899) );
  NAND2X0 U33494 ( .IN1(n29934), .IN2(n29942), .QN(n29908) );
  INVX0 U33495 ( .INP(n29930), .ZN(n29941) );
  NAND2X0 U33496 ( .IN1(n34285), .IN2(n29941), .QN(n29903) );
  INVX0 U33497 ( .INP(n29902), .ZN(n29907) );
  OA22X1 U33498 ( .IN1(n29895), .IN2(n29919), .IN3(n29903), .IN4(n29907), .Q(
        n29897) );
  NAND2X0 U33499 ( .IN1(\s1/msel/gnt_p0 [0]), .IN2(\s1/msel/gnt_p0 [1]), .QN(
        n29896) );
  INVX0 U33500 ( .INP(n29949), .ZN(n29959) );
  NOR2X0 U33501 ( .IN1(\s1/msel/gnt_p0 [0]), .IN2(n29959), .QN(n29918) );
  AOI22X1 U33502 ( .IN1(n29897), .IN2(n29896), .IN3(n29918), .IN4(n34285), 
        .QN(n29898) );
  OA21X1 U33503 ( .IN1(n29899), .IN2(n29908), .IN3(n29898), .Q(n29900) );
  AO22X1 U33504 ( .IN1(\s1/msel/gnt_p0 [2]), .IN2(n29901), .IN3(n29917), .IN4(
        n29900), .Q(n17999) );
  OA21X1 U33505 ( .IN1(n29905), .IN2(n29908), .IN3(n29902), .Q(n29904) );
  OA22X1 U33506 ( .IN1(n29904), .IN2(n29903), .IN3(n29929), .IN4(n29919), .Q(
        n29916) );
  NAND3X0 U33507 ( .IN1(n29959), .IN2(\s1/msel/gnt_p0 [1]), .IN3(n29941), .QN(
        n29906) );
  NAND2X0 U33508 ( .IN1(n29906), .IN2(n29905), .QN(n29911) );
  NAND4X0 U33509 ( .IN1(\s1/msel/gnt_p0 [1]), .IN2(n29942), .IN3(n29934), 
        .IN4(n29911), .QN(n29915) );
  NAND2X0 U33510 ( .IN1(n29909), .IN2(n29907), .QN(n29914) );
  INVX0 U33511 ( .INP(n29908), .ZN(n29910) );
  AOI21X1 U33512 ( .IN1(n29910), .IN2(n29909), .IN3(n29958), .QN(n29913) );
  INVX0 U33513 ( .INP(n29911), .ZN(n29912) );
  AO221X1 U33514 ( .IN1(n29914), .IN2(n29913), .IN3(n29914), .IN4(n29912), 
        .IN5(n34454), .Q(n29920) );
  OA221X1 U33515 ( .IN1(\s1/msel/gnt_p0 [2]), .IN2(n29916), .IN3(
        \s1/msel/gnt_p0 [2]), .IN4(n29915), .IN5(n29920), .Q(n29928) );
  OA21X1 U33516 ( .IN1(n29928), .IN2(n29918), .IN3(n29917), .Q(n29927) );
  NOR2X0 U33517 ( .IN1(n29919), .IN2(n29933), .QN(n29925) );
  INVX0 U33518 ( .INP(n29920), .ZN(n29922) );
  NAND2X0 U33519 ( .IN1(n29945), .IN2(n34233), .QN(n29921) );
  NAND3X0 U33520 ( .IN1(n29922), .IN2(n29942), .IN3(n29921), .QN(n29923) );
  NAND2X0 U33521 ( .IN1(n29923), .IN2(\s1/msel/gnt_p0 [2]), .QN(n29924) );
  NOR2X0 U33522 ( .IN1(n29925), .IN2(n29924), .QN(n29926) );
  OAI22X1 U33523 ( .IN1(n29928), .IN2(n34285), .IN3(n29927), .IN4(n29926), 
        .QN(n17998) );
  OA21X1 U33524 ( .IN1(n29945), .IN2(n29942), .IN3(n29929), .Q(n29946) );
  OA21X1 U33525 ( .IN1(n29946), .IN2(n29944), .IN3(n29941), .Q(n29943) );
  OA21X1 U33526 ( .IN1(n29930), .IN2(\s1/msel/gnt_p0 [0]), .IN3(n29959), .Q(
        n29932) );
  NOR2X0 U33527 ( .IN1(n29932), .IN2(n29931), .QN(n29936) );
  NAND2X0 U33528 ( .IN1(n29934), .IN2(n29933), .QN(n29935) );
  NOR2X0 U33529 ( .IN1(n29936), .IN2(n29935), .QN(n29938) );
  INVX0 U33530 ( .INP(n29946), .ZN(n29937) );
  NOR2X0 U33531 ( .IN1(n29938), .IN2(n29937), .QN(n29939) );
  OA22X1 U33532 ( .IN1(\s1/msel/gnt_p0 [1]), .IN2(n29943), .IN3(n29944), .IN4(
        n29939), .Q(n29956) );
  OA21X1 U33533 ( .IN1(n29941), .IN2(n29949), .IN3(n29940), .Q(n29950) );
  OA21X1 U33534 ( .IN1(n29947), .IN2(n29950), .IN3(n29942), .Q(n29953) );
  OR4X1 U33535 ( .IN1(n34285), .IN2(n34233), .IN3(n29945), .IN4(n29953), .Q(
        n29955) );
  OR2X1 U33536 ( .IN1(n29943), .IN2(n29949), .Q(n29952) );
  AO221X1 U33537 ( .IN1(n29946), .IN2(n29945), .IN3(n29946), .IN4(n34233), 
        .IN5(n29944), .Q(n29948) );
  AO221X1 U33538 ( .IN1(n29950), .IN2(n29949), .IN3(n29950), .IN4(n29948), 
        .IN5(n29947), .Q(n29951) );
  OA221X1 U33539 ( .IN1(\s1/msel/gnt_p0 [1]), .IN2(n29953), .IN3(n34285), 
        .IN4(n29952), .IN5(n29951), .Q(n29954) );
  OA222X1 U33540 ( .IN1(\s1/msel/gnt_p0 [2]), .IN2(n29956), .IN3(
        \s1/msel/gnt_p0 [2]), .IN4(n29955), .IN5(n29954), .IN6(n34454), .Q(
        n29961) );
  AO221X1 U33541 ( .IN1(n34233), .IN2(n34454), .IN3(n34233), .IN4(n29957), 
        .IN5(n29961), .Q(n29967) );
  NAND4X0 U33542 ( .IN1(\s1/msel/gnt_p0 [2]), .IN2(\s1/msel/gnt_p0 [0]), .IN3(
        n29958), .IN4(\s1/msel/gnt_p0 [1]), .QN(n29966) );
  NOR2X0 U33543 ( .IN1(\s1/msel/gnt_p0 [1]), .IN2(n29959), .QN(n29960) );
  NOR2X0 U33544 ( .IN1(n29960), .IN2(\s1/msel/gnt_p0 [2]), .QN(n29964) );
  NAND2X0 U33545 ( .IN1(n29962), .IN2(n29961), .QN(n29963) );
  NAND2X0 U33546 ( .IN1(n29964), .IN2(n29963), .QN(n29965) );
  NAND3X0 U33547 ( .IN1(n29967), .IN2(n29966), .IN3(n29965), .QN(n17997) );
  NOR2X0 U33548 ( .IN1(n29979), .IN2(n29971), .QN(n29977) );
  NOR2X0 U33549 ( .IN1(n29971), .IN2(n29983), .QN(n29986) );
  OA22X1 U33550 ( .IN1(\s1/msel/gnt_p2 [1]), .IN2(n29969), .IN3(n29986), .IN4(
        n29968), .Q(n29976) );
  INVX0 U33551 ( .INP(n29970), .ZN(n29978) );
  OA21X1 U33552 ( .IN1(n29972), .IN2(n29971), .IN3(n29978), .Q(n29984) );
  INVX0 U33553 ( .INP(n29984), .ZN(n29973) );
  OA21X1 U33554 ( .IN1(n29977), .IN2(n29973), .IN3(n29996), .Q(n29975) );
  OA22X1 U33555 ( .IN1(n29977), .IN2(n29976), .IN3(n29975), .IN4(n29974), .Q(
        n29995) );
  OR2X1 U33556 ( .IN1(n29983), .IN2(n29978), .Q(n29987) );
  NAND2X0 U33557 ( .IN1(n29979), .IN2(n29987), .QN(n29982) );
  AO221X1 U33558 ( .IN1(n29982), .IN2(n29981), .IN3(n29982), .IN4(n29980), 
        .IN5(\s1/msel/gnt_p2 [2]), .Q(n29994) );
  NOR2X0 U33559 ( .IN1(n29984), .IN2(n29983), .QN(n29985) );
  NOR2X0 U33560 ( .IN1(n29985), .IN2(n34385), .QN(n29992) );
  INVX0 U33561 ( .INP(n29986), .ZN(n29988) );
  NAND3X0 U33562 ( .IN1(n29989), .IN2(n29988), .IN3(n29987), .QN(n29990) );
  NAND2X0 U33563 ( .IN1(\s1/msel/gnt_p2 [1]), .IN2(n29990), .QN(n29991) );
  NOR2X0 U33564 ( .IN1(n29992), .IN2(n29991), .QN(n29993) );
  OA22X1 U33565 ( .IN1(n29995), .IN2(n34437), .IN3(n29994), .IN4(n29993), .Q(
        n30007) );
  AND3X1 U33566 ( .IN1(\s1/msel/gnt_p2 [2]), .IN2(\s1/msel/gnt_p2 [0]), .IN3(
        n29996), .Q(n30006) );
  NAND2X0 U33567 ( .IN1(n29998), .IN2(n29997), .QN(n30001) );
  NAND3X0 U33568 ( .IN1(n30007), .IN2(n34385), .IN3(n29999), .QN(n30000) );
  NAND3X0 U33569 ( .IN1(n30001), .IN2(n30000), .IN3(\s1/msel/gnt_p2 [2]), .QN(
        n30002) );
  OA221X1 U33570 ( .IN1(n30004), .IN2(n30003), .IN3(n30004), .IN4(n30007), 
        .IN5(n30002), .Q(n30005) );
  AO221X1 U33571 ( .IN1(n30007), .IN2(\s1/msel/gnt_p2 [1]), .IN3(n30007), 
        .IN4(n30006), .IN5(n30005), .Q(n17995) );
  NOR2X0 U33572 ( .IN1(n30008), .IN2(n34379), .QN(n30009) );
  MUX21X1 U33573 ( .IN1(n34308), .IN2(s15_data_o[0]), .S(n30009), .Q(n17993)
         );
  MUX21X1 U33574 ( .IN1(n34523), .IN2(s15_data_o[1]), .S(n30009), .Q(n17992)
         );
  MUX21X1 U33575 ( .IN1(n34337), .IN2(s15_data_o[2]), .S(n30009), .Q(n17991)
         );
  MUX21X1 U33576 ( .IN1(n34524), .IN2(s15_data_o[3]), .S(n30009), .Q(n17990)
         );
  MUX21X1 U33577 ( .IN1(n34626), .IN2(s15_data_o[4]), .S(n30009), .Q(n17989)
         );
  MUX21X1 U33578 ( .IN1(n34563), .IN2(s15_data_o[5]), .S(n30009), .Q(n17988)
         );
  MUX21X1 U33579 ( .IN1(n34479), .IN2(s15_data_o[6]), .S(n30009), .Q(n17987)
         );
  MUX21X1 U33580 ( .IN1(n34647), .IN2(s15_data_o[7]), .S(n30009), .Q(n17986)
         );
  MUX21X1 U33581 ( .IN1(n34605), .IN2(s15_data_o[8]), .S(n30009), .Q(n17985)
         );
  MUX21X1 U33582 ( .IN1(n34373), .IN2(s15_data_o[9]), .S(n30009), .Q(n17984)
         );
  MUX21X1 U33583 ( .IN1(n34307), .IN2(s15_data_o[10]), .S(n30009), .Q(n17983)
         );
  MUX21X1 U33584 ( .IN1(n34484), .IN2(s15_data_o[11]), .S(n30009), .Q(n17982)
         );
  MUX21X1 U33585 ( .IN1(n34615), .IN2(s15_data_o[12]), .S(n30009), .Q(n17981)
         );
  MUX21X1 U33586 ( .IN1(n34576), .IN2(s15_data_o[13]), .S(n30009), .Q(n17980)
         );
  MUX21X1 U33587 ( .IN1(n34478), .IN2(s15_data_o[14]), .S(n30009), .Q(n17979)
         );
  MUX21X1 U33588 ( .IN1(n34641), .IN2(s15_data_o[15]), .S(n30009), .Q(n17978)
         );
  NOR2X0 U33589 ( .IN1(\s2/msel/gnt_p3 [0]), .IN2(n34395), .QN(n30056) );
  OA22X1 U33590 ( .IN1(n30051), .IN2(\s2/msel/gnt_p3 [0]), .IN3(n30024), .IN4(
        \s2/msel/gnt_p3 [1]), .Q(n30010) );
  NOR2X0 U33591 ( .IN1(n30056), .IN2(n30010), .QN(n30015) );
  INVX0 U33592 ( .INP(n30073), .ZN(n30086) );
  INVX0 U33593 ( .INP(n30051), .ZN(n30088) );
  MUX21X1 U33594 ( .IN1(n30086), .IN2(n30088), .S(\s2/msel/gnt_p3 [0]), .Q(
        n30047) );
  INVX0 U33595 ( .INP(n30087), .ZN(n30060) );
  NAND2X0 U33596 ( .IN1(\s2/msel/gnt_p3 [1]), .IN2(n30060), .QN(n30011) );
  NOR2X0 U33597 ( .IN1(n34277), .IN2(n34395), .QN(n30074) );
  INVX0 U33598 ( .INP(n30074), .ZN(n30064) );
  OAI221X1 U33599 ( .IN1(\s2/msel/gnt_p3 [1]), .IN2(n30047), .IN3(
        \s2/msel/gnt_p3 [0]), .IN4(n30011), .IN5(n30064), .QN(n30013) );
  INVX0 U33600 ( .INP(n30012), .ZN(n30072) );
  NAND2X0 U33601 ( .IN1(n30013), .IN2(n30072), .QN(n30014) );
  NOR2X0 U33602 ( .IN1(n30015), .IN2(n30014), .QN(n30021) );
  NOR2X0 U33603 ( .IN1(\s2/msel/gnt_p3 [0]), .IN2(\s2/msel/gnt_p3 [1]), .QN(
        n30026) );
  AO22X1 U33604 ( .IN1(n30056), .IN2(n30082), .IN3(n30070), .IN4(n30026), .Q(
        n30083) );
  INVX0 U33605 ( .INP(n30083), .ZN(n30018) );
  NAND2X0 U33606 ( .IN1(\s2/msel/gnt_p3 [1]), .IN2(n30055), .QN(n30043) );
  OA21X1 U33607 ( .IN1(\s2/msel/gnt_p3 [1]), .IN2(n30061), .IN3(n30043), .Q(
        n30085) );
  OR2X1 U33608 ( .IN1(\s2/msel/gnt_p3 [1]), .IN2(n30036), .Q(n30016) );
  NAND4X0 U33609 ( .IN1(n30018), .IN2(n30085), .IN3(n30017), .IN4(n30016), 
        .QN(n30019) );
  OA222X1 U33610 ( .IN1(\s2/msel/gnt_p3 [2]), .IN2(n30021), .IN3(
        \s2/msel/gnt_p3 [2]), .IN4(n30020), .IN5(n34548), .IN6(n30019), .Q(
        n17977) );
  NOR2X0 U33611 ( .IN1(\s2/msel/gnt_p3 [1]), .IN2(n34277), .QN(n30022) );
  NOR2X0 U33612 ( .IN1(n30056), .IN2(n30022), .QN(n30037) );
  NOR2X0 U33613 ( .IN1(n30024), .IN2(n30037), .QN(n30030) );
  NOR2X0 U33614 ( .IN1(\s2/msel/gnt_p3 [1]), .IN2(n30087), .QN(n30054) );
  OA21X1 U33615 ( .IN1(n30054), .IN2(n30023), .IN3(n30036), .Q(n30031) );
  INVX0 U33616 ( .INP(n30038), .ZN(n30025) );
  NOR2X0 U33617 ( .IN1(n30031), .IN2(n30025), .QN(n30027) );
  OAI21X1 U33618 ( .IN1(n34395), .IN2(n30025), .IN3(n30024), .QN(n30029) );
  INVX0 U33619 ( .INP(n30026), .ZN(n30075) );
  OA222X1 U33620 ( .IN1(n30027), .IN2(n30026), .IN3(n30027), .IN4(n30029), 
        .IN5(n30075), .IN6(n30051), .Q(n30028) );
  NOR2X0 U33621 ( .IN1(n30030), .IN2(n30028), .QN(n30042) );
  NOR2X0 U33622 ( .IN1(\s2/msel/gnt_p3 [0]), .IN2(n30044), .QN(n30071) );
  NAND2X0 U33623 ( .IN1(n30071), .IN2(n34395), .QN(n30034) );
  NAND2X0 U33624 ( .IN1(n30039), .IN2(n30029), .QN(n30033) );
  NOR2X0 U33625 ( .IN1(n30074), .IN2(n30030), .QN(n30032) );
  AO222X1 U33626 ( .IN1(n30034), .IN2(n30033), .IN3(n30034), .IN4(n30032), 
        .IN5(n30033), .IN6(n30031), .Q(n30035) );
  OA21X1 U33627 ( .IN1(n30037), .IN2(n30036), .IN3(n30035), .Q(n30041) );
  NAND3X0 U33628 ( .IN1(n30039), .IN2(n30056), .IN3(n30038), .QN(n30040) );
  OA221X1 U33629 ( .IN1(\s2/msel/gnt_p3 [2]), .IN2(n30042), .IN3(n34548), 
        .IN4(n30041), .IN5(n30040), .Q(n30050) );
  OR2X1 U33630 ( .IN1(n30070), .IN2(n30050), .Q(n30046) );
  OA21X1 U33631 ( .IN1(n30044), .IN2(n30050), .IN3(n30043), .Q(n30045) );
  OA221X1 U33632 ( .IN1(\s2/msel/gnt_p3 [0]), .IN2(n30046), .IN3(n34277), 
        .IN4(n30045), .IN5(\s2/msel/gnt_p3 [2]), .Q(n30049) );
  OA21X1 U33633 ( .IN1(n30064), .IN2(n30072), .IN3(n34548), .Q(n30091) );
  OA21X1 U33634 ( .IN1(n30050), .IN2(n30047), .IN3(n30091), .Q(n30048) );
  OAI22X1 U33635 ( .IN1(n30050), .IN2(n34395), .IN3(n30049), .IN4(n30048), 
        .QN(n17976) );
  OA21X1 U33636 ( .IN1(n30082), .IN2(n34277), .IN3(n30061), .Q(n30063) );
  OA21X1 U33637 ( .IN1(n30070), .IN2(n30063), .IN3(n30072), .Q(n30053) );
  OA21X1 U33638 ( .IN1(n30087), .IN2(n30053), .IN3(n30051), .Q(n30078) );
  AND3X1 U33639 ( .IN1(n30086), .IN2(n30061), .IN3(n30072), .Q(n30052) );
  NOR2X0 U33640 ( .IN1(n30053), .IN2(n30052), .QN(n30058) );
  NOR2X0 U33641 ( .IN1(n30070), .IN2(n30082), .QN(n30057) );
  OA221X1 U33642 ( .IN1(n30058), .IN2(n30055), .IN3(n30058), .IN4(n30057), 
        .IN5(n30054), .Q(n30067) );
  AO21X1 U33643 ( .IN1(n30088), .IN2(n30073), .IN3(n30055), .Q(n30059) );
  OA221X1 U33644 ( .IN1(n30058), .IN2(n30057), .IN3(n30058), .IN4(n30059), 
        .IN5(n30056), .Q(n30066) );
  INVX0 U33645 ( .INP(n30059), .ZN(n30081) );
  NAND2X0 U33646 ( .IN1(n30073), .IN2(n30060), .QN(n30069) );
  AND2X1 U33647 ( .IN1(n30061), .IN2(n30069), .Q(n30062) );
  OA22X1 U33648 ( .IN1(n30082), .IN2(n30081), .IN3(n30063), .IN4(n30062), .Q(
        n30076) );
  NOR3X0 U33649 ( .IN1(n30070), .IN2(n30076), .IN3(n30064), .QN(n30065) );
  NOR4X0 U33650 ( .IN1(\s2/msel/gnt_p3 [2]), .IN2(n30067), .IN3(n30066), .IN4(
        n30065), .QN(n30068) );
  OA21X1 U33651 ( .IN1(n30078), .IN2(n30075), .IN3(n30068), .Q(n30095) );
  AO221X1 U33652 ( .IN1(n30072), .IN2(n30071), .IN3(n30072), .IN4(n30070), 
        .IN5(n30069), .Q(n30080) );
  NAND2X0 U33653 ( .IN1(n30074), .IN2(n30073), .QN(n30077) );
  OA22X1 U33654 ( .IN1(n30078), .IN2(n30077), .IN3(n30076), .IN4(n30075), .Q(
        n30079) );
  OA221X1 U33655 ( .IN1(n30082), .IN2(n30081), .IN3(n30082), .IN4(n30080), 
        .IN5(n30079), .Q(n30084) );
  AO221X1 U33656 ( .IN1(\s2/msel/gnt_p3 [2]), .IN2(n30084), .IN3(n34548), 
        .IN4(n34277), .IN5(n30083), .Q(n30094) );
  OA21X1 U33657 ( .IN1(n30085), .IN2(n34277), .IN3(\s2/msel/gnt_p3 [2]), .Q(
        n30093) );
  AO221X1 U33658 ( .IN1(\s2/msel/gnt_p3 [1]), .IN2(n30087), .IN3(n34395), 
        .IN4(n30086), .IN5(n30095), .Q(n30090) );
  NAND3X0 U33659 ( .IN1(\s2/msel/gnt_p3 [0]), .IN2(n30088), .IN3(n34395), .QN(
        n30089) );
  AND3X1 U33660 ( .IN1(n30091), .IN2(n30090), .IN3(n30089), .Q(n30092) );
  OAI22X1 U33661 ( .IN1(n30095), .IN2(n30094), .IN3(n30093), .IN4(n30092), 
        .QN(n17975) );
  NAND3X0 U33662 ( .IN1(n13607), .IN2(m5s2_cyc), .IN3(n34307), .QN(n30134) );
  NAND2X0 U33663 ( .IN1(n34383), .IN2(n30134), .QN(n30159) );
  NAND3X0 U33664 ( .IN1(n13555), .IN2(m6s2_cyc), .IN3(n34615), .QN(n30121) );
  NAND3X0 U33665 ( .IN1(n13474), .IN2(m7s2_cyc), .IN3(n34478), .QN(n30132) );
  NAND2X0 U33666 ( .IN1(n30121), .IN2(n30132), .QN(n30101) );
  NAND2X0 U33667 ( .IN1(\s2/msel/gnt_p1 [1]), .IN2(n30132), .QN(n30158) );
  OA21X1 U33668 ( .IN1(n30159), .IN2(n30101), .IN3(n30158), .Q(n30096) );
  NAND3X0 U33669 ( .IN1(n13867), .IN2(m0s2_cyc), .IN3(n34308), .QN(n30131) );
  NAND3X0 U33670 ( .IN1(n13815), .IN2(m1s2_cyc), .IN3(n34337), .QN(n30133) );
  NAND2X0 U33671 ( .IN1(n30131), .IN2(n30133), .QN(n30109) );
  NAND3X0 U33672 ( .IN1(n13763), .IN2(m2s2_cyc), .IN3(n34626), .QN(n30130) );
  NAND3X0 U33673 ( .IN1(n13711), .IN2(m3s2_cyc), .IN3(n34479), .QN(n30129) );
  NAND2X0 U33674 ( .IN1(n30130), .IN2(n30129), .QN(n30113) );
  NOR2X0 U33675 ( .IN1(n30109), .IN2(n30113), .QN(n34085) );
  NOR2X0 U33676 ( .IN1(n30096), .IN2(n34085), .QN(n30098) );
  NAND3X0 U33677 ( .IN1(n13659), .IN2(m4s2_cyc), .IN3(n34605), .QN(n30112) );
  INVX0 U33678 ( .INP(n30112), .ZN(n30143) );
  INVX0 U33679 ( .INP(n30121), .ZN(n30148) );
  MUX21X1 U33680 ( .IN1(n30143), .IN2(n30148), .S(\s2/msel/gnt_p1 [1]), .Q(
        n30161) );
  NAND2X0 U33681 ( .IN1(n34241), .IN2(n30161), .QN(n30097) );
  NAND2X0 U33682 ( .IN1(n30098), .IN2(n30097), .QN(n30105) );
  OA21X1 U33683 ( .IN1(\s2/msel/gnt_p1 [0]), .IN2(n30131), .IN3(n30133), .Q(
        n30120) );
  NOR2X0 U33684 ( .IN1(n34241), .IN2(n34383), .QN(n30100) );
  INVX0 U33685 ( .INP(n30113), .ZN(n30099) );
  OA22X1 U33686 ( .IN1(\s2/msel/gnt_p1 [1]), .IN2(n30120), .IN3(n30100), .IN4(
        n30099), .Q(n30104) );
  AND2X1 U33687 ( .IN1(n30134), .IN2(n30112), .Q(n30107) );
  INVX0 U33688 ( .INP(n30101), .ZN(n30110) );
  AND2X1 U33689 ( .IN1(n30107), .IN2(n30110), .Q(n34086) );
  AO221X1 U33690 ( .IN1(\s2/msel/gnt_p1 [0]), .IN2(n30129), .IN3(n34241), 
        .IN4(n30130), .IN5(n34383), .Q(n30102) );
  NAND2X0 U33691 ( .IN1(n30102), .IN2(n34438), .QN(n30118) );
  NOR2X0 U33692 ( .IN1(n34086), .IN2(n30118), .QN(n30103) );
  AO22X1 U33693 ( .IN1(\s2/msel/gnt_p1 [2]), .IN2(n30105), .IN3(n30104), .IN4(
        n30103), .Q(n17974) );
  INVX0 U33694 ( .INP(n30109), .ZN(n30106) );
  OA21X1 U33695 ( .IN1(n30107), .IN2(n30113), .IN3(n30106), .Q(n30108) );
  NAND2X0 U33696 ( .IN1(n30110), .IN2(n34383), .QN(n30111) );
  OA22X1 U33697 ( .IN1(n30108), .IN2(n30158), .IN3(n30113), .IN4(n30111), .Q(
        n30117) );
  NAND2X0 U33698 ( .IN1(n30110), .IN2(n30109), .QN(n30116) );
  NAND4X0 U33699 ( .IN1(n30134), .IN2(n30112), .IN3(n30116), .IN4(n30111), 
        .QN(n30115) );
  NAND2X0 U33700 ( .IN1(n34383), .IN2(n30113), .QN(n30114) );
  NAND4X0 U33701 ( .IN1(n34438), .IN2(n30129), .IN3(n30115), .IN4(n30114), 
        .QN(n30119) );
  OA221X1 U33702 ( .IN1(n34438), .IN2(n30117), .IN3(n34438), .IN4(n30116), 
        .IN5(n30119), .Q(n30128) );
  AO21X1 U33703 ( .IN1(n30120), .IN2(n30119), .IN3(n30118), .Q(n30127) );
  NOR2X0 U33704 ( .IN1(n34383), .IN2(n30121), .QN(n30122) );
  NAND2X0 U33705 ( .IN1(n30122), .IN2(n34241), .QN(n30125) );
  NAND2X0 U33706 ( .IN1(n30143), .IN2(n34241), .QN(n30123) );
  NAND3X0 U33707 ( .IN1(n30123), .IN2(n30134), .IN3(n30128), .QN(n30124) );
  NAND3X0 U33708 ( .IN1(n30125), .IN2(n30124), .IN3(\s2/msel/gnt_p1 [2]), .QN(
        n30126) );
  AO22X1 U33709 ( .IN1(\s2/msel/gnt_p1 [1]), .IN2(n30128), .IN3(n30127), .IN4(
        n30126), .Q(n17973) );
  NOR2X0 U33710 ( .IN1(\s2/msel/gnt_p1 [1]), .IN2(n30131), .QN(n30156) );
  INVX0 U33711 ( .INP(n30130), .ZN(n30146) );
  OA21X1 U33712 ( .IN1(n30143), .IN2(n30134), .IN3(n30129), .Q(n30149) );
  OAI21X1 U33713 ( .IN1(n30146), .IN2(n30149), .IN3(n30133), .QN(n30150) );
  NAND3X0 U33714 ( .IN1(\s2/msel/gnt_p1 [1]), .IN2(n30150), .IN3(n30131), .QN(
        n30141) );
  NAND2X0 U33715 ( .IN1(n30131), .IN2(n30130), .QN(n30135) );
  INVX0 U33716 ( .INP(n30131), .ZN(n30144) );
  OA21X1 U33717 ( .IN1(n30144), .IN2(n30133), .IN3(n30132), .Q(n30145) );
  OA21X1 U33718 ( .IN1(n34241), .IN2(n30135), .IN3(n30145), .Q(n30137) );
  OA21X1 U33719 ( .IN1(n30148), .IN2(n30137), .IN3(n30134), .Q(n30142) );
  NAND2X0 U33720 ( .IN1(n34241), .IN2(n34383), .QN(n30139) );
  AND2X1 U33721 ( .IN1(n30145), .IN2(n30143), .Q(n30136) );
  OA22X1 U33722 ( .IN1(n30137), .IN2(n30136), .IN3(n30149), .IN4(n30135), .Q(
        n30138) );
  OA22X1 U33723 ( .IN1(n30142), .IN2(n30139), .IN3(n30148), .IN4(n30138), .Q(
        n30140) );
  NAND3X0 U33724 ( .IN1(n30141), .IN2(n30140), .IN3(\s2/msel/gnt_p1 [2]), .QN(
        n30155) );
  OR4X1 U33725 ( .IN1(n34383), .IN2(n34241), .IN3(n30142), .IN4(n30143), .Q(
        n30153) );
  AO221X1 U33726 ( .IN1(n30145), .IN2(n30144), .IN3(n30145), .IN4(n34241), 
        .IN5(n30143), .Q(n30147) );
  AO221X1 U33727 ( .IN1(n30149), .IN2(n30148), .IN3(n30149), .IN4(n30147), 
        .IN5(n30146), .Q(n30152) );
  NAND2X0 U33728 ( .IN1(n30150), .IN2(n34383), .QN(n30151) );
  NAND4X0 U33729 ( .IN1(n34438), .IN2(n30153), .IN3(n30152), .IN4(n30151), 
        .QN(n30154) );
  NAND2X0 U33730 ( .IN1(n30155), .IN2(n30154), .QN(n30160) );
  AO221X1 U33731 ( .IN1(n30157), .IN2(n30156), .IN3(n30157), .IN4(n30160), 
        .IN5(\s2/msel/gnt_p1 [2]), .Q(n30164) );
  NAND4X0 U33732 ( .IN1(\s2/msel/gnt_p1 [2]), .IN2(\s2/msel/gnt_p1 [0]), .IN3(
        n30159), .IN4(n30158), .QN(n30163) );
  AO221X1 U33733 ( .IN1(n34241), .IN2(n34438), .IN3(n34241), .IN4(n30161), 
        .IN5(n30160), .Q(n30162) );
  NAND3X0 U33734 ( .IN1(n30164), .IN2(n30163), .IN3(n30162), .QN(n17972) );
  NAND3X0 U33735 ( .IN1(n13633), .IN2(n13607), .IN3(m5s2_cyc), .QN(n30219) );
  NAND3X0 U33736 ( .IN1(n13529), .IN2(n13474), .IN3(m7s2_cyc), .QN(n30215) );
  MUX21X1 U33737 ( .IN1(n30219), .IN2(n30215), .S(\s2/msel/gnt_p0 [1]), .Q(
        n30234) );
  NAND3X0 U33738 ( .IN1(n13581), .IN2(n13555), .IN3(m6s2_cyc), .QN(n30212) );
  NAND2X0 U33739 ( .IN1(n30212), .IN2(n30215), .QN(n30177) );
  NAND2X0 U33740 ( .IN1(n34670), .IN2(n30177), .QN(n30167) );
  NAND3X0 U33741 ( .IN1(n13685), .IN2(n13659), .IN3(m4s2_cyc), .QN(n30211) );
  INVX0 U33742 ( .INP(n30211), .ZN(n30222) );
  INVX0 U33743 ( .INP(n30212), .ZN(n30218) );
  MUX21X1 U33744 ( .IN1(n30222), .IN2(n30218), .S(\s2/msel/gnt_p0 [1]), .Q(
        n30232) );
  NAND2X0 U33745 ( .IN1(n34554), .IN2(n30232), .QN(n30166) );
  NAND3X0 U33746 ( .IN1(n13789), .IN2(n13763), .IN3(m2s2_cyc), .QN(n30200) );
  NAND3X0 U33747 ( .IN1(n13900), .IN2(n13867), .IN3(m0s2_cyc), .QN(n30203) );
  NAND3X0 U33748 ( .IN1(n13737), .IN2(n13711), .IN3(m3s2_cyc), .QN(n30202) );
  NAND3X0 U33749 ( .IN1(n13841), .IN2(n13815), .IN3(m1s2_cyc), .QN(n30209) );
  NAND4X0 U33750 ( .IN1(n30200), .IN2(n30203), .IN3(n30202), .IN4(n30209), 
        .QN(n30165) );
  NAND4X0 U33751 ( .IN1(n30234), .IN2(n30167), .IN3(n30166), .IN4(n30165), 
        .QN(n30174) );
  NAND2X0 U33752 ( .IN1(\s2/msel/gnt_p0 [0]), .IN2(\s2/msel/gnt_p0 [1]), .QN(
        n30216) );
  INVX0 U33753 ( .INP(n30216), .ZN(n30169) );
  INVX0 U33754 ( .INP(n30200), .ZN(n30226) );
  INVX0 U33755 ( .INP(n30202), .ZN(n30208) );
  NOR2X0 U33756 ( .IN1(n30226), .IN2(n30208), .QN(n30176) );
  NOR2X0 U33757 ( .IN1(\s2/msel/gnt_p0 [0]), .IN2(n34670), .QN(n30193) );
  AO22X1 U33758 ( .IN1(n30209), .IN2(n30176), .IN3(n30193), .IN4(n30202), .Q(
        n30168) );
  NAND2X0 U33759 ( .IN1(n30211), .IN2(n30219), .QN(n30175) );
  OA22X1 U33760 ( .IN1(n30169), .IN2(n30168), .IN3(n30175), .IN4(n30177), .Q(
        n30173) );
  NOR3X0 U33761 ( .IN1(\s2/msel/gnt_p0 [1]), .IN2(\s2/msel/gnt_p0 [0]), .IN3(
        n30203), .QN(n30171) );
  NAND2X0 U33762 ( .IN1(n30193), .IN2(n30226), .QN(n30170) );
  NAND2X0 U33763 ( .IN1(n30208), .IN2(n30169), .QN(n30230) );
  NAND3X0 U33764 ( .IN1(n30170), .IN2(n30230), .IN3(n34291), .QN(n30192) );
  NOR2X0 U33765 ( .IN1(n30171), .IN2(n30192), .QN(n30172) );
  AO22X1 U33766 ( .IN1(\s2/msel/gnt_p0 [2]), .IN2(n30174), .IN3(n30173), .IN4(
        n30172), .Q(n17971) );
  NAND2X0 U33767 ( .IN1(n30193), .IN2(n30208), .QN(n30182) );
  NAND4X0 U33768 ( .IN1(n30200), .IN2(n30212), .IN3(n30202), .IN4(n30215), 
        .QN(n30183) );
  NAND2X0 U33769 ( .IN1(n30176), .IN2(n30175), .QN(n30184) );
  NAND4X0 U33770 ( .IN1(n34670), .IN2(n30209), .IN3(n30183), .IN4(n30184), 
        .QN(n30181) );
  INVX0 U33771 ( .INP(n30177), .ZN(n30179) );
  NAND2X0 U33772 ( .IN1(n30203), .IN2(n30209), .QN(n30178) );
  NAND2X0 U33773 ( .IN1(n30179), .IN2(n30178), .QN(n30186) );
  NAND4X0 U33774 ( .IN1(\s2/msel/gnt_p0 [1]), .IN2(n30219), .IN3(n30211), 
        .IN4(n30186), .QN(n30180) );
  NAND3X0 U33775 ( .IN1(n30182), .IN2(n30181), .IN3(n30180), .QN(n30191) );
  NOR2X0 U33776 ( .IN1(n30183), .IN2(\s2/msel/gnt_p0 [1]), .QN(n30189) );
  NAND3X0 U33777 ( .IN1(n30203), .IN2(n30209), .IN3(n30184), .QN(n30185) );
  NAND3X0 U33778 ( .IN1(\s2/msel/gnt_p0 [1]), .IN2(n30215), .IN3(n30185), .QN(
        n30187) );
  NAND2X0 U33779 ( .IN1(n30187), .IN2(n30186), .QN(n30188) );
  NOR2X0 U33780 ( .IN1(n30189), .IN2(n30188), .QN(n30190) );
  MUX21X1 U33781 ( .IN1(n30191), .IN2(n30190), .S(\s2/msel/gnt_p0 [2]), .Q(
        n30199) );
  AO221X1 U33782 ( .IN1(n30199), .IN2(\s2/msel/gnt_p0 [0]), .IN3(n30199), 
        .IN4(n30203), .IN5(n30192), .Q(n30198) );
  NAND2X0 U33783 ( .IN1(n30193), .IN2(n30218), .QN(n30196) );
  NAND2X0 U33784 ( .IN1(n30222), .IN2(n34554), .QN(n30194) );
  NAND3X0 U33785 ( .IN1(n30194), .IN2(n30199), .IN3(n30219), .QN(n30195) );
  NAND3X0 U33786 ( .IN1(n30196), .IN2(n30195), .IN3(\s2/msel/gnt_p0 [2]), .QN(
        n30197) );
  AO22X1 U33787 ( .IN1(\s2/msel/gnt_p0 [1]), .IN2(n30199), .IN3(n30198), .IN4(
        n30197), .Q(n17970) );
  NOR2X0 U33788 ( .IN1(n30222), .IN2(n30219), .QN(n30207) );
  NAND3X0 U33789 ( .IN1(n30207), .IN2(n30200), .IN3(n30203), .QN(n30205) );
  NAND2X0 U33790 ( .IN1(n30200), .IN2(n30203), .QN(n30201) );
  AO221X1 U33791 ( .IN1(n30202), .IN2(n30222), .IN3(n30202), .IN4(n34554), 
        .IN5(n30201), .Q(n30204) );
  INVX0 U33792 ( .INP(n30203), .ZN(n30231) );
  OA21X1 U33793 ( .IN1(n30231), .IN2(n30209), .IN3(n30215), .Q(n30217) );
  NAND3X0 U33794 ( .IN1(n30205), .IN2(n30204), .IN3(n30217), .QN(n30206) );
  NAND2X0 U33795 ( .IN1(n30206), .IN2(n30212), .QN(n30229) );
  NOR2X0 U33796 ( .IN1(n30208), .IN2(n30207), .QN(n30225) );
  OA21X1 U33797 ( .IN1(n30226), .IN2(n30225), .IN3(n30209), .Q(n30220) );
  OR3X1 U33798 ( .IN1(n34670), .IN2(n30231), .IN3(n30220), .Q(n30228) );
  INVX0 U33799 ( .INP(n30209), .ZN(n30210) );
  NOR2X0 U33800 ( .IN1(\s2/msel/gnt_p0 [0]), .IN2(n30210), .QN(n30214) );
  NAND2X0 U33801 ( .IN1(n30212), .IN2(n30211), .QN(n30213) );
  AO221X1 U33802 ( .IN1(n30215), .IN2(n30231), .IN3(n30215), .IN4(n30214), 
        .IN5(n30213), .Q(n30224) );
  AO221X1 U33803 ( .IN1(n30219), .IN2(n30218), .IN3(n30219), .IN4(n30217), 
        .IN5(n30216), .Q(n30221) );
  OA22X1 U33804 ( .IN1(n30222), .IN2(n30221), .IN3(\s2/msel/gnt_p0 [1]), .IN4(
        n30220), .Q(n30223) );
  OA221X1 U33805 ( .IN1(n30226), .IN2(n30225), .IN3(n30226), .IN4(n30224), 
        .IN5(n30223), .Q(n30227) );
  OA222X1 U33806 ( .IN1(n34291), .IN2(n30229), .IN3(n34291), .IN4(n30228), 
        .IN5(n30227), .IN6(\s2/msel/gnt_p0 [2]), .Q(n30233) );
  OA221X1 U33807 ( .IN1(n30233), .IN2(n30231), .IN3(n30233), .IN4(n34670), 
        .IN5(n30230), .Q(n30237) );
  OA21X1 U33808 ( .IN1(n34291), .IN2(n30232), .IN3(n34554), .Q(n30236) );
  OA21X1 U33809 ( .IN1(n34291), .IN2(n30234), .IN3(n30233), .Q(n30235) );
  OAI22X1 U33810 ( .IN1(\s2/msel/gnt_p0 [2]), .IN2(n30237), .IN3(n30236), 
        .IN4(n30235), .QN(n17969) );
  NAND2X0 U33811 ( .IN1(\s2/msel/gnt_p2 [1]), .IN2(n30283), .QN(n30321) );
  NAND2X0 U33812 ( .IN1(n34268), .IN2(n30289), .QN(n30322) );
  MUX21X1 U33813 ( .IN1(n30296), .IN2(n30312), .S(\s2/msel/gnt_p2 [1]), .Q(
        n30325) );
  NOR2X0 U33814 ( .IN1(\s2/msel/gnt_p2 [0]), .IN2(n30325), .QN(n30238) );
  AO221X1 U33815 ( .IN1(n30321), .IN2(n30322), .IN3(n30321), .IN4(n30251), 
        .IN5(n30238), .Q(n30245) );
  INVX0 U33816 ( .INP(n30284), .ZN(n30239) );
  NAND2X0 U33817 ( .IN1(\s2/msel/gnt_p2 [0]), .IN2(n30239), .QN(n30317) );
  OA21X1 U33818 ( .IN1(\s2/msel/gnt_p2 [0]), .IN2(n30297), .IN3(n30317), .Q(
        n30270) );
  NOR2X0 U33819 ( .IN1(\s2/msel/gnt_p2 [1]), .IN2(n30270), .QN(n30243) );
  NAND2X0 U33820 ( .IN1(\s2/msel/gnt_p2 [0]), .IN2(n34268), .QN(n30256) );
  NAND2X0 U33821 ( .IN1(n34609), .IN2(n34268), .QN(n30301) );
  OR2X1 U33822 ( .IN1(n30239), .IN2(n30301), .Q(n30255) );
  AND2X1 U33823 ( .IN1(n30256), .IN2(n30255), .Q(n30240) );
  OA22X1 U33824 ( .IN1(n30260), .IN2(n34268), .IN3(n30240), .IN4(n30254), .Q(
        n30242) );
  NAND2X0 U33825 ( .IN1(\s2/msel/gnt_p2 [1]), .IN2(n34609), .QN(n30263) );
  INVX0 U33826 ( .INP(n30263), .ZN(n30274) );
  INVX0 U33827 ( .INP(n30314), .ZN(n30288) );
  NAND2X0 U33828 ( .IN1(n30274), .IN2(n30288), .QN(n30241) );
  NAND3X0 U33829 ( .IN1(\s2/msel/gnt_p2 [0]), .IN2(\s2/msel/gnt_p2 [1]), .IN3(
        n30260), .QN(n30320) );
  NAND3X0 U33830 ( .IN1(n30241), .IN2(n30320), .IN3(n34391), .QN(n30268) );
  NOR4X0 U33831 ( .IN1(n30243), .IN2(n34088), .IN3(n30242), .IN4(n30268), .QN(
        n30244) );
  AO221X1 U33832 ( .IN1(\s2/msel/gnt_p2 [2]), .IN2(n34089), .IN3(
        \s2/msel/gnt_p2 [2]), .IN4(n30245), .IN5(n30244), .Q(n17968) );
  INVX0 U33833 ( .INP(n30247), .ZN(n30246) );
  AND2X1 U33834 ( .IN1(n30254), .IN2(n30246), .Q(n30250) );
  NAND2X0 U33835 ( .IN1(n34268), .IN2(n30314), .QN(n30295) );
  OA221X1 U33836 ( .IN1(n30251), .IN2(n30246), .IN3(n30251), .IN4(n30295), 
        .IN5(n30289), .Q(n30261) );
  OR2X1 U33837 ( .IN1(n30261), .IN2(n30301), .Q(n30249) );
  NOR2X0 U33838 ( .IN1(n30247), .IN2(n30252), .QN(n30259) );
  OA22X1 U33839 ( .IN1(n30259), .IN2(n30321), .IN3(n30251), .IN4(n30256), .Q(
        n30248) );
  AO222X1 U33840 ( .IN1(n30250), .IN2(n30249), .IN3(n30250), .IN4(n30289), 
        .IN5(n30249), .IN6(n30248), .Q(n30267) );
  INVX0 U33841 ( .INP(n30251), .ZN(n30253) );
  NOR2X0 U33842 ( .IN1(n30253), .IN2(n30252), .QN(n30258) );
  NOR2X0 U33843 ( .IN1(n30258), .IN2(n30254), .QN(n30257) );
  OA221X1 U33844 ( .IN1(n30257), .IN2(n30256), .IN3(n30257), .IN4(n30255), 
        .IN5(n34391), .Q(n30266) );
  NOR3X0 U33845 ( .IN1(n30260), .IN2(n30259), .IN3(n30258), .QN(n30264) );
  NAND2X0 U33846 ( .IN1(n30296), .IN2(\s2/msel/gnt_p2 [0]), .QN(n30285) );
  OR2X1 U33847 ( .IN1(n34268), .IN2(n30285), .Q(n30292) );
  INVX0 U33848 ( .INP(n30261), .ZN(n30262) );
  OA22X1 U33849 ( .IN1(n30264), .IN2(n30263), .IN3(n30292), .IN4(n30262), .Q(
        n30265) );
  NAND2X0 U33850 ( .IN1(n30266), .IN2(n30265), .QN(n30269) );
  OA21X1 U33851 ( .IN1(n30267), .IN2(n34391), .IN3(n30269), .Q(n30279) );
  AO21X1 U33852 ( .IN1(n30270), .IN2(n30269), .IN3(n30268), .Q(n30278) );
  INVX0 U33853 ( .INP(n30296), .ZN(n30281) );
  NOR2X0 U33854 ( .IN1(\s2/msel/gnt_p2 [0]), .IN2(n30281), .QN(n30306) );
  NOR2X0 U33855 ( .IN1(\s2/msel/gnt_p2 [0]), .IN2(n30306), .QN(n30272) );
  NAND2X0 U33856 ( .IN1(n30279), .IN2(n30289), .QN(n30271) );
  NOR2X0 U33857 ( .IN1(n30272), .IN2(n30271), .QN(n30273) );
  NOR2X0 U33858 ( .IN1(n30273), .IN2(n34391), .QN(n30276) );
  INVX0 U33859 ( .INP(n30312), .ZN(n30291) );
  NAND2X0 U33860 ( .IN1(n30291), .IN2(n30274), .QN(n30275) );
  NAND2X0 U33861 ( .IN1(n30276), .IN2(n30275), .QN(n30277) );
  AO22X1 U33862 ( .IN1(\s2/msel/gnt_p2 [1]), .IN2(n30279), .IN3(n30278), .IN4(
        n30277), .Q(n17967) );
  INVX0 U33863 ( .INP(n30297), .ZN(n30316) );
  OA21X1 U33864 ( .IN1(n30289), .IN2(n30281), .IN3(n30280), .Q(n30300) );
  OA21X1 U33865 ( .IN1(n30288), .IN2(n30300), .IN3(n30284), .Q(n30287) );
  OR3X1 U33866 ( .IN1(n34268), .IN2(n30316), .IN3(n30287), .Q(n30282) );
  NAND2X0 U33867 ( .IN1(\s2/msel/gnt_p2 [2]), .IN2(n30282), .QN(n30313) );
  NAND2X0 U33868 ( .IN1(n30314), .IN2(n30297), .QN(n30290) );
  OA21X1 U33869 ( .IN1(n30284), .IN2(n30316), .IN3(n30283), .Q(n30304) );
  OAI221X1 U33870 ( .IN1(n30290), .IN2(n30285), .IN3(n30290), .IN4(n30300), 
        .IN5(n30304), .QN(n30311) );
  NAND3X0 U33871 ( .IN1(n30286), .IN2(n30312), .IN3(n30296), .QN(n30299) );
  OA21X1 U33872 ( .IN1(n30288), .IN2(n30299), .IN3(n30287), .Q(n30294) );
  OA221X1 U33873 ( .IN1(n30291), .IN2(n30304), .IN3(n30291), .IN4(n30290), 
        .IN5(n30289), .Q(n30293) );
  OA22X1 U33874 ( .IN1(n30294), .IN2(n30301), .IN3(n30293), .IN4(n30292), .Q(
        n30309) );
  NAND2X0 U33875 ( .IN1(\s2/msel/gnt_p2 [0]), .IN2(n30295), .QN(n30303) );
  NAND4X0 U33876 ( .IN1(\s2/msel/gnt_p2 [0]), .IN2(n30297), .IN3(n30312), 
        .IN4(n30296), .QN(n30298) );
  NAND3X0 U33877 ( .IN1(n30300), .IN2(n30299), .IN3(n30298), .QN(n30302) );
  NAND3X0 U33878 ( .IN1(n30303), .IN2(n30302), .IN3(n30301), .QN(n30308) );
  INVX0 U33879 ( .INP(n30304), .ZN(n30305) );
  NAND4X0 U33880 ( .IN1(\s2/msel/gnt_p2 [1]), .IN2(n30306), .IN3(n30305), 
        .IN4(n30312), .QN(n30307) );
  NAND4X0 U33881 ( .IN1(n30309), .IN2(n34391), .IN3(n30308), .IN4(n30307), 
        .QN(n30310) );
  OA221X1 U33882 ( .IN1(n30313), .IN2(n30312), .IN3(n30313), .IN4(n30311), 
        .IN5(n30310), .Q(n30315) );
  NAND3X0 U33883 ( .IN1(\s2/msel/gnt_p2 [1]), .IN2(n30315), .IN3(n30314), .QN(
        n30319) );
  INVX0 U33884 ( .INP(n30315), .ZN(n30323) );
  AO221X1 U33885 ( .IN1(n30317), .IN2(n30316), .IN3(n30317), .IN4(n30323), 
        .IN5(\s2/msel/gnt_p2 [1]), .Q(n30318) );
  NAND3X0 U33886 ( .IN1(n30320), .IN2(n30319), .IN3(n30318), .QN(n30328) );
  NAND3X0 U33887 ( .IN1(n30322), .IN2(\s2/msel/gnt_p2 [2]), .IN3(n30321), .QN(
        n30324) );
  NAND2X0 U33888 ( .IN1(n30324), .IN2(n30323), .QN(n30327) );
  AO21X1 U33889 ( .IN1(\s2/msel/gnt_p2 [2]), .IN2(n30325), .IN3(
        \s2/msel/gnt_p2 [0]), .Q(n30326) );
  AO22X1 U33890 ( .IN1(n34391), .IN2(n30328), .IN3(n30327), .IN4(n30326), .Q(
        n17966) );
  NOR2X0 U33891 ( .IN1(n30329), .IN2(n34379), .QN(n30330) );
  MUX21X1 U33892 ( .IN1(n34309), .IN2(s15_data_o[0]), .S(n30330), .Q(n17965)
         );
  MUX21X1 U33893 ( .IN1(n34485), .IN2(s15_data_o[1]), .S(n30330), .Q(n17964)
         );
  MUX21X1 U33894 ( .IN1(n34310), .IN2(s15_data_o[2]), .S(n30330), .Q(n17963)
         );
  MUX21X1 U33895 ( .IN1(n34486), .IN2(s15_data_o[3]), .S(n30330), .Q(n17962)
         );
  MUX21X1 U33896 ( .IN1(n34637), .IN2(s15_data_o[4]), .S(n30330), .Q(n17961)
         );
  MUX21X1 U33897 ( .IN1(n34595), .IN2(s15_data_o[5]), .S(n30330), .Q(n17960)
         );
  MUX21X1 U33898 ( .IN1(n34616), .IN2(s15_data_o[6]), .S(n30330), .Q(n17959)
         );
  MUX21X1 U33899 ( .IN1(n34564), .IN2(s15_data_o[7]), .S(n30330), .Q(n17958)
         );
  MUX21X1 U33900 ( .IN1(n34236), .IN2(s15_data_o[8]), .S(n30330), .Q(n17957)
         );
  MUX21X1 U33901 ( .IN1(n34487), .IN2(s15_data_o[9]), .S(n30330), .Q(n17956)
         );
  MUX21X1 U33902 ( .IN1(n34361), .IN2(s15_data_o[10]), .S(n30330), .Q(n17955)
         );
  MUX21X1 U33903 ( .IN1(n34551), .IN2(s15_data_o[11]), .S(n30330), .Q(n17954)
         );
  MUX21X1 U33904 ( .IN1(n34311), .IN2(s15_data_o[12]), .S(n30330), .Q(n17953)
         );
  MUX21X1 U33905 ( .IN1(n34488), .IN2(s15_data_o[13]), .S(n30330), .Q(n17952)
         );
  MUX21X1 U33906 ( .IN1(n34312), .IN2(s15_data_o[14]), .S(n30330), .Q(n17951)
         );
  MUX21X1 U33907 ( .IN1(n34489), .IN2(s15_data_o[15]), .S(n30330), .Q(n17950)
         );
  NOR2X0 U33908 ( .IN1(\s3/msel/gnt_p3 [0]), .IN2(\s3/msel/gnt_p3 [1]), .QN(
        n30396) );
  NAND2X0 U33909 ( .IN1(n30396), .IN2(n30375), .QN(n30343) );
  NOR2X0 U33910 ( .IN1(n30345), .IN2(n30343), .QN(n30333) );
  NAND2X0 U33911 ( .IN1(\s3/msel/gnt_p3 [0]), .IN2(\s3/msel/gnt_p3 [1]), .QN(
        n30402) );
  INVX0 U33912 ( .INP(n30402), .ZN(n30404) );
  NAND2X0 U33913 ( .IN1(\s3/msel/gnt_p3 [1]), .IN2(n34665), .QN(n30376) );
  INVX0 U33914 ( .INP(n30376), .ZN(n30331) );
  NOR2X0 U33915 ( .IN1(n30386), .IN2(n34665), .QN(n30368) );
  INVX0 U33916 ( .INP(n30393), .ZN(n30366) );
  OA21X1 U33917 ( .IN1(n30331), .IN2(n30368), .IN3(n30366), .Q(n30332) );
  NOR3X0 U33918 ( .IN1(n30333), .IN2(n30404), .IN3(n30332), .QN(n30335) );
  INVX0 U33919 ( .INP(n30408), .ZN(n30387) );
  INVX0 U33920 ( .INP(n30375), .ZN(n30410) );
  MUX21X1 U33921 ( .IN1(n30387), .IN2(n30410), .S(\s3/msel/gnt_p3 [0]), .Q(
        n30357) );
  OA222X1 U33922 ( .IN1(n30376), .IN2(n30386), .IN3(n30357), .IN4(
        \s3/msel/gnt_p3 [1]), .IN5(n30402), .IN6(n30393), .Q(n30334) );
  NOR3X0 U33923 ( .IN1(n30336), .IN2(n30335), .IN3(n30334), .QN(n30339) );
  INVX0 U33924 ( .INP(n30374), .ZN(n30364) );
  NAND2X0 U33925 ( .IN1(\s3/msel/gnt_p3 [1]), .IN2(n30364), .QN(n30358) );
  OA21X1 U33926 ( .IN1(\s3/msel/gnt_p3 [1]), .IN2(n30365), .IN3(n30358), .Q(
        n30414) );
  MUX21X1 U33927 ( .IN1(n30388), .IN2(n30398), .S(\s3/msel/gnt_p3 [1]), .Q(
        n30416) );
  OA22X1 U33928 ( .IN1(\s3/msel/gnt_p3 [0]), .IN2(n30416), .IN3(n30345), .IN4(
        n30353), .Q(n30337) );
  NAND2X0 U33929 ( .IN1(n34404), .IN2(n30340), .QN(n30349) );
  NAND3X0 U33930 ( .IN1(n30414), .IN2(n30337), .IN3(n30349), .QN(n30338) );
  MUX21X1 U33931 ( .IN1(n30339), .IN2(n30338), .S(\s3/msel/gnt_p3 [2]), .Q(
        n17949) );
  OA221X1 U33932 ( .IN1(n30347), .IN2(n34404), .IN3(n30347), .IN4(n30398), 
        .IN5(n30344), .Q(n30348) );
  INVX0 U33933 ( .INP(n30340), .ZN(n30341) );
  OA222X1 U33934 ( .IN1(n34404), .IN2(n30353), .IN3(n30374), .IN4(n30410), 
        .IN5(n30396), .IN6(n30341), .Q(n30342) );
  OA22X1 U33935 ( .IN1(n30348), .IN2(n30343), .IN3(n30342), .IN4(n30347), .Q(
        n30356) );
  AO221X1 U33936 ( .IN1(\s3/msel/gnt_p3 [1]), .IN2(\s3/msel/gnt_p3 [0]), .IN3(
        n34404), .IN4(n34665), .IN5(n30344), .Q(n30355) );
  INVX0 U33937 ( .INP(n30365), .ZN(n30399) );
  NAND2X0 U33938 ( .IN1(n30399), .IN2(n30376), .QN(n30346) );
  NAND2X0 U33939 ( .IN1(n30346), .IN2(n30345), .QN(n30352) );
  OA22X1 U33940 ( .IN1(n30348), .IN2(n30402), .IN3(n30347), .IN4(n30376), .Q(
        n30351) );
  OA22X1 U33941 ( .IN1(n30399), .IN2(n30349), .IN3(n30374), .IN4(n30376), .Q(
        n30350) );
  OA221X1 U33942 ( .IN1(n30353), .IN2(n30352), .IN3(n30353), .IN4(n30351), 
        .IN5(n30350), .Q(n30354) );
  OA222X1 U33943 ( .IN1(\s3/msel/gnt_p3 [2]), .IN2(n30356), .IN3(
        \s3/msel/gnt_p3 [2]), .IN4(n30355), .IN5(n30354), .IN6(n34458), .Q(
        n30361) );
  OA21X1 U33944 ( .IN1(n30366), .IN2(n30402), .IN3(n34458), .Q(n30413) );
  OA21X1 U33945 ( .IN1(n30361), .IN2(n30357), .IN3(n30413), .Q(n30363) );
  INVX0 U33946 ( .INP(n30388), .ZN(n30381) );
  OA22X1 U33947 ( .IN1(n30381), .IN2(n30361), .IN3(n34404), .IN4(n30398), .Q(
        n30360) );
  OA21X1 U33948 ( .IN1(n30399), .IN2(n30361), .IN3(n30358), .Q(n30359) );
  OA221X1 U33949 ( .IN1(\s3/msel/gnt_p3 [0]), .IN2(n30360), .IN3(n34665), 
        .IN4(n30359), .IN5(\s3/msel/gnt_p3 [2]), .Q(n30362) );
  OAI22X1 U33950 ( .IN1(n30363), .IN2(n30362), .IN3(n34404), .IN4(n30361), 
        .QN(n17948) );
  INVX0 U33951 ( .INP(n30386), .ZN(n30409) );
  NAND3X0 U33952 ( .IN1(n30364), .IN2(n30388), .IN3(n30398), .QN(n30372) );
  INVX0 U33953 ( .INP(n30372), .ZN(n30369) );
  NAND2X0 U33954 ( .IN1(n30366), .IN2(n30365), .QN(n30367) );
  AND2X1 U33955 ( .IN1(n30398), .IN2(\s3/msel/gnt_p3 [0]), .Q(n30395) );
  AO221X1 U33956 ( .IN1(n30388), .IN2(n30399), .IN3(n30388), .IN4(n30395), 
        .IN5(n30393), .Q(n30370) );
  OA21X1 U33957 ( .IN1(n30408), .IN2(n30367), .IN3(n30370), .Q(n30373) );
  OA21X1 U33958 ( .IN1(n30369), .IN2(n30373), .IN3(n30368), .Q(n30407) );
  AOI21X1 U33959 ( .IN1(n30409), .IN2(n30370), .IN3(n30410), .QN(n30385) );
  INVX0 U33960 ( .INP(n30396), .ZN(n30371) );
  AO221X1 U33961 ( .IN1(n30385), .IN2(n30386), .IN3(n30385), .IN4(n30372), 
        .IN5(n30371), .Q(n30384) );
  INVX0 U33962 ( .INP(n30373), .ZN(n30378) );
  OA21X1 U33963 ( .IN1(n30387), .IN2(n30375), .IN3(n30374), .Q(n30379) );
  NAND2X0 U33964 ( .IN1(n30388), .IN2(n30398), .QN(n30377) );
  AO221X1 U33965 ( .IN1(n30378), .IN2(n30379), .IN3(n30378), .IN4(n30377), 
        .IN5(n30376), .Q(n30383) );
  INVX0 U33966 ( .INP(n30379), .ZN(n30391) );
  AOI21X1 U33967 ( .IN1(n30398), .IN2(n30391), .IN3(n30399), .QN(n30380) );
  OR3X1 U33968 ( .IN1(n30381), .IN2(n30380), .IN3(n30402), .Q(n30382) );
  NAND4X0 U33969 ( .IN1(n34458), .IN2(n30384), .IN3(n30383), .IN4(n30382), 
        .QN(n30406) );
  NOR2X0 U33970 ( .IN1(n30387), .IN2(n30385), .QN(n30403) );
  NOR2X0 U33971 ( .IN1(n30399), .IN2(\s3/msel/gnt_p3 [0]), .QN(n30390) );
  NOR2X0 U33972 ( .IN1(n30387), .IN2(n30386), .QN(n30392) );
  NAND2X0 U33973 ( .IN1(n30388), .IN2(n30392), .QN(n30389) );
  NOR2X0 U33974 ( .IN1(n30390), .IN2(n30389), .QN(n30394) );
  AO21X1 U33975 ( .IN1(n30393), .IN2(n30392), .IN3(n30391), .Q(n30397) );
  OA22X1 U33976 ( .IN1(\s3/msel/gnt_p3 [1]), .IN2(n30395), .IN3(n30394), .IN4(
        n30397), .Q(n30401) );
  OA221X1 U33977 ( .IN1(n30399), .IN2(n30398), .IN3(n30399), .IN4(n30397), 
        .IN5(n30396), .Q(n30400) );
  AO221X1 U33978 ( .IN1(n30404), .IN2(n30403), .IN3(n30402), .IN4(n30401), 
        .IN5(n30400), .Q(n30405) );
  OA22X1 U33979 ( .IN1(n30407), .IN2(n30406), .IN3(n34458), .IN4(n30405), .Q(
        n30415) );
  OAI221X1 U33980 ( .IN1(n34404), .IN2(n30409), .IN3(\s3/msel/gnt_p3 [1]), 
        .IN4(n30408), .IN5(n30415), .QN(n30412) );
  NAND3X0 U33981 ( .IN1(\s3/msel/gnt_p3 [0]), .IN2(n30410), .IN3(n34404), .QN(
        n30411) );
  NAND3X0 U33982 ( .IN1(n30413), .IN2(n30412), .IN3(n30411), .QN(n30419) );
  NOR2X0 U33983 ( .IN1(n30414), .IN2(n34665), .QN(n30418) );
  OA221X1 U33984 ( .IN1(\s3/msel/gnt_p3 [0]), .IN2(\s3/msel/gnt_p3 [2]), .IN3(
        \s3/msel/gnt_p3 [0]), .IN4(n30416), .IN5(n30415), .Q(n30417) );
  AO221X1 U33985 ( .IN1(n30419), .IN2(n30418), .IN3(n30419), .IN4(n34458), 
        .IN5(n30417), .Q(n17947) );
  NOR2X0 U33986 ( .IN1(n30427), .IN2(n30435), .QN(n30420) );
  NOR4X0 U33987 ( .IN1(n30446), .IN2(n30445), .IN3(n30420), .IN4(n34388), .QN(
        n30433) );
  NAND2X0 U33988 ( .IN1(n30434), .IN2(n30421), .QN(n30426) );
  NAND2X0 U33989 ( .IN1(n30423), .IN2(n30422), .QN(n30424) );
  AO22X1 U33990 ( .IN1(n30425), .IN2(n30441), .IN3(n30426), .IN4(n30424), .Q(
        n30432) );
  AO22X1 U33991 ( .IN1(n30427), .IN2(n30426), .IN3(n34658), .IN4(n30440), .Q(
        n30428) );
  OA22X1 U33992 ( .IN1(n19079), .IN2(n30430), .IN3(n30429), .IN4(n30428), .Q(
        n30431) );
  AO222X1 U33993 ( .IN1(n34418), .IN2(n30433), .IN3(n34418), .IN4(n30432), 
        .IN5(n30431), .IN6(\s3/msel/gnt_p1 [2]), .Q(n30454) );
  INVX0 U33994 ( .INP(n30434), .ZN(n30436) );
  OA21X1 U33995 ( .IN1(n30436), .IN2(n30435), .IN3(n30454), .Q(n30443) );
  AO21X1 U33996 ( .IN1(n30438), .IN2(n30443), .IN3(n30437), .Q(n30453) );
  NAND2X0 U33997 ( .IN1(n30440), .IN2(n30439), .QN(n30451) );
  NAND2X0 U33998 ( .IN1(n30442), .IN2(n30441), .QN(n30450) );
  INVX0 U33999 ( .INP(n30443), .ZN(n30444) );
  NOR2X0 U34000 ( .IN1(n30445), .IN2(n30444), .QN(n30448) );
  NAND2X0 U34001 ( .IN1(n30446), .IN2(n34658), .QN(n30447) );
  NAND2X0 U34002 ( .IN1(n30448), .IN2(n30447), .QN(n30449) );
  NAND4X0 U34003 ( .IN1(\s3/msel/gnt_p1 [2]), .IN2(n30451), .IN3(n30450), 
        .IN4(n30449), .QN(n30452) );
  AO22X1 U34004 ( .IN1(\s3/msel/gnt_p1 [1]), .IN2(n30454), .IN3(n30453), .IN4(
        n30452), .Q(n17945) );
  AND3X1 U34005 ( .IN1(n13634), .IN2(n13608), .IN3(m5s3_cyc), .Q(n30510) );
  NAND3X0 U34006 ( .IN1(n13530), .IN2(n13475), .IN3(m7s3_cyc), .QN(n30502) );
  AOI21X1 U34007 ( .IN1(n30502), .IN2(\s3/msel/gnt_p0 [1]), .IN3(n34413), .QN(
        n30483) );
  OA21X1 U34008 ( .IN1(\s3/msel/gnt_p0 [1]), .IN2(n30510), .IN3(n30483), .Q(
        n30535) );
  INVX0 U34009 ( .INP(n30535), .ZN(n30466) );
  NOR2X0 U34010 ( .IN1(\s3/msel/gnt_p0 [0]), .IN2(n34263), .QN(n30467) );
  AND3X1 U34011 ( .IN1(n13790), .IN2(n13764), .IN3(m2s3_cyc), .Q(n30520) );
  NAND2X0 U34012 ( .IN1(n30467), .IN2(n30520), .QN(n30455) );
  NAND3X0 U34013 ( .IN1(n13738), .IN2(n13712), .IN3(m3s3_cyc), .QN(n30456) );
  INVX0 U34014 ( .INP(n30456), .ZN(n30501) );
  NOR2X0 U34015 ( .IN1(n34393), .IN2(n34263), .QN(n30458) );
  NAND2X0 U34016 ( .IN1(n30501), .IN2(n30458), .QN(n30533) );
  NAND3X0 U34017 ( .IN1(n30455), .IN2(n30533), .IN3(n34413), .QN(n30489) );
  NOR2X0 U34018 ( .IN1(n30520), .IN2(n30501), .QN(n30472) );
  NAND3X0 U34019 ( .IN1(n13842), .IN2(n13816), .IN3(m1s3_cyc), .QN(n30503) );
  AND2X1 U34020 ( .IN1(n34263), .IN2(n30503), .Q(n30473) );
  AO22X1 U34021 ( .IN1(n30472), .IN2(n30473), .IN3(n30467), .IN4(n30456), .Q(
        n30457) );
  NAND3X0 U34022 ( .IN1(n13902), .IN2(n13868), .IN3(m0s3_cyc), .QN(n30514) );
  OR2X1 U34023 ( .IN1(n34393), .IN2(n30503), .Q(n30530) );
  OA21X1 U34024 ( .IN1(\s3/msel/gnt_p0 [0]), .IN2(n30514), .IN3(n30530), .Q(
        n30490) );
  OAI22X1 U34025 ( .IN1(n30458), .IN2(n30457), .IN3(\s3/msel/gnt_p0 [1]), 
        .IN4(n30490), .QN(n30459) );
  NOR2X0 U34026 ( .IN1(n30489), .IN2(n30459), .QN(n30461) );
  NAND3X0 U34027 ( .IN1(n13582), .IN2(n13556), .IN3(m6s3_cyc), .QN(n30512) );
  NAND2X0 U34028 ( .IN1(n30512), .IN2(n30502), .QN(n30462) );
  INVX0 U34029 ( .INP(n30462), .ZN(n30469) );
  NAND3X0 U34030 ( .IN1(n13686), .IN2(n13660), .IN3(m4s3_cyc), .QN(n30523) );
  INVX0 U34031 ( .INP(n30523), .ZN(n30504) );
  NOR2X0 U34032 ( .IN1(n30504), .IN2(n30510), .QN(n30470) );
  NAND2X0 U34033 ( .IN1(n30469), .IN2(n30470), .QN(n30460) );
  NAND2X0 U34034 ( .IN1(n30461), .IN2(n30460), .QN(n30465) );
  NAND2X0 U34035 ( .IN1(n34263), .IN2(n30462), .QN(n30477) );
  MUX21X1 U34036 ( .IN1(n30523), .IN2(n30512), .S(\s3/msel/gnt_p0 [1]), .Q(
        n30500) );
  AO221X1 U34037 ( .IN1(n30477), .IN2(\s3/msel/gnt_p0 [0]), .IN3(n30477), 
        .IN4(n30500), .IN5(n34413), .Q(n30464) );
  AND3X1 U34038 ( .IN1(\s3/msel/gnt_p0 [2]), .IN2(n30514), .IN3(n30503), .Q(
        n30481) );
  NAND2X0 U34039 ( .IN1(n30472), .IN2(n30481), .QN(n30463) );
  NAND4X0 U34040 ( .IN1(n30466), .IN2(n30465), .IN3(n30464), .IN4(n30463), 
        .QN(n17943) );
  NAND2X0 U34041 ( .IN1(n30467), .IN2(n30501), .QN(n30476) );
  NAND2X0 U34042 ( .IN1(n30514), .IN2(n30503), .QN(n30468) );
  NAND2X0 U34043 ( .IN1(n30469), .IN2(n30468), .QN(n30484) );
  NAND3X0 U34044 ( .IN1(\s3/msel/gnt_p0 [1]), .IN2(n30470), .IN3(n30484), .QN(
        n30475) );
  NAND2X0 U34045 ( .IN1(n30469), .IN2(n30472), .QN(n30479) );
  INVX0 U34046 ( .INP(n30470), .ZN(n30471) );
  NAND2X0 U34047 ( .IN1(n30472), .IN2(n30471), .QN(n30478) );
  NAND3X0 U34048 ( .IN1(n30479), .IN2(n30478), .IN3(n30473), .QN(n30474) );
  NAND3X0 U34049 ( .IN1(n30476), .IN2(n30475), .IN3(n30474), .QN(n30488) );
  NOR2X0 U34050 ( .IN1(\s3/msel/gnt_p0 [0]), .IN2(\s3/msel/gnt_p0 [1]), .QN(
        n30528) );
  INVX0 U34051 ( .INP(n30528), .ZN(n30521) );
  NOR2X0 U34052 ( .IN1(n30479), .IN2(n30521), .QN(n30487) );
  NAND2X0 U34053 ( .IN1(\s3/msel/gnt_p0 [0]), .IN2(n30477), .QN(n30482) );
  OA21X1 U34054 ( .IN1(\s3/msel/gnt_p0 [1]), .IN2(n30479), .IN3(n30478), .Q(
        n30480) );
  AO22X1 U34055 ( .IN1(n30483), .IN2(n30482), .IN3(n30481), .IN4(n30480), .Q(
        n30485) );
  NAND2X0 U34056 ( .IN1(n30485), .IN2(n30484), .QN(n30486) );
  NOR2X0 U34057 ( .IN1(n30487), .IN2(n30486), .QN(n30491) );
  AO21X1 U34058 ( .IN1(n34413), .IN2(n30488), .IN3(n30491), .Q(n30499) );
  AO21X1 U34059 ( .IN1(n30490), .IN2(n30499), .IN3(n30489), .Q(n30498) );
  AO221X1 U34060 ( .IN1(\s3/msel/gnt_p0 [0]), .IN2(n30502), .IN3(n34393), 
        .IN4(n30512), .IN5(n34263), .Q(n30496) );
  INVX0 U34061 ( .INP(n30491), .ZN(n30492) );
  NOR2X0 U34062 ( .IN1(n30510), .IN2(n30492), .QN(n30494) );
  NAND2X0 U34063 ( .IN1(n30504), .IN2(n34393), .QN(n30493) );
  NAND2X0 U34064 ( .IN1(n30494), .IN2(n30493), .QN(n30495) );
  NAND3X0 U34065 ( .IN1(\s3/msel/gnt_p0 [2]), .IN2(n30496), .IN3(n30495), .QN(
        n30497) );
  AO22X1 U34066 ( .IN1(\s3/msel/gnt_p0 [1]), .IN2(n30499), .IN3(n30498), .IN4(
        n30497), .Q(n17942) );
  AO21X1 U34067 ( .IN1(\s3/msel/gnt_p0 [2]), .IN2(n30500), .IN3(
        \s3/msel/gnt_p0 [0]), .Q(n30538) );
  INVX0 U34068 ( .INP(n30514), .ZN(n30531) );
  NAND2X0 U34069 ( .IN1(n30523), .IN2(n30512), .QN(n30515) );
  AO21X1 U34070 ( .IN1(n30510), .IN2(n30523), .IN3(n30501), .Q(n30513) );
  INVX0 U34071 ( .INP(n30513), .ZN(n30505) );
  OA21X1 U34072 ( .IN1(n34393), .IN2(n30515), .IN3(n30505), .Q(n30518) );
  OA21X1 U34073 ( .IN1(n30520), .IN2(n30518), .IN3(n30503), .Q(n30522) );
  OR3X1 U34074 ( .IN1(n34263), .IN2(n30531), .IN3(n30522), .Q(n30509) );
  OA21X1 U34075 ( .IN1(n30531), .IN2(n30503), .IN3(n30502), .Q(n30516) );
  AO221X1 U34076 ( .IN1(n30505), .IN2(n30504), .IN3(n30505), .IN4(n34393), 
        .IN5(n30520), .Q(n30507) );
  INVX0 U34077 ( .INP(n30512), .ZN(n30506) );
  AO221X1 U34078 ( .IN1(n30516), .IN2(n30531), .IN3(n30516), .IN4(n30507), 
        .IN5(n30506), .Q(n30508) );
  NAND3X0 U34079 ( .IN1(\s3/msel/gnt_p0 [2]), .IN2(n30509), .IN3(n30508), .QN(
        n30529) );
  INVX0 U34080 ( .INP(n30516), .ZN(n30511) );
  AO21X1 U34081 ( .IN1(n30512), .IN2(n30511), .IN3(n30510), .Q(n30527) );
  NOR2X0 U34082 ( .IN1(n30514), .IN2(n30513), .QN(n30517) );
  OA22X1 U34083 ( .IN1(n30518), .IN2(n30517), .IN3(n30516), .IN4(n30515), .Q(
        n30519) );
  OA22X1 U34084 ( .IN1(n30522), .IN2(n30521), .IN3(n30520), .IN4(n30519), .Q(
        n30525) );
  NAND4X0 U34085 ( .IN1(\s3/msel/gnt_p0 [1]), .IN2(\s3/msel/gnt_p0 [0]), .IN3(
        n30523), .IN4(n30527), .QN(n30524) );
  NAND3X0 U34086 ( .IN1(n30525), .IN2(n34413), .IN3(n30524), .QN(n30526) );
  OA221X1 U34087 ( .IN1(n30529), .IN2(n30528), .IN3(n30529), .IN4(n30527), 
        .IN5(n30526), .Q(n30537) );
  INVX0 U34088 ( .INP(n30537), .ZN(n30532) );
  OA222X1 U34089 ( .IN1(n30532), .IN2(n30531), .IN3(n30532), .IN4(n34263), 
        .IN5(\s3/msel/gnt_p0 [1]), .IN6(n30530), .Q(n30534) );
  NAND2X0 U34090 ( .IN1(n30534), .IN2(n30533), .QN(n30536) );
  AO222X1 U34091 ( .IN1(n30538), .IN2(n30537), .IN3(n34413), .IN4(n30536), 
        .IN5(n30535), .IN6(\s3/msel/gnt_p0 [0]), .Q(n17941) );
  MUX21X1 U34092 ( .IN1(n30549), .IN2(n30594), .S(\s3/msel/gnt_p2 [1]), .Q(
        n30620) );
  INVX0 U34093 ( .INP(n30620), .ZN(n30540) );
  NAND2X0 U34094 ( .IN1(\s3/msel/gnt_p2 [1]), .IN2(n30579), .QN(n30558) );
  OR2X1 U34095 ( .IN1(n30557), .IN2(n30618), .Q(n30539) );
  AO22X1 U34096 ( .IN1(n34416), .IN2(n30540), .IN3(n30558), .IN4(n30539), .Q(
        n30547) );
  OR2X1 U34097 ( .IN1(n30580), .IN2(n34416), .Q(n30613) );
  OA21X1 U34098 ( .IN1(\s3/msel/gnt_p2 [0]), .IN2(n30591), .IN3(n30613), .Q(
        n30568) );
  NOR2X0 U34099 ( .IN1(\s3/msel/gnt_p2 [1]), .IN2(n30568), .QN(n30545) );
  INVX0 U34100 ( .INP(n30541), .ZN(n30561) );
  AND2X1 U34101 ( .IN1(n34287), .IN2(n30580), .Q(n30554) );
  AOI22X1 U34102 ( .IN1(\s3/msel/gnt_p2 [1]), .IN2(n30576), .IN3(n30561), 
        .IN4(n30554), .QN(n30543) );
  INVX0 U34103 ( .INP(n30610), .ZN(n30584) );
  NOR2X0 U34104 ( .IN1(\s3/msel/gnt_p2 [0]), .IN2(n34287), .QN(n30569) );
  NAND2X0 U34105 ( .IN1(\s3/msel/gnt_p2 [1]), .IN2(\s3/msel/gnt_p2 [0]), .QN(
        n30552) );
  OA21X1 U34106 ( .IN1(n30552), .IN2(n30576), .IN3(n34650), .Q(n30616) );
  INVX0 U34107 ( .INP(n30616), .ZN(n30542) );
  AO21X1 U34108 ( .IN1(n30584), .IN2(n30569), .IN3(n30542), .Q(n30567) );
  NOR4X0 U34109 ( .IN1(n30545), .IN2(n30544), .IN3(n30543), .IN4(n30567), .QN(
        n30546) );
  AO221X1 U34110 ( .IN1(\s3/msel/gnt_p2 [2]), .IN2(n30548), .IN3(
        \s3/msel/gnt_p2 [2]), .IN4(n30547), .IN5(n30546), .Q(n17940) );
  NAND4X0 U34111 ( .IN1(n30591), .IN2(n30580), .IN3(n30549), .IN4(n30577), 
        .QN(n30556) );
  NAND3X0 U34112 ( .IN1(n30549), .IN2(n30577), .IN3(n30557), .QN(n30550) );
  NAND3X0 U34113 ( .IN1(n30576), .IN2(n30556), .IN3(n30550), .QN(n30555) );
  NAND2X0 U34114 ( .IN1(n30561), .IN2(n30550), .QN(n30553) );
  OA21X1 U34115 ( .IN1(n30557), .IN2(n30551), .IN3(n30577), .Q(n30563) );
  NOR2X0 U34116 ( .IN1(n30597), .IN2(n30552), .QN(n30608) );
  AO222X1 U34117 ( .IN1(n30555), .IN2(n30569), .IN3(n30554), .IN4(n30553), 
        .IN5(n30563), .IN6(n30608), .Q(n30566) );
  INVX0 U34118 ( .INP(n30556), .ZN(n30559) );
  OA22X1 U34119 ( .IN1(n30559), .IN2(n30558), .IN3(\s3/msel/gnt_p2 [1]), .IN4(
        n30557), .Q(n30564) );
  NOR2X0 U34120 ( .IN1(\s3/msel/gnt_p2 [1]), .IN2(\s3/msel/gnt_p2 [0]), .QN(
        n30602) );
  INVX0 U34121 ( .INP(n30602), .ZN(n30589) );
  NOR2X0 U34122 ( .IN1(n30561), .IN2(n30560), .QN(n30562) );
  AO221X1 U34123 ( .IN1(n30564), .IN2(n30563), .IN3(n30564), .IN4(n30589), 
        .IN5(n30562), .Q(n30565) );
  MUX21X1 U34124 ( .IN1(n30566), .IN2(n30565), .S(\s3/msel/gnt_p2 [2]), .Q(
        n30575) );
  AO21X1 U34125 ( .IN1(n30568), .IN2(n30575), .IN3(n30567), .Q(n30574) );
  INVX0 U34126 ( .INP(n30594), .ZN(n30599) );
  NAND2X0 U34127 ( .IN1(n30569), .IN2(n30599), .QN(n30572) );
  NAND2X0 U34128 ( .IN1(n30597), .IN2(n34416), .QN(n30570) );
  NAND3X0 U34129 ( .IN1(n30577), .IN2(n30575), .IN3(n30570), .QN(n30571) );
  NAND3X0 U34130 ( .IN1(n30572), .IN2(n30571), .IN3(\s3/msel/gnt_p2 [2]), .QN(
        n30573) );
  AO22X1 U34131 ( .IN1(\s3/msel/gnt_p2 [1]), .IN2(n30575), .IN3(n30574), .IN4(
        n30573), .Q(n17939) );
  NOR2X0 U34132 ( .IN1(n30597), .IN2(n30599), .QN(n30582) );
  INVX0 U34133 ( .INP(n30579), .ZN(n30617) );
  NAND3X0 U34134 ( .IN1(n30610), .IN2(n30582), .IN3(n30617), .QN(n30578) );
  OA21X1 U34135 ( .IN1(n30597), .IN2(n30577), .IN3(n30576), .Q(n30598) );
  OA21X1 U34136 ( .IN1(n30584), .IN2(n30598), .IN3(n30580), .Q(n30595) );
  NAND2X0 U34137 ( .IN1(n30578), .IN2(n30595), .QN(n30590) );
  INVX0 U34138 ( .INP(n30591), .ZN(n30612) );
  OA21X1 U34139 ( .IN1(n30612), .IN2(n30580), .IN3(n30579), .Q(n30601) );
  INVX0 U34140 ( .INP(n30582), .ZN(n30581) );
  NOR2X0 U34141 ( .IN1(n30601), .IN2(n30581), .QN(n30587) );
  NAND3X0 U34142 ( .IN1(n30582), .IN2(\s3/msel/gnt_p2 [0]), .IN3(n30591), .QN(
        n30583) );
  NAND2X0 U34143 ( .IN1(n30583), .IN2(n30598), .QN(n30586) );
  NOR2X0 U34144 ( .IN1(n30584), .IN2(\s3/msel/gnt_p2 [1]), .QN(n30585) );
  OA22X1 U34145 ( .IN1(n30587), .IN2(n30586), .IN3(n30585), .IN4(n34416), .Q(
        n30588) );
  AO221X1 U34146 ( .IN1(n30602), .IN2(n30590), .IN3(n30589), .IN4(n30588), 
        .IN5(\s3/msel/gnt_p2 [2]), .Q(n30609) );
  NAND2X0 U34147 ( .IN1(n30610), .IN2(n30591), .QN(n30596) );
  NOR2X0 U34148 ( .IN1(n34416), .IN2(n30596), .QN(n30593) );
  INVX0 U34149 ( .INP(n30601), .ZN(n30592) );
  AO221X1 U34150 ( .IN1(n30594), .IN2(n30593), .IN3(n30594), .IN4(n30592), 
        .IN5(n30618), .Q(n30607) );
  OR3X1 U34151 ( .IN1(n34287), .IN2(n30612), .IN3(n30595), .Q(n30605) );
  AO221X1 U34152 ( .IN1(n30598), .IN2(n30597), .IN3(n30598), .IN4(n34416), 
        .IN5(n30596), .Q(n30600) );
  AO21X1 U34153 ( .IN1(n30601), .IN2(n30600), .IN3(n30599), .Q(n30604) );
  NAND2X0 U34154 ( .IN1(n30602), .IN2(n30607), .QN(n30603) );
  NAND4X0 U34155 ( .IN1(\s3/msel/gnt_p2 [2]), .IN2(n30605), .IN3(n30604), 
        .IN4(n30603), .QN(n30606) );
  OA221X1 U34156 ( .IN1(n30609), .IN2(n30608), .IN3(n30609), .IN4(n30607), 
        .IN5(n30606), .Q(n30619) );
  NAND3X0 U34157 ( .IN1(\s3/msel/gnt_p2 [1]), .IN2(n30619), .IN3(n30610), .QN(
        n30615) );
  INVX0 U34158 ( .INP(n30619), .ZN(n30611) );
  AO221X1 U34159 ( .IN1(n30613), .IN2(n30612), .IN3(n30613), .IN4(n30611), 
        .IN5(\s3/msel/gnt_p2 [1]), .Q(n30614) );
  NAND3X0 U34160 ( .IN1(n30616), .IN2(n30615), .IN3(n30614), .QN(n30623) );
  OA221X1 U34161 ( .IN1(\s3/msel/gnt_p2 [1]), .IN2(n30618), .IN3(n34287), 
        .IN4(n30617), .IN5(\s3/msel/gnt_p2 [0]), .Q(n30622) );
  OA221X1 U34162 ( .IN1(\s3/msel/gnt_p2 [0]), .IN2(\s3/msel/gnt_p2 [2]), .IN3(
        \s3/msel/gnt_p2 [0]), .IN4(n30620), .IN5(n30619), .Q(n30621) );
  AO221X1 U34163 ( .IN1(n30623), .IN2(n34650), .IN3(n30623), .IN4(n30622), 
        .IN5(n30621), .Q(n17938) );
  NOR2X0 U34164 ( .IN1(n30624), .IN2(n34379), .QN(n30625) );
  MUX21X1 U34165 ( .IN1(n34340), .IN2(s15_data_o[0]), .S(n30625), .Q(n17937)
         );
  MUX21X1 U34166 ( .IN1(n34490), .IN2(s15_data_o[1]), .S(n30625), .Q(n17936)
         );
  MUX21X1 U34167 ( .IN1(n34315), .IN2(s15_data_o[2]), .S(n30625), .Q(n17935)
         );
  MUX21X1 U34168 ( .IN1(n34491), .IN2(s15_data_o[3]), .S(n30625), .Q(n17934)
         );
  MUX21X1 U34169 ( .IN1(n34627), .IN2(s15_data_o[4]), .S(n30625), .Q(n17933)
         );
  MUX21X1 U34170 ( .IN1(n34577), .IN2(s15_data_o[5]), .S(n30625), .Q(n17932)
         );
  MUX21X1 U34171 ( .IN1(n34617), .IN2(s15_data_o[6]), .S(n30625), .Q(n17931)
         );
  MUX21X1 U34172 ( .IN1(n34578), .IN2(s15_data_o[7]), .S(n30625), .Q(n17930)
         );
  MUX21X1 U34173 ( .IN1(n34338), .IN2(s15_data_o[8]), .S(n30625), .Q(n17929)
         );
  MUX21X1 U34174 ( .IN1(n34525), .IN2(s15_data_o[9]), .S(n30625), .Q(n17928)
         );
  MUX21X1 U34175 ( .IN1(n34313), .IN2(s15_data_o[10]), .S(n30625), .Q(n17927)
         );
  MUX21X1 U34176 ( .IN1(n34492), .IN2(s15_data_o[11]), .S(n30625), .Q(n17926)
         );
  MUX21X1 U34177 ( .IN1(n34339), .IN2(s15_data_o[12]), .S(n30625), .Q(n17925)
         );
  MUX21X1 U34178 ( .IN1(n34526), .IN2(s15_data_o[13]), .S(n30625), .Q(n17924)
         );
  MUX21X1 U34179 ( .IN1(n34314), .IN2(s15_data_o[14]), .S(n30625), .Q(n17923)
         );
  MUX21X1 U34180 ( .IN1(n34527), .IN2(s15_data_o[15]), .S(n30625), .Q(n17922)
         );
  NOR2X0 U34181 ( .IN1(\s4/msel/gnt_p3 [1]), .IN2(n30681), .QN(n30634) );
  NOR2X0 U34182 ( .IN1(n34656), .IN2(n30690), .QN(n30654) );
  NOR2X0 U34183 ( .IN1(n30634), .IN2(n30654), .QN(n30715) );
  INVX0 U34184 ( .INP(n30626), .ZN(n30638) );
  OA221X1 U34185 ( .IN1(\s4/msel/gnt_p3 [1]), .IN2(n30678), .IN3(n34656), 
        .IN4(n30679), .IN5(\s4/msel/gnt_p3 [2]), .Q(n30703) );
  NAND2X0 U34186 ( .IN1(\s4/msel/gnt_p3 [0]), .IN2(\s4/msel/gnt_p3 [2]), .QN(
        n30716) );
  INVX0 U34187 ( .INP(n30716), .ZN(n30665) );
  OA22X1 U34188 ( .IN1(\s4/msel/gnt_p3 [1]), .IN2(n30638), .IN3(n30703), .IN4(
        n30665), .Q(n30627) );
  NAND2X0 U34189 ( .IN1(n30715), .IN2(n30627), .QN(n30633) );
  NOR2X0 U34190 ( .IN1(\s4/msel/gnt_p3 [1]), .IN2(n34455), .QN(n30648) );
  INVX0 U34191 ( .INP(n30648), .ZN(n30704) );
  NAND2X0 U34192 ( .IN1(n34656), .IN2(n30705), .QN(n30646) );
  NAND2X0 U34193 ( .IN1(n34455), .IN2(\s4/msel/gnt_p3 [1]), .QN(n30656) );
  OA221X1 U34194 ( .IN1(n30707), .IN2(n30704), .IN3(n30707), .IN4(n30646), 
        .IN5(n30656), .Q(n30628) );
  NOR2X0 U34195 ( .IN1(n34455), .IN2(n34656), .QN(n30697) );
  INVX0 U34196 ( .INP(n30697), .ZN(n30629) );
  OA21X1 U34197 ( .IN1(n30666), .IN2(n30628), .IN3(n30629), .Q(n30631) );
  INVX0 U34198 ( .INP(n30667), .ZN(n30706) );
  INVX0 U34199 ( .INP(n30705), .ZN(n30640) );
  MUX21X1 U34200 ( .IN1(n30706), .IN2(n30640), .S(\s4/msel/gnt_p3 [0]), .Q(
        n30655) );
  OA222X1 U34201 ( .IN1(n30629), .IN2(n30666), .IN3(n30655), .IN4(
        \s4/msel/gnt_p3 [1]), .IN5(n30656), .IN6(n30707), .Q(n30630) );
  NOR3X0 U34202 ( .IN1(n34101), .IN2(n30631), .IN3(n30630), .QN(n30632) );
  OA22X1 U34203 ( .IN1(n34100), .IN2(n30633), .IN3(\s4/msel/gnt_p3 [2]), .IN4(
        n30632), .Q(n17921) );
  INVX0 U34204 ( .INP(n30634), .ZN(n30676) );
  INVX0 U34205 ( .INP(n30641), .ZN(n30635) );
  INVX0 U34206 ( .INP(n30679), .ZN(n30673) );
  AO221X1 U34207 ( .IN1(n30635), .IN2(\s4/msel/gnt_p3 [1]), .IN3(n30635), 
        .IN4(n30673), .IN5(n30647), .Q(n30644) );
  NAND4X0 U34208 ( .IN1(n30667), .IN2(n30705), .IN3(n30676), .IN4(n30644), 
        .QN(n30637) );
  NAND2X0 U34209 ( .IN1(n34455), .IN2(n30681), .QN(n30669) );
  AO21X1 U34210 ( .IN1(n30669), .IN2(n30704), .IN3(n30638), .Q(n30636) );
  AND3X1 U34211 ( .IN1(\s4/msel/gnt_p3 [2]), .IN2(n30637), .IN3(n30636), .Q(
        n30653) );
  NAND2X0 U34212 ( .IN1(n30697), .IN2(n30667), .QN(n30674) );
  AND2X1 U34213 ( .IN1(n30674), .IN2(n30690), .Q(n30639) );
  OA22X1 U34214 ( .IN1(n30640), .IN2(n30639), .IN3(n34656), .IN4(n30638), .Q(
        n30643) );
  AO221X1 U34215 ( .IN1(n30643), .IN2(n30642), .IN3(n30643), .IN4(n30656), 
        .IN5(n30641), .Q(n30651) );
  INVX0 U34216 ( .INP(n30644), .ZN(n30645) );
  AO221X1 U34217 ( .IN1(n30646), .IN2(n30656), .IN3(n30646), .IN4(n30682), 
        .IN5(n30645), .Q(n30650) );
  NAND2X0 U34218 ( .IN1(n30648), .IN2(n30647), .QN(n30649) );
  AND4X1 U34219 ( .IN1(n30651), .IN2(n34465), .IN3(n30650), .IN4(n30649), .Q(
        n30652) );
  AO221X1 U34220 ( .IN1(n30653), .IN2(n30656), .IN3(n30653), .IN4(n30690), 
        .IN5(n30652), .Q(n30661) );
  INVX0 U34221 ( .INP(n30661), .ZN(n30659) );
  AO21X1 U34222 ( .IN1(n30659), .IN2(n30681), .IN3(n30654), .Q(n30664) );
  AO21X1 U34223 ( .IN1(\s4/msel/gnt_p3 [1]), .IN2(n30673), .IN3(n34465), .Q(
        n30660) );
  OA22X1 U34224 ( .IN1(n30668), .IN2(n30656), .IN3(n30661), .IN4(n30655), .Q(
        n30657) );
  NAND2X0 U34225 ( .IN1(n30666), .IN2(n30697), .QN(n30709) );
  NAND3X0 U34226 ( .IN1(n30657), .IN2(n34465), .IN3(n30709), .QN(n30658) );
  OA221X1 U34227 ( .IN1(n30660), .IN2(n30659), .IN3(n30660), .IN4(n30678), 
        .IN5(n30658), .Q(n30663) );
  NOR2X0 U34228 ( .IN1(n34656), .IN2(n30661), .QN(n30662) );
  AO221X1 U34229 ( .IN1(n30665), .IN2(n30664), .IN3(n30716), .IN4(n30663), 
        .IN5(n30662), .Q(n17920) );
  INVX0 U34230 ( .INP(n30681), .ZN(n30694) );
  OA221X1 U34231 ( .IN1(n30694), .IN2(\s4/msel/gnt_p3 [0]), .IN3(n30694), 
        .IN4(n30679), .IN5(n30678), .Q(n30695) );
  NOR2X0 U34232 ( .IN1(n30666), .IN2(n30695), .QN(n30683) );
  OA21X1 U34233 ( .IN1(n30707), .IN2(n30683), .IN3(n30705), .Q(n30677) );
  NAND2X0 U34234 ( .IN1(n30668), .IN2(n30667), .QN(n30671) );
  NAND2X0 U34235 ( .IN1(n30678), .IN2(n30669), .QN(n30670) );
  OA21X1 U34236 ( .IN1(n30706), .IN2(n30705), .IN3(n30690), .Q(n30680) );
  OA221X1 U34237 ( .IN1(n30671), .IN2(n30682), .IN3(n30671), .IN4(n30670), 
        .IN5(n30680), .Q(n30672) );
  OA22X1 U34238 ( .IN1(n30677), .IN2(n30674), .IN3(n30673), .IN4(n30672), .Q(
        n30675) );
  NAND3X0 U34239 ( .IN1(n30676), .IN2(n30675), .IN3(\s4/msel/gnt_p3 [2]), .QN(
        n30702) );
  NOR2X0 U34240 ( .IN1(n30677), .IN2(\s4/msel/gnt_p3 [0]), .QN(n30687) );
  NAND2X0 U34241 ( .IN1(n30679), .IN2(n30678), .QN(n30689) );
  NOR2X0 U34242 ( .IN1(n30680), .IN2(n30689), .QN(n30693) );
  AND3X1 U34243 ( .IN1(n30682), .IN2(n30681), .IN3(n30706), .Q(n30684) );
  NOR2X0 U34244 ( .IN1(n30684), .IN2(n30683), .QN(n30688) );
  NOR2X0 U34245 ( .IN1(n30693), .IN2(n30688), .QN(n30685) );
  NAND2X0 U34246 ( .IN1(\s4/msel/gnt_p3 [1]), .IN2(n30685), .QN(n30686) );
  NAND2X0 U34247 ( .IN1(n30687), .IN2(n30686), .QN(n30700) );
  INVX0 U34248 ( .INP(n30688), .ZN(n30692) );
  OR2X1 U34249 ( .IN1(n30690), .IN2(n30689), .Q(n30691) );
  AO21X1 U34250 ( .IN1(n30692), .IN2(n30691), .IN3(n30707), .Q(n30699) );
  AO21X1 U34251 ( .IN1(n30695), .IN2(n30694), .IN3(n30693), .Q(n30696) );
  NAND2X0 U34252 ( .IN1(n30697), .IN2(n30696), .QN(n30698) );
  NAND4X0 U34253 ( .IN1(n30700), .IN2(n34465), .IN3(n30699), .IN4(n30698), 
        .QN(n30701) );
  NAND2X0 U34254 ( .IN1(n30702), .IN2(n30701), .QN(n30714) );
  NOR2X0 U34255 ( .IN1(\s4/msel/gnt_p3 [0]), .IN2(n30703), .QN(n30713) );
  NOR2X0 U34256 ( .IN1(n30705), .IN2(n30704), .QN(n30711) );
  AO221X1 U34257 ( .IN1(\s4/msel/gnt_p3 [1]), .IN2(n30707), .IN3(n34656), 
        .IN4(n30706), .IN5(n30714), .Q(n30708) );
  NAND2X0 U34258 ( .IN1(n30709), .IN2(n30708), .QN(n30710) );
  NOR2X0 U34259 ( .IN1(n30711), .IN2(n30710), .QN(n30712) );
  OAI222X1 U34260 ( .IN1(n30716), .IN2(n30715), .IN3(n30714), .IN4(n30713), 
        .IN5(n30712), .IN6(\s4/msel/gnt_p3 [2]), .QN(n17919) );
  NAND2X0 U34261 ( .IN1(n30718), .IN2(n30717), .QN(n30728) );
  INVX0 U34262 ( .INP(n30723), .ZN(n30719) );
  NAND2X0 U34263 ( .IN1(n30719), .IN2(n30721), .QN(n30736) );
  NAND2X0 U34264 ( .IN1(n30721), .IN2(n30720), .QN(n30730) );
  NAND3X0 U34265 ( .IN1(n30736), .IN2(n30730), .IN3(n30722), .QN(n30727) );
  OA21X1 U34266 ( .IN1(n30724), .IN2(n30723), .IN3(n30754), .Q(n30737) );
  NAND3X0 U34267 ( .IN1(\s4/msel/gnt_p1 [1]), .IN2(n30737), .IN3(n30725), .QN(
        n30726) );
  NAND3X0 U34268 ( .IN1(n30728), .IN2(n30727), .IN3(n30726), .QN(n30739) );
  NAND2X0 U34269 ( .IN1(n34246), .IN2(n34389), .QN(n30768) );
  NAND2X0 U34270 ( .IN1(n30729), .IN2(n34246), .QN(n30734) );
  OR2X1 U34271 ( .IN1(\s4/msel/gnt_p1 [1]), .IN2(n30736), .Q(n30731) );
  NAND4X0 U34272 ( .IN1(n30751), .IN2(n30753), .IN3(n30731), .IN4(n30730), 
        .QN(n30732) );
  NAND3X0 U34273 ( .IN1(n30734), .IN2(n30733), .IN3(n30732), .QN(n30735) );
  OA221X1 U34274 ( .IN1(n30768), .IN2(n30737), .IN3(n30768), .IN4(n30736), 
        .IN5(n30735), .Q(n30738) );
  MUX21X1 U34275 ( .IN1(n30739), .IN2(n30738), .S(\s4/msel/gnt_p1 [2]), .Q(
        n30748) );
  AO21X1 U34276 ( .IN1(n30741), .IN2(n30748), .IN3(n30740), .Q(n30747) );
  AO221X1 U34277 ( .IN1(\s4/msel/gnt_p1 [0]), .IN2(n30752), .IN3(n34246), 
        .IN4(n30742), .IN5(n34389), .Q(n30745) );
  NAND2X0 U34278 ( .IN1(n30762), .IN2(n34246), .QN(n30743) );
  NAND3X0 U34279 ( .IN1(n30743), .IN2(n30748), .IN3(n30754), .QN(n30744) );
  NAND3X0 U34280 ( .IN1(\s4/msel/gnt_p1 [2]), .IN2(n30745), .IN3(n30744), .QN(
        n30746) );
  AO22X1 U34281 ( .IN1(\s4/msel/gnt_p1 [1]), .IN2(n30748), .IN3(n30747), .IN4(
        n30746), .Q(n17917) );
  OA21X1 U34282 ( .IN1(n30762), .IN2(n30754), .IN3(n30749), .Q(n30767) );
  OAI21X1 U34283 ( .IN1(n30764), .IN2(n30767), .IN3(n30753), .QN(n30769) );
  NAND3X0 U34284 ( .IN1(\s4/msel/gnt_p1 [1]), .IN2(n30769), .IN3(n30751), .QN(
        n30760) );
  NAND2X0 U34285 ( .IN1(n30751), .IN2(n30750), .QN(n30755) );
  OA21X1 U34286 ( .IN1(n30777), .IN2(n30753), .IN3(n30752), .Q(n30763) );
  OA21X1 U34287 ( .IN1(n34246), .IN2(n30755), .IN3(n30763), .Q(n30757) );
  OA21X1 U34288 ( .IN1(n30766), .IN2(n30757), .IN3(n30754), .Q(n30761) );
  AND2X1 U34289 ( .IN1(n30763), .IN2(n30762), .Q(n30756) );
  OA22X1 U34290 ( .IN1(n30757), .IN2(n30756), .IN3(n30767), .IN4(n30755), .Q(
        n30758) );
  OA22X1 U34291 ( .IN1(n30761), .IN2(n30768), .IN3(n30766), .IN4(n30758), .Q(
        n30759) );
  NAND3X0 U34292 ( .IN1(n30760), .IN2(n30759), .IN3(\s4/msel/gnt_p1 [2]), .QN(
        n30775) );
  OR4X1 U34293 ( .IN1(n34389), .IN2(n34246), .IN3(n30761), .IN4(n30762), .Q(
        n30773) );
  AO221X1 U34294 ( .IN1(n30763), .IN2(n30777), .IN3(n30763), .IN4(n34246), 
        .IN5(n30762), .Q(n30765) );
  AO221X1 U34295 ( .IN1(n30767), .IN2(n30766), .IN3(n30767), .IN4(n30765), 
        .IN5(n30764), .Q(n30772) );
  INVX0 U34296 ( .INP(n30768), .ZN(n30770) );
  NAND2X0 U34297 ( .IN1(n30770), .IN2(n30769), .QN(n30771) );
  NAND4X0 U34298 ( .IN1(n34459), .IN2(n30773), .IN3(n30772), .IN4(n30771), 
        .QN(n30774) );
  NAND2X0 U34299 ( .IN1(n30775), .IN2(n30774), .QN(n30780) );
  OA222X1 U34300 ( .IN1(n30780), .IN2(n30777), .IN3(n30780), .IN4(n34389), 
        .IN5(\s4/msel/gnt_p1 [1]), .IN6(n30776), .Q(n30779) );
  AO21X1 U34301 ( .IN1(n30779), .IN2(n30778), .IN3(\s4/msel/gnt_p1 [2]), .Q(
        n30784) );
  AO221X1 U34302 ( .IN1(n34246), .IN2(n34459), .IN3(n34246), .IN4(n30781), 
        .IN5(n30780), .Q(n30783) );
  NAND3X0 U34303 ( .IN1(n30784), .IN2(n30783), .IN3(n30782), .QN(n17916) );
  NAND3X0 U34304 ( .IN1(n13627), .IN2(n13601), .IN3(m5s4_cyc), .QN(n30830) );
  NAND2X0 U34305 ( .IN1(n34232), .IN2(n30830), .QN(n30787) );
  NAND3X0 U34306 ( .IN1(n13575), .IN2(n13549), .IN3(m6s4_cyc), .QN(n30839) );
  NAND3X0 U34307 ( .IN1(n13523), .IN2(n13464), .IN3(m7s4_cyc), .QN(n30836) );
  NAND2X0 U34308 ( .IN1(n30839), .IN2(n30836), .QN(n30798) );
  OR2X1 U34309 ( .IN1(n30787), .IN2(n30798), .Q(n30785) );
  INVX0 U34310 ( .INP(n30836), .ZN(n30832) );
  NAND2X0 U34311 ( .IN1(n34232), .IN2(\s4/msel/gnt_p0 [0]), .QN(n30875) );
  INVX0 U34312 ( .INP(n30839), .ZN(n30851) );
  OR2X1 U34313 ( .IN1(n30875), .IN2(n30851), .Q(n30860) );
  NAND2X0 U34314 ( .IN1(\s4/msel/gnt_p0 [1]), .IN2(n30836), .QN(n30788) );
  OA21X1 U34315 ( .IN1(n30832), .IN2(n30860), .IN3(n30788), .Q(n30803) );
  NAND3X0 U34316 ( .IN1(n13679), .IN2(n13653), .IN3(m4s4_cyc), .QN(n30840) );
  INVX0 U34317 ( .INP(n30840), .ZN(n30858) );
  MUX21X1 U34318 ( .IN1(n30858), .IN2(n30851), .S(\s4/msel/gnt_p0 [1]), .Q(
        n30880) );
  NAND3X0 U34319 ( .IN1(n13888), .IN2(n13861), .IN3(m0s4_cyc), .QN(n30872) );
  INVX0 U34320 ( .INP(n30872), .ZN(n30849) );
  NAND3X0 U34321 ( .IN1(n13835), .IN2(n13809), .IN3(m1s4_cyc), .QN(n30876) );
  INVX0 U34322 ( .INP(n30876), .ZN(n30834) );
  NOR2X0 U34323 ( .IN1(n30849), .IN2(n30834), .QN(n30799) );
  NAND3X0 U34324 ( .IN1(n13783), .IN2(n13757), .IN3(m2s4_cyc), .QN(n30871) );
  NAND3X0 U34325 ( .IN1(n13731), .IN2(n13705), .IN3(m3s4_cyc), .QN(n30852) );
  NAND2X0 U34326 ( .IN1(n30871), .IN2(n30852), .QN(n30801) );
  INVX0 U34327 ( .INP(n30801), .ZN(n30807) );
  AO222X1 U34328 ( .IN1(n30785), .IN2(n30803), .IN3(n34378), .IN4(n30880), 
        .IN5(n30799), .IN6(n30807), .Q(n30786) );
  NAND2X0 U34329 ( .IN1(\s4/msel/gnt_p0 [2]), .IN2(n30786), .QN(n30797) );
  NAND4X0 U34330 ( .IN1(\s4/msel/gnt_p0 [2]), .IN2(\s4/msel/gnt_p0 [0]), .IN3(
        n30788), .IN4(n30787), .QN(n30882) );
  NAND2X0 U34331 ( .IN1(\s4/msel/gnt_p0 [0]), .IN2(\s4/msel/gnt_p0 [1]), .QN(
        n30792) );
  NOR2X0 U34332 ( .IN1(n30852), .IN2(n30792), .QN(n30873) );
  NOR2X0 U34333 ( .IN1(\s4/msel/gnt_p0 [2]), .IN2(n30873), .QN(n30790) );
  INVX0 U34334 ( .INP(n30871), .ZN(n30833) );
  NOR2X0 U34335 ( .IN1(\s4/msel/gnt_p0 [0]), .IN2(n34232), .QN(n30821) );
  NAND2X0 U34336 ( .IN1(n30833), .IN2(n30821), .QN(n30789) );
  NAND2X0 U34337 ( .IN1(n30790), .IN2(n30789), .QN(n30819) );
  MUX21X1 U34338 ( .IN1(n30872), .IN2(n30876), .S(\s4/msel/gnt_p0 [0]), .Q(
        n30820) );
  INVX0 U34339 ( .INP(n30830), .ZN(n30837) );
  NOR2X0 U34340 ( .IN1(n30837), .IN2(n30858), .QN(n30800) );
  INVX0 U34341 ( .INP(n30800), .ZN(n30806) );
  OAI22X1 U34342 ( .IN1(\s4/msel/gnt_p0 [1]), .IN2(n30820), .IN3(n30806), 
        .IN4(n30798), .QN(n30791) );
  NOR2X0 U34343 ( .IN1(n30819), .IN2(n30791), .QN(n30795) );
  INVX0 U34344 ( .INP(n30852), .ZN(n30813) );
  INVX0 U34345 ( .INP(n30821), .ZN(n30861) );
  OA21X1 U34346 ( .IN1(n30875), .IN2(n30833), .IN3(n30861), .Q(n30843) );
  NAND2X0 U34347 ( .IN1(n34378), .IN2(n34232), .QN(n30853) );
  OR2X1 U34348 ( .IN1(n30853), .IN2(n30834), .Q(n30805) );
  OA22X1 U34349 ( .IN1(n30813), .IN2(n30843), .IN3(n30805), .IN4(n30801), .Q(
        n30793) );
  NAND2X0 U34350 ( .IN1(n30793), .IN2(n30792), .QN(n30794) );
  NAND2X0 U34351 ( .IN1(n30795), .IN2(n30794), .QN(n30796) );
  NAND3X0 U34352 ( .IN1(n30797), .IN2(n30882), .IN3(n30796), .QN(n17915) );
  NOR2X0 U34353 ( .IN1(n30801), .IN2(n30798), .QN(n30808) );
  NOR2X0 U34354 ( .IN1(n30799), .IN2(n30798), .QN(n30812) );
  NOR2X0 U34355 ( .IN1(n30808), .IN2(n30812), .QN(n30804) );
  OA221X1 U34356 ( .IN1(n30801), .IN2(n30800), .IN3(n30801), .IN4(n30860), 
        .IN5(n30799), .Q(n30802) );
  OA22X1 U34357 ( .IN1(n30804), .IN2(n30853), .IN3(n30803), .IN4(n30802), .Q(
        n30818) );
  NAND2X0 U34358 ( .IN1(n30805), .IN2(n30875), .QN(n30811) );
  NAND2X0 U34359 ( .IN1(n30807), .IN2(n30806), .QN(n30810) );
  INVX0 U34360 ( .INP(n30808), .ZN(n30809) );
  NAND3X0 U34361 ( .IN1(n30811), .IN2(n30810), .IN3(n30809), .QN(n30816) );
  OR4X1 U34362 ( .IN1(n34232), .IN2(n30858), .IN3(n30837), .IN4(n30812), .Q(
        n30815) );
  NAND2X0 U34363 ( .IN1(n30813), .IN2(n30821), .QN(n30814) );
  NAND4X0 U34364 ( .IN1(n34457), .IN2(n30816), .IN3(n30815), .IN4(n30814), 
        .QN(n30817) );
  OA21X1 U34365 ( .IN1(n30818), .IN2(n34457), .IN3(n30817), .Q(n30829) );
  AO21X1 U34366 ( .IN1(n30829), .IN2(n30820), .IN3(n30819), .Q(n30828) );
  NAND2X0 U34367 ( .IN1(n30821), .IN2(n30851), .QN(n30826) );
  INVX0 U34368 ( .INP(n30829), .ZN(n30822) );
  NOR2X0 U34369 ( .IN1(n30837), .IN2(n30822), .QN(n30824) );
  NAND2X0 U34370 ( .IN1(n34378), .IN2(n30858), .QN(n30823) );
  NAND2X0 U34371 ( .IN1(n30824), .IN2(n30823), .QN(n30825) );
  NAND3X0 U34372 ( .IN1(n30826), .IN2(n30825), .IN3(\s4/msel/gnt_p0 [2]), .QN(
        n30827) );
  AO22X1 U34373 ( .IN1(\s4/msel/gnt_p0 [1]), .IN2(n30829), .IN3(n30828), .IN4(
        n30827), .Q(n17914) );
  OA21X1 U34374 ( .IN1(n30858), .IN2(n30830), .IN3(n30852), .Q(n30859) );
  NOR2X0 U34375 ( .IN1(n30851), .IN2(n30858), .QN(n30844) );
  NAND2X0 U34376 ( .IN1(\s4/msel/gnt_p0 [0]), .IN2(n30844), .QN(n30831) );
  OA221X1 U34377 ( .IN1(n30833), .IN2(n30859), .IN3(n30833), .IN4(n30831), 
        .IN5(n30876), .Q(n30848) );
  NAND2X0 U34378 ( .IN1(n30832), .IN2(n30844), .QN(n30846) );
  AO221X1 U34379 ( .IN1(n30848), .IN2(n30833), .IN3(n30848), .IN4(n30846), 
        .IN5(n30853), .Q(n30842) );
  NAND2X0 U34380 ( .IN1(n30871), .IN2(n30872), .QN(n30857) );
  NOR2X0 U34381 ( .IN1(n34378), .IN2(n30857), .QN(n30838) );
  NAND2X0 U34382 ( .IN1(n30834), .IN2(n30872), .QN(n30835) );
  NAND2X0 U34383 ( .IN1(n30836), .IN2(n30835), .QN(n30856) );
  AO221X1 U34384 ( .IN1(n30839), .IN2(n30838), .IN3(n30839), .IN4(n30856), 
        .IN5(n30837), .Q(n30850) );
  NAND3X0 U34385 ( .IN1(\s4/msel/gnt_p0 [1]), .IN2(n30840), .IN3(n30850), .QN(
        n30841) );
  NAND3X0 U34386 ( .IN1(n34457), .IN2(n30842), .IN3(n30841), .QN(n30870) );
  INVX0 U34387 ( .INP(n30843), .ZN(n30869) );
  NAND2X0 U34388 ( .IN1(n30876), .IN2(n34378), .QN(n30845) );
  NAND3X0 U34389 ( .IN1(n30845), .IN2(n30872), .IN3(n30844), .QN(n30847) );
  NAND3X0 U34390 ( .IN1(n30859), .IN2(n30847), .IN3(n30846), .QN(n30868) );
  OR3X1 U34391 ( .IN1(n34232), .IN2(n30849), .IN3(n30848), .Q(n30866) );
  INVX0 U34392 ( .INP(n30850), .ZN(n30855) );
  OR3X1 U34393 ( .IN1(n30857), .IN2(n30852), .IN3(n30851), .Q(n30854) );
  AO21X1 U34394 ( .IN1(n30855), .IN2(n30854), .IN3(n30853), .Q(n30865) );
  INVX0 U34395 ( .INP(n30856), .ZN(n30863) );
  AO22X1 U34396 ( .IN1(n30863), .IN2(n30862), .IN3(n30861), .IN4(n30860), .Q(
        n30864) );
  NAND4X0 U34397 ( .IN1(\s4/msel/gnt_p0 [2]), .IN2(n30866), .IN3(n30865), 
        .IN4(n30864), .QN(n30867) );
  OA221X1 U34398 ( .IN1(n30870), .IN2(n30869), .IN3(n30870), .IN4(n30868), 
        .IN5(n30867), .Q(n30878) );
  OA221X1 U34399 ( .IN1(\s4/msel/gnt_p0 [1]), .IN2(n30872), .IN3(n34232), 
        .IN4(n30871), .IN5(n30878), .Q(n30874) );
  NOR2X0 U34400 ( .IN1(n30874), .IN2(n30873), .QN(n30877) );
  AO221X1 U34401 ( .IN1(n30877), .IN2(n30876), .IN3(n30877), .IN4(n30875), 
        .IN5(\s4/msel/gnt_p0 [2]), .Q(n30883) );
  INVX0 U34402 ( .INP(n30878), .ZN(n30879) );
  AO221X1 U34403 ( .IN1(n34378), .IN2(n34457), .IN3(n34378), .IN4(n30880), 
        .IN5(n30879), .Q(n30881) );
  NAND3X0 U34404 ( .IN1(n30883), .IN2(n30882), .IN3(n30881), .QN(n17913) );
  NAND2X0 U34405 ( .IN1(n30884), .IN2(n30910), .QN(n30886) );
  OA221X1 U34406 ( .IN1(\s4/msel/gnt_p2 [1]), .IN2(n30927), .IN3(
        \s4/msel/gnt_p2 [1]), .IN4(n30945), .IN5(n30930), .Q(n30885) );
  NAND3X0 U34407 ( .IN1(\s4/msel/gnt_p2 [2]), .IN2(n30886), .IN3(n30885), .QN(
        n30895) );
  NOR2X0 U34408 ( .IN1(\s4/msel/gnt_p2 [0]), .IN2(\s4/msel/gnt_p2 [1]), .QN(
        n30953) );
  INVX0 U34409 ( .INP(n30953), .ZN(n30939) );
  NOR2X0 U34410 ( .IN1(\s4/msel/gnt_p2 [0]), .IN2(n34279), .QN(n30903) );
  NAND2X0 U34411 ( .IN1(n30949), .IN2(n30903), .QN(n30917) );
  OA21X1 U34412 ( .IN1(n30939), .IN2(n30900), .IN3(n30917), .Q(n30969) );
  INVX0 U34413 ( .INP(n30969), .ZN(n30894) );
  NOR2X0 U34414 ( .IN1(n34408), .IN2(n34279), .QN(n30899) );
  AND2X1 U34415 ( .IN1(n34279), .IN2(n30931), .Q(n30901) );
  AO22X1 U34416 ( .IN1(n30910), .IN2(n30901), .IN3(n30903), .IN4(n30926), .Q(
        n30887) );
  NOR2X0 U34417 ( .IN1(n30899), .IN2(n30887), .QN(n30892) );
  OR2X1 U34418 ( .IN1(n34408), .IN2(n30931), .Q(n30964) );
  OA21X1 U34419 ( .IN1(\s4/msel/gnt_p2 [0]), .IN2(n30941), .IN3(n30964), .Q(
        n30920) );
  NOR2X0 U34420 ( .IN1(\s4/msel/gnt_p2 [1]), .IN2(n30920), .QN(n30891) );
  NAND2X0 U34421 ( .IN1(n30928), .IN2(n30903), .QN(n30889) );
  NAND2X0 U34422 ( .IN1(n30899), .IN2(n30888), .QN(n30967) );
  NAND2X0 U34423 ( .IN1(n30889), .IN2(n30967), .QN(n30919) );
  NOR4X0 U34424 ( .IN1(n30892), .IN2(n30891), .IN3(n30890), .IN4(n30919), .QN(
        n30893) );
  AO222X1 U34425 ( .IN1(\s4/msel/gnt_p2 [2]), .IN2(n30895), .IN3(
        \s4/msel/gnt_p2 [2]), .IN4(n30894), .IN5(n30895), .IN6(n30893), .Q(
        n17912) );
  NAND2X0 U34426 ( .IN1(n30947), .IN2(n34408), .QN(n30916) );
  NAND4X0 U34427 ( .IN1(n30927), .IN2(n30941), .IN3(n30931), .IN4(n30900), 
        .QN(n30905) );
  NAND2X0 U34428 ( .IN1(n30930), .IN2(n30945), .QN(n30906) );
  NAND3X0 U34429 ( .IN1(n30927), .IN2(n30900), .IN3(n30906), .QN(n30896) );
  NAND3X0 U34430 ( .IN1(n30926), .IN2(n30905), .IN3(n30896), .QN(n30904) );
  NAND2X0 U34431 ( .IN1(n30910), .IN2(n30896), .QN(n30902) );
  INVX0 U34432 ( .INP(n30927), .ZN(n30942) );
  NOR2X0 U34433 ( .IN1(\s4/msel/gnt_p2 [1]), .IN2(n30928), .QN(n30935) );
  INVX0 U34434 ( .INP(n30906), .ZN(n30897) );
  OA21X1 U34435 ( .IN1(n30935), .IN2(n30909), .IN3(n30897), .Q(n30898) );
  NOR2X0 U34436 ( .IN1(n30942), .IN2(n30898), .QN(n30912) );
  AND2X1 U34437 ( .IN1(n30900), .IN2(n30899), .Q(n30959) );
  AO222X1 U34438 ( .IN1(n30904), .IN2(n30903), .IN3(n30902), .IN4(n30901), 
        .IN5(n30912), .IN6(n30959), .Q(n30915) );
  INVX0 U34439 ( .INP(n30905), .ZN(n30908) );
  NAND2X0 U34440 ( .IN1(\s4/msel/gnt_p2 [1]), .IN2(n30930), .QN(n30907) );
  OA22X1 U34441 ( .IN1(n30908), .IN2(n30907), .IN3(\s4/msel/gnt_p2 [1]), .IN4(
        n30906), .Q(n30913) );
  NOR2X0 U34442 ( .IN1(n30910), .IN2(n30909), .QN(n30911) );
  AO221X1 U34443 ( .IN1(n30913), .IN2(n30912), .IN3(n30913), .IN4(n30939), 
        .IN5(n30911), .Q(n30914) );
  MUX21X1 U34444 ( .IN1(n30915), .IN2(n30914), .S(\s4/msel/gnt_p2 [2]), .Q(
        n30921) );
  NAND3X0 U34445 ( .IN1(n30916), .IN2(n30921), .IN3(n30927), .QN(n30918) );
  NAND2X0 U34446 ( .IN1(n30918), .IN2(n30917), .QN(n30924) );
  AO21X1 U34447 ( .IN1(n30920), .IN2(n30921), .IN3(n30919), .Q(n30923) );
  AND2X1 U34448 ( .IN1(n30921), .IN2(\s4/msel/gnt_p2 [1]), .Q(n30922) );
  AO221X1 U34449 ( .IN1(\s4/msel/gnt_p2 [2]), .IN2(n30924), .IN3(n34607), 
        .IN4(n30923), .IN5(n30922), .Q(n17911) );
  INVX0 U34450 ( .INP(n30930), .ZN(n30925) );
  OA221X1 U34451 ( .IN1(\s4/msel/gnt_p2 [1]), .IN2(n30942), .IN3(n34279), 
        .IN4(n30925), .IN5(\s4/msel/gnt_p2 [0]), .Q(n30974) );
  NAND3X0 U34452 ( .IN1(n30961), .IN2(n30925), .IN3(n30933), .QN(n30929) );
  OA21X1 U34453 ( .IN1(n30947), .IN2(n30927), .IN3(n30926), .Q(n30948) );
  OA21X1 U34454 ( .IN1(n30928), .IN2(n30948), .IN3(n30931), .Q(n30952) );
  NAND2X0 U34455 ( .IN1(n30929), .IN2(n30952), .QN(n30940) );
  INVX0 U34456 ( .INP(n30941), .ZN(n30963) );
  OA21X1 U34457 ( .IN1(n30963), .IN2(n30931), .IN3(n30930), .Q(n30951) );
  INVX0 U34458 ( .INP(n30933), .ZN(n30932) );
  NOR2X0 U34459 ( .IN1(n30951), .IN2(n30932), .QN(n30937) );
  NAND3X0 U34460 ( .IN1(n30933), .IN2(\s4/msel/gnt_p2 [0]), .IN3(n30941), .QN(
        n30934) );
  NAND2X0 U34461 ( .IN1(n30934), .IN2(n30948), .QN(n30936) );
  OA22X1 U34462 ( .IN1(n30937), .IN2(n30936), .IN3(n30935), .IN4(n34408), .Q(
        n30938) );
  AO221X1 U34463 ( .IN1(n30953), .IN2(n30940), .IN3(n30939), .IN4(n30938), 
        .IN5(\s4/msel/gnt_p2 [2]), .Q(n30960) );
  NAND2X0 U34464 ( .IN1(n30961), .IN2(n30941), .QN(n30946) );
  NOR2X0 U34465 ( .IN1(n34408), .IN2(n30946), .QN(n30944) );
  INVX0 U34466 ( .INP(n30951), .ZN(n30943) );
  AO221X1 U34467 ( .IN1(n30945), .IN2(n30944), .IN3(n30945), .IN4(n30943), 
        .IN5(n30942), .Q(n30958) );
  AO221X1 U34468 ( .IN1(n30948), .IN2(n30947), .IN3(n30948), .IN4(n34408), 
        .IN5(n30946), .Q(n30950) );
  AO21X1 U34469 ( .IN1(n30951), .IN2(n30950), .IN3(n30949), .Q(n30956) );
  OR3X1 U34470 ( .IN1(n34279), .IN2(n30963), .IN3(n30952), .Q(n30955) );
  NAND2X0 U34471 ( .IN1(n30953), .IN2(n30958), .QN(n30954) );
  NAND4X0 U34472 ( .IN1(\s4/msel/gnt_p2 [2]), .IN2(n30956), .IN3(n30955), 
        .IN4(n30954), .QN(n30957) );
  OA221X1 U34473 ( .IN1(n30960), .IN2(n30959), .IN3(n30960), .IN4(n30958), 
        .IN5(n30957), .Q(n30968) );
  NAND3X0 U34474 ( .IN1(\s4/msel/gnt_p2 [1]), .IN2(n30968), .IN3(n30961), .QN(
        n30966) );
  INVX0 U34475 ( .INP(n30968), .ZN(n30962) );
  AO221X1 U34476 ( .IN1(n30964), .IN2(n30963), .IN3(n30964), .IN4(n30962), 
        .IN5(\s4/msel/gnt_p2 [1]), .Q(n30965) );
  NAND3X0 U34477 ( .IN1(n30967), .IN2(n30966), .IN3(n30965), .QN(n30973) );
  NOR2X0 U34478 ( .IN1(\s4/msel/gnt_p2 [0]), .IN2(\s4/msel/gnt_p2 [2]), .QN(
        n30971) );
  NAND2X0 U34479 ( .IN1(n30969), .IN2(n30968), .QN(n30970) );
  NOR2X0 U34480 ( .IN1(n30971), .IN2(n30970), .QN(n30972) );
  AO221X1 U34481 ( .IN1(\s4/msel/gnt_p2 [2]), .IN2(n30974), .IN3(n34607), 
        .IN4(n30973), .IN5(n30972), .Q(n17910) );
  NOR2X0 U34482 ( .IN1(n30975), .IN2(n34379), .QN(n30976) );
  MUX21X1 U34483 ( .IN1(n34344), .IN2(s15_data_o[0]), .S(n30976), .Q(n17909)
         );
  MUX21X1 U34484 ( .IN1(n34493), .IN2(s15_data_o[1]), .S(n30976), .Q(n17908)
         );
  MUX21X1 U34485 ( .IN1(n34343), .IN2(s15_data_o[2]), .S(n30976), .Q(n17907)
         );
  MUX21X1 U34486 ( .IN1(n34494), .IN2(s15_data_o[3]), .S(n30976), .Q(n17906)
         );
  MUX21X1 U34487 ( .IN1(n34587), .IN2(s15_data_o[4]), .S(n30976), .Q(n17905)
         );
  MUX21X1 U34488 ( .IN1(n34370), .IN2(s15_data_o[5]), .S(n30976), .Q(n17904)
         );
  MUX21X1 U34489 ( .IN1(n34317), .IN2(s15_data_o[6]), .S(n30976), .Q(n17903)
         );
  MUX21X1 U34490 ( .IN1(n34495), .IN2(s15_data_o[7]), .S(n30976), .Q(n17902)
         );
  MUX21X1 U34491 ( .IN1(n34235), .IN2(s15_data_o[8]), .S(n30976), .Q(n17901)
         );
  MUX21X1 U34492 ( .IN1(n34496), .IN2(s15_data_o[9]), .S(n30976), .Q(n17900)
         );
  MUX21X1 U34493 ( .IN1(n34342), .IN2(s15_data_o[10]), .S(n30976), .Q(n17899)
         );
  MUX21X1 U34494 ( .IN1(n34528), .IN2(s15_data_o[11]), .S(n30976), .Q(n17898)
         );
  MUX21X1 U34495 ( .IN1(n34341), .IN2(s15_data_o[12]), .S(n30976), .Q(n17897)
         );
  MUX21X1 U34496 ( .IN1(n34529), .IN2(s15_data_o[13]), .S(n30976), .Q(n17896)
         );
  MUX21X1 U34497 ( .IN1(n34316), .IN2(s15_data_o[14]), .S(n30976), .Q(n17895)
         );
  MUX21X1 U34498 ( .IN1(n34530), .IN2(s15_data_o[15]), .S(n30976), .Q(n17894)
         );
  INVX0 U34499 ( .INP(n31057), .ZN(n31020) );
  INVX0 U34500 ( .INP(n31021), .ZN(n31058) );
  MUX21X1 U34501 ( .IN1(n31020), .IN2(n31058), .S(\s5/msel/gnt_p3 [0]), .Q(
        n31006) );
  NOR2X0 U34502 ( .IN1(n34409), .IN2(n34227), .QN(n31043) );
  INVX0 U34503 ( .INP(n31043), .ZN(n31018) );
  OA221X1 U34504 ( .IN1(\s5/msel/gnt_p3 [1]), .IN2(n31006), .IN3(n34227), 
        .IN4(n30977), .IN5(n31018), .Q(n30981) );
  INVX0 U34505 ( .INP(n30991), .ZN(n30979) );
  NOR2X0 U34506 ( .IN1(\s5/msel/gnt_p3 [0]), .IN2(\s5/msel/gnt_p3 [1]), .QN(
        n31017) );
  NAND2X0 U34507 ( .IN1(n31017), .IN2(n31021), .QN(n30990) );
  NAND2X0 U34508 ( .IN1(\s5/msel/gnt_p3 [1]), .IN2(n31036), .QN(n30978) );
  OA221X1 U34509 ( .IN1(n30979), .IN2(n34409), .IN3(n30979), .IN4(n30990), 
        .IN5(n30978), .Q(n30980) );
  NOR3X0 U34510 ( .IN1(n30982), .IN2(n30981), .IN3(n30980), .QN(n30988) );
  NOR2X0 U34511 ( .IN1(\s5/msel/gnt_p3 [1]), .IN2(n31008), .QN(n31033) );
  NOR2X0 U34512 ( .IN1(n31007), .IN2(n31033), .QN(n30999) );
  NAND2X0 U34513 ( .IN1(n30983), .IN2(n30991), .QN(n30986) );
  INVX0 U34514 ( .INP(n31023), .ZN(n31029) );
  NAND2X0 U34515 ( .IN1(n31029), .IN2(n34227), .QN(n31055) );
  NOR2X0 U34516 ( .IN1(n34409), .IN2(n34275), .QN(n31063) );
  INVX0 U34517 ( .INP(n31063), .ZN(n30984) );
  INVX0 U34518 ( .INP(n31038), .ZN(n31022) );
  AO221X1 U34519 ( .IN1(\s5/msel/gnt_p3 [1]), .IN2(n31046), .IN3(n34227), 
        .IN4(n31022), .IN5(n34275), .Q(n31015) );
  NAND2X0 U34520 ( .IN1(n30984), .IN2(n31015), .QN(n30985) );
  NAND4X0 U34521 ( .IN1(n30999), .IN2(n30986), .IN3(n31055), .IN4(n30985), 
        .QN(n30987) );
  OA21X1 U34522 ( .IN1(\s5/msel/gnt_p3 [2]), .IN2(n30988), .IN3(n30987), .Q(
        n17893) );
  OA21X1 U34523 ( .IN1(n31008), .IN2(n30992), .IN3(n30991), .Q(n30993) );
  OA222X1 U34524 ( .IN1(n34227), .IN2(n31001), .IN3(n31019), .IN4(n31058), 
        .IN5(n30997), .IN6(n31017), .Q(n30989) );
  OA22X1 U34525 ( .IN1(n30993), .IN2(n30990), .IN3(n30989), .IN4(n30992), .Q(
        n31005) );
  INVX0 U34526 ( .INP(n31017), .ZN(n31044) );
  NAND2X0 U34527 ( .IN1(n31018), .IN2(n31044), .QN(n31032) );
  OR2X1 U34528 ( .IN1(n31032), .IN2(n30991), .Q(n31004) );
  NAND2X0 U34529 ( .IN1(n34409), .IN2(n31023), .QN(n31037) );
  NOR2X0 U34530 ( .IN1(n31036), .IN2(n31037), .QN(n30996) );
  OA22X1 U34531 ( .IN1(n30993), .IN2(n31018), .IN3(n34227), .IN4(n30992), .Q(
        n30994) );
  NAND2X0 U34532 ( .IN1(n31004), .IN2(n30994), .QN(n30995) );
  NOR2X0 U34533 ( .IN1(n30996), .IN2(n30995), .QN(n31002) );
  OA21X1 U34534 ( .IN1(n31001), .IN2(n31053), .IN3(n30997), .Q(n30998) );
  OA22X1 U34535 ( .IN1(n30999), .IN2(n31032), .IN3(n30998), .IN4(n31037), .Q(
        n31000) );
  OA21X1 U34536 ( .IN1(n31002), .IN2(n31001), .IN3(n31000), .Q(n31003) );
  OA222X1 U34537 ( .IN1(\s5/msel/gnt_p3 [2]), .IN2(n31005), .IN3(
        \s5/msel/gnt_p3 [2]), .IN4(n31004), .IN5(n31003), .IN6(n34275), .Q(
        n31009) );
  OR2X1 U34538 ( .IN1(n34227), .IN2(n31009), .Q(n31014) );
  NAND2X0 U34539 ( .IN1(n31016), .IN2(n31043), .QN(n31061) );
  AO221X1 U34540 ( .IN1(n31061), .IN2(n31009), .IN3(n31061), .IN4(n31006), 
        .IN5(\s5/msel/gnt_p3 [2]), .Q(n31013) );
  NAND2X0 U34541 ( .IN1(\s5/msel/gnt_p3 [1]), .IN2(n31007), .QN(n31056) );
  OA21X1 U34542 ( .IN1(n31029), .IN2(n31009), .IN3(n31056), .Q(n31011) );
  OA22X1 U34543 ( .IN1(n31022), .IN2(n31009), .IN3(n34227), .IN4(n31008), .Q(
        n31010) );
  AO221X1 U34544 ( .IN1(\s5/msel/gnt_p3 [0]), .IN2(n31011), .IN3(n34409), 
        .IN4(n31010), .IN5(n34275), .Q(n31012) );
  NAND3X0 U34545 ( .IN1(n31014), .IN2(n31013), .IN3(n31012), .QN(n17892) );
  NAND2X0 U34546 ( .IN1(n34409), .IN2(n31015), .QN(n31066) );
  OA21X1 U34547 ( .IN1(n31046), .IN2(n34409), .IN3(n31023), .Q(n31047) );
  NOR2X0 U34548 ( .IN1(n31022), .IN2(n31047), .QN(n31028) );
  AO221X1 U34549 ( .IN1(n31053), .IN2(n31016), .IN3(n31053), .IN4(n31028), 
        .IN5(n31058), .Q(n31042) );
  NAND2X0 U34550 ( .IN1(n31017), .IN2(n31042), .QN(n31027) );
  NOR2X0 U34551 ( .IN1(n31022), .IN2(n31018), .QN(n31025) );
  OA21X1 U34552 ( .IN1(n31021), .IN2(n31020), .IN3(n31019), .Q(n31034) );
  OR3X1 U34553 ( .IN1(n31046), .IN2(n31022), .IN3(n31034), .Q(n31031) );
  NAND2X0 U34554 ( .IN1(n31031), .IN2(n31023), .QN(n31024) );
  NAND2X0 U34555 ( .IN1(n31025), .IN2(n31024), .QN(n31026) );
  NAND3X0 U34556 ( .IN1(n31027), .IN2(n34275), .IN3(n31026), .QN(n31054) );
  OAI21X1 U34557 ( .IN1(n31057), .IN2(n31029), .IN3(n31028), .QN(n31030) );
  NAND3X0 U34558 ( .IN1(n31036), .IN2(n31031), .IN3(n31030), .QN(n31052) );
  NOR2X0 U34559 ( .IN1(n31033), .IN2(n31032), .QN(n31041) );
  NAND2X0 U34560 ( .IN1(n31057), .IN2(n31053), .QN(n31035) );
  OA21X1 U34561 ( .IN1(n31036), .IN2(n31035), .IN3(n31034), .Q(n31045) );
  NAND4X0 U34562 ( .IN1(n31038), .IN2(n31057), .IN3(n31037), .IN4(n31053), 
        .QN(n31039) );
  NAND2X0 U34563 ( .IN1(n31045), .IN2(n31039), .QN(n31040) );
  NAND2X0 U34564 ( .IN1(n31041), .IN2(n31040), .QN(n31050) );
  NAND3X0 U34565 ( .IN1(n31043), .IN2(n31057), .IN3(n31042), .QN(n31049) );
  AO221X1 U34566 ( .IN1(n31047), .IN2(n31046), .IN3(n31047), .IN4(n31045), 
        .IN5(n31044), .Q(n31048) );
  NAND4X0 U34567 ( .IN1(\s5/msel/gnt_p3 [2]), .IN2(n31050), .IN3(n31049), 
        .IN4(n31048), .QN(n31051) );
  OA221X1 U34568 ( .IN1(n31054), .IN2(n31053), .IN3(n31054), .IN4(n31052), 
        .IN5(n31051), .Q(n31065) );
  NAND2X0 U34569 ( .IN1(n31056), .IN2(n31055), .QN(n31064) );
  OAI21X1 U34570 ( .IN1(n31057), .IN2(\s5/msel/gnt_p3 [1]), .IN3(n31065), .QN(
        n31060) );
  NAND3X0 U34571 ( .IN1(\s5/msel/gnt_p3 [0]), .IN2(n31058), .IN3(n34227), .QN(
        n31059) );
  NAND3X0 U34572 ( .IN1(n31061), .IN2(n31060), .IN3(n31059), .QN(n31062) );
  AO222X1 U34573 ( .IN1(n31066), .IN2(n31065), .IN3(n31064), .IN4(n31063), 
        .IN5(n31062), .IN6(n34275), .Q(n17891) );
  NAND3X0 U34574 ( .IN1(n13550), .IN2(m6s5_cyc), .IN3(n34341), .QN(n31116) );
  NAND3X0 U34575 ( .IN1(n13465), .IN2(m7s5_cyc), .IN3(n34316), .QN(n31120) );
  NAND2X0 U34576 ( .IN1(n31116), .IN2(n31120), .QN(n31092) );
  NAND3X0 U34577 ( .IN1(n13602), .IN2(m5s5_cyc), .IN3(n34342), .QN(n31126) );
  NAND2X0 U34578 ( .IN1(n34252), .IN2(n31126), .QN(n31071) );
  NAND2X0 U34579 ( .IN1(\s5/msel/gnt_p1 [1]), .IN2(n31120), .QN(n31072) );
  AO22X1 U34580 ( .IN1(n34657), .IN2(n31072), .IN3(n34252), .IN4(n31092), .Q(
        n31097) );
  OA21X1 U34581 ( .IN1(n31092), .IN2(n31071), .IN3(n31097), .Q(n31067) );
  NAND3X0 U34582 ( .IN1(n13810), .IN2(m1s5_cyc), .IN3(n34343), .QN(n31148) );
  NAND3X0 U34583 ( .IN1(n13862), .IN2(m0s5_cyc), .IN3(n34344), .QN(n31144) );
  NAND2X0 U34584 ( .IN1(n31148), .IN2(n31144), .QN(n31091) );
  AND3X1 U34585 ( .IN1(n13758), .IN2(m2s5_cyc), .IN3(n34587), .Q(n31128) );
  NAND3X0 U34586 ( .IN1(n13706), .IN2(m3s5_cyc), .IN3(n34317), .QN(n31130) );
  INVX0 U34587 ( .INP(n31130), .ZN(n31118) );
  NOR2X0 U34588 ( .IN1(n31128), .IN2(n31118), .QN(n31088) );
  INVX0 U34589 ( .INP(n31088), .ZN(n31093) );
  NOR2X0 U34590 ( .IN1(n31091), .IN2(n31093), .QN(n34108) );
  NOR2X0 U34591 ( .IN1(n31067), .IN2(n34108), .QN(n31069) );
  NAND3X0 U34592 ( .IN1(n13654), .IN2(m4s5_cyc), .IN3(n34235), .QN(n31115) );
  INVX0 U34593 ( .INP(n31115), .ZN(n31129) );
  INVX0 U34594 ( .INP(n31116), .ZN(n31137) );
  MUX21X1 U34595 ( .IN1(n31129), .IN2(n31137), .S(\s5/msel/gnt_p1 [1]), .Q(
        n31156) );
  NAND2X0 U34596 ( .IN1(n34657), .IN2(n31156), .QN(n31068) );
  NAND2X0 U34597 ( .IN1(n31069), .IN2(n31068), .QN(n31070) );
  NAND2X0 U34598 ( .IN1(\s5/msel/gnt_p1 [2]), .IN2(n31070), .QN(n31079) );
  NAND4X0 U34599 ( .IN1(\s5/msel/gnt_p1 [2]), .IN2(\s5/msel/gnt_p1 [0]), .IN3(
        n31072), .IN4(n31071), .QN(n31157) );
  AND2X1 U34600 ( .IN1(n34252), .IN2(n31148), .Q(n31085) );
  NAND2X0 U34601 ( .IN1(n31088), .IN2(n31085), .QN(n31073) );
  OA21X1 U34602 ( .IN1(n31118), .IN2(n34252), .IN3(n31073), .Q(n31077) );
  NAND2X0 U34603 ( .IN1(n31115), .IN2(n31126), .QN(n31089) );
  NOR2X0 U34604 ( .IN1(n31092), .IN2(n31089), .QN(n34109) );
  MUX21X1 U34605 ( .IN1(n31144), .IN2(n31148), .S(\s5/msel/gnt_p1 [0]), .Q(
        n31102) );
  NOR2X0 U34606 ( .IN1(\s5/msel/gnt_p1 [1]), .IN2(n31102), .QN(n31076) );
  NAND2X0 U34607 ( .IN1(\s5/msel/gnt_p1 [0]), .IN2(\s5/msel/gnt_p1 [1]), .QN(
        n31104) );
  NOR2X0 U34608 ( .IN1(n31130), .IN2(n31104), .QN(n31147) );
  NOR2X0 U34609 ( .IN1(\s5/msel/gnt_p1 [2]), .IN2(n31147), .QN(n31075) );
  NOR2X0 U34610 ( .IN1(\s5/msel/gnt_p1 [0]), .IN2(n34252), .QN(n31103) );
  NAND2X0 U34611 ( .IN1(n31128), .IN2(n31103), .QN(n31074) );
  NAND2X0 U34612 ( .IN1(n31075), .IN2(n31074), .QN(n31101) );
  OR4X1 U34613 ( .IN1(n31077), .IN2(n34109), .IN3(n31076), .IN4(n31101), .Q(
        n31078) );
  NAND3X0 U34614 ( .IN1(n31079), .IN2(n31157), .IN3(n31078), .QN(n17890) );
  INVX0 U34615 ( .INP(n31092), .ZN(n31080) );
  AO21X1 U34616 ( .IN1(n34252), .IN2(n31080), .IN3(n31089), .Q(n31082) );
  INVX0 U34617 ( .INP(n31082), .ZN(n31081) );
  NAND2X0 U34618 ( .IN1(n31080), .IN2(n31091), .QN(n31083) );
  AO21X1 U34619 ( .IN1(n31081), .IN2(n31083), .IN3(n31118), .Q(n31087) );
  NAND2X0 U34620 ( .IN1(n31088), .IN2(n31082), .QN(n31086) );
  NOR2X0 U34621 ( .IN1(n31129), .IN2(n31104), .QN(n31142) );
  NAND2X0 U34622 ( .IN1(n31126), .IN2(n31083), .QN(n31094) );
  INVX0 U34623 ( .INP(n31094), .ZN(n31084) );
  AO222X1 U34624 ( .IN1(n31087), .IN2(n31103), .IN3(n31086), .IN4(n31085), 
        .IN5(n31142), .IN6(n31084), .Q(n31100) );
  NOR2X0 U34625 ( .IN1(\s5/msel/gnt_p1 [1]), .IN2(n34657), .QN(n31150) );
  OA21X1 U34626 ( .IN1(n31150), .IN2(n31089), .IN3(n31088), .Q(n31090) );
  NOR2X0 U34627 ( .IN1(n31091), .IN2(n31090), .QN(n31098) );
  NOR2X0 U34628 ( .IN1(n31093), .IN2(n31092), .QN(n31095) );
  NOR2X0 U34629 ( .IN1(n31095), .IN2(n31094), .QN(n31096) );
  NAND2X0 U34630 ( .IN1(n34657), .IN2(n34252), .QN(n31134) );
  OA22X1 U34631 ( .IN1(n31098), .IN2(n31097), .IN3(n31096), .IN4(n31134), .Q(
        n31099) );
  MUX21X1 U34632 ( .IN1(n31100), .IN2(n31099), .S(\s5/msel/gnt_p1 [2]), .Q(
        n31114) );
  AO21X1 U34633 ( .IN1(n31114), .IN2(n31102), .IN3(n31101), .Q(n31113) );
  INVX0 U34634 ( .INP(n31103), .ZN(n31105) );
  OA22X1 U34635 ( .IN1(n31116), .IN2(n31105), .IN3(n31120), .IN4(n31104), .Q(
        n31111) );
  INVX0 U34636 ( .INP(n31114), .ZN(n31107) );
  INVX0 U34637 ( .INP(n31126), .ZN(n31106) );
  NOR2X0 U34638 ( .IN1(n31107), .IN2(n31106), .QN(n31109) );
  NAND2X0 U34639 ( .IN1(n34657), .IN2(n31129), .QN(n31108) );
  NAND2X0 U34640 ( .IN1(n31109), .IN2(n31108), .QN(n31110) );
  NAND3X0 U34641 ( .IN1(\s5/msel/gnt_p1 [2]), .IN2(n31111), .IN3(n31110), .QN(
        n31112) );
  AO22X1 U34642 ( .IN1(\s5/msel/gnt_p1 [1]), .IN2(n31114), .IN3(n31113), .IN4(
        n31112), .Q(n17889) );
  NOR2X0 U34643 ( .IN1(n31128), .IN2(n34252), .QN(n31145) );
  NAND2X0 U34644 ( .IN1(n31116), .IN2(n31115), .QN(n31121) );
  NOR2X0 U34645 ( .IN1(n31129), .IN2(n31126), .QN(n31117) );
  NOR2X0 U34646 ( .IN1(n31118), .IN2(n31117), .QN(n31119) );
  OA21X1 U34647 ( .IN1(n34657), .IN2(n31121), .IN3(n31119), .Q(n31123) );
  INVX0 U34648 ( .INP(n31144), .ZN(n31133) );
  AND2X1 U34649 ( .IN1(n31133), .IN2(n31119), .Q(n31122) );
  OA21X1 U34650 ( .IN1(n31133), .IN2(n31148), .IN3(n31120), .Q(n31131) );
  OA22X1 U34651 ( .IN1(n31123), .IN2(n31122), .IN3(n31131), .IN4(n31121), .Q(
        n31124) );
  OA21X1 U34652 ( .IN1(n31128), .IN2(n31123), .IN3(n31148), .Q(n31127) );
  OA22X1 U34653 ( .IN1(n31128), .IN2(n31124), .IN3(n31127), .IN4(n31134), .Q(
        n31125) );
  NAND2X0 U34654 ( .IN1(n31125), .IN2(n34371), .QN(n31143) );
  OA21X1 U34655 ( .IN1(n31137), .IN2(n31131), .IN3(n31126), .Q(n31135) );
  INVX0 U34656 ( .INP(n31135), .ZN(n31141) );
  OR3X1 U34657 ( .IN1(n34252), .IN2(n31133), .IN3(n31127), .Q(n31139) );
  AO221X1 U34658 ( .IN1(n31130), .IN2(n31129), .IN3(n31130), .IN4(n34657), 
        .IN5(n31128), .Q(n31132) );
  OA21X1 U34659 ( .IN1(n31133), .IN2(n31132), .IN3(n31131), .Q(n31136) );
  OA22X1 U34660 ( .IN1(n31137), .IN2(n31136), .IN3(n31135), .IN4(n31134), .Q(
        n31138) );
  NAND3X0 U34661 ( .IN1(\s5/msel/gnt_p1 [2]), .IN2(n31139), .IN3(n31138), .QN(
        n31140) );
  OA221X1 U34662 ( .IN1(n31143), .IN2(n31142), .IN3(n31143), .IN4(n31141), 
        .IN5(n31140), .Q(n31154) );
  OA21X1 U34663 ( .IN1(n31145), .IN2(n31144), .IN3(n31154), .Q(n31146) );
  NOR2X0 U34664 ( .IN1(n31147), .IN2(n31146), .QN(n31152) );
  INVX0 U34665 ( .INP(n31148), .ZN(n31149) );
  NAND2X0 U34666 ( .IN1(n31150), .IN2(n31149), .QN(n31151) );
  NAND2X0 U34667 ( .IN1(n31152), .IN2(n31151), .QN(n31153) );
  NAND2X0 U34668 ( .IN1(n31153), .IN2(n34371), .QN(n31159) );
  INVX0 U34669 ( .INP(n31154), .ZN(n31155) );
  AO221X1 U34670 ( .IN1(n34657), .IN2(n34371), .IN3(n34657), .IN4(n31156), 
        .IN5(n31155), .Q(n31158) );
  NAND3X0 U34671 ( .IN1(n31159), .IN2(n31158), .IN3(n31157), .QN(n17888) );
  NAND3X0 U34672 ( .IN1(n13628), .IN2(n13602), .IN3(m5s5_cyc), .QN(n31202) );
  NAND2X0 U34673 ( .IN1(n34415), .IN2(n31202), .QN(n31162) );
  NAND3X0 U34674 ( .IN1(n13576), .IN2(n13550), .IN3(m6s5_cyc), .QN(n31216) );
  NAND3X0 U34675 ( .IN1(n13524), .IN2(n13465), .IN3(m7s5_cyc), .QN(n31205) );
  NAND2X0 U34676 ( .IN1(n31216), .IN2(n31205), .QN(n31178) );
  OR2X1 U34677 ( .IN1(n31162), .IN2(n31178), .Q(n31160) );
  NAND2X0 U34678 ( .IN1(\s5/msel/gnt_p0 [1]), .IN2(n31205), .QN(n31163) );
  OA21X1 U34679 ( .IN1(n34398), .IN2(n31178), .IN3(n31163), .Q(n31184) );
  NAND3X0 U34680 ( .IN1(n13680), .IN2(n13654), .IN3(m4s5_cyc), .QN(n31215) );
  INVX0 U34681 ( .INP(n31215), .ZN(n31217) );
  INVX0 U34682 ( .INP(n31216), .ZN(n31218) );
  MUX21X1 U34683 ( .IN1(n31217), .IN2(n31218), .S(\s5/msel/gnt_p0 [1]), .Q(
        n31244) );
  NAND3X0 U34684 ( .IN1(n13890), .IN2(n13862), .IN3(m0s5_cyc), .QN(n31237) );
  INVX0 U34685 ( .INP(n31237), .ZN(n31204) );
  NAND3X0 U34686 ( .IN1(n13836), .IN2(n13810), .IN3(m1s5_cyc), .QN(n31203) );
  INVX0 U34687 ( .INP(n31203), .ZN(n31167) );
  NOR2X0 U34688 ( .IN1(n31204), .IN2(n31167), .QN(n31183) );
  NAND3X0 U34689 ( .IN1(n13784), .IN2(n13758), .IN3(m2s5_cyc), .QN(n31236) );
  INVX0 U34690 ( .INP(n31236), .ZN(n31227) );
  NAND3X0 U34691 ( .IN1(n13732), .IN2(n13706), .IN3(m3s5_cyc), .QN(n31201) );
  INVX0 U34692 ( .INP(n31201), .ZN(n31180) );
  NOR2X0 U34693 ( .IN1(n31227), .IN2(n31180), .QN(n31175) );
  AO222X1 U34694 ( .IN1(n31160), .IN2(n31184), .IN3(n34398), .IN4(n31244), 
        .IN5(n31183), .IN6(n31175), .Q(n31161) );
  NAND2X0 U34695 ( .IN1(\s5/msel/gnt_p0 [2]), .IN2(n31161), .QN(n31173) );
  NAND4X0 U34696 ( .IN1(\s5/msel/gnt_p0 [2]), .IN2(\s5/msel/gnt_p0 [0]), .IN3(
        n31163), .IN4(n31162), .QN(n31246) );
  NAND2X0 U34697 ( .IN1(\s5/msel/gnt_p0 [0]), .IN2(\s5/msel/gnt_p0 [1]), .QN(
        n31168) );
  NOR2X0 U34698 ( .IN1(n31201), .IN2(n31168), .QN(n31238) );
  NOR2X0 U34699 ( .IN1(\s5/msel/gnt_p0 [2]), .IN2(n31238), .QN(n31165) );
  NOR2X0 U34700 ( .IN1(\s5/msel/gnt_p0 [0]), .IN2(n34415), .QN(n31195) );
  NAND2X0 U34701 ( .IN1(n31227), .IN2(n31195), .QN(n31164) );
  NAND2X0 U34702 ( .IN1(n31165), .IN2(n31164), .QN(n31190) );
  NAND2X0 U34703 ( .IN1(\s5/msel/gnt_p0 [0]), .IN2(n31167), .QN(n31240) );
  OA21X1 U34704 ( .IN1(\s5/msel/gnt_p0 [0]), .IN2(n31237), .IN3(n31240), .Q(
        n31191) );
  NAND2X0 U34705 ( .IN1(n31202), .IN2(n31215), .QN(n31174) );
  OAI22X1 U34706 ( .IN1(\s5/msel/gnt_p0 [1]), .IN2(n31191), .IN3(n31174), 
        .IN4(n31178), .QN(n31166) );
  NOR2X0 U34707 ( .IN1(n31190), .IN2(n31166), .QN(n31171) );
  NOR2X0 U34708 ( .IN1(\s5/msel/gnt_p0 [0]), .IN2(\s5/msel/gnt_p0 [1]), .QN(
        n31234) );
  INVX0 U34709 ( .INP(n31234), .ZN(n31225) );
  NOR2X0 U34710 ( .IN1(n31167), .IN2(n31225), .QN(n31176) );
  NOR2X0 U34711 ( .IN1(\s5/msel/gnt_p0 [1]), .IN2(n34398), .QN(n31177) );
  AO21X1 U34712 ( .IN1(n31177), .IN2(n31236), .IN3(n31195), .Q(n31224) );
  AOI22X1 U34713 ( .IN1(n31176), .IN2(n31175), .IN3(n31201), .IN4(n31224), 
        .QN(n31169) );
  NAND2X0 U34714 ( .IN1(n31169), .IN2(n31168), .QN(n31170) );
  NAND2X0 U34715 ( .IN1(n31171), .IN2(n31170), .QN(n31172) );
  NAND3X0 U34716 ( .IN1(n31173), .IN2(n31246), .IN3(n31172), .QN(n17887) );
  INVX0 U34717 ( .INP(n31202), .ZN(n31212) );
  NOR2X0 U34718 ( .IN1(n31183), .IN2(n31178), .QN(n31185) );
  NOR4X0 U34719 ( .IN1(n31217), .IN2(n31212), .IN3(n31185), .IN4(n34415), .QN(
        n31189) );
  NAND2X0 U34720 ( .IN1(n31175), .IN2(n31174), .QN(n31182) );
  OA21X1 U34721 ( .IN1(n31177), .IN2(n31176), .IN3(n31182), .Q(n31179) );
  OR4X1 U34722 ( .IN1(n31178), .IN2(\s5/msel/gnt_p0 [1]), .IN3(n31227), .IN4(
        n31180), .Q(n31181) );
  AO22X1 U34723 ( .IN1(n31180), .IN2(n31195), .IN3(n31179), .IN4(n31181), .Q(
        n31188) );
  OA221X1 U34724 ( .IN1(n31184), .IN2(n31183), .IN3(n31184), .IN4(n31182), 
        .IN5(n31181), .Q(n31187) );
  INVX0 U34725 ( .INP(n31185), .ZN(n31186) );
  AO222X1 U34726 ( .IN1(n34258), .IN2(n31189), .IN3(n34258), .IN4(n31188), 
        .IN5(n18198), .IN6(\s5/msel/gnt_p0 [2]), .Q(n31200) );
  AO21X1 U34727 ( .IN1(n31191), .IN2(n31200), .IN3(n31190), .Q(n31199) );
  NOR2X0 U34728 ( .IN1(\s5/msel/gnt_p0 [0]), .IN2(n31215), .QN(n31193) );
  NAND2X0 U34729 ( .IN1(n31200), .IN2(n31202), .QN(n31192) );
  NOR2X0 U34730 ( .IN1(n31193), .IN2(n31192), .QN(n31194) );
  NOR2X0 U34731 ( .IN1(n31194), .IN2(n34258), .QN(n31197) );
  NAND2X0 U34732 ( .IN1(n31218), .IN2(n31195), .QN(n31196) );
  NAND2X0 U34733 ( .IN1(n31197), .IN2(n31196), .QN(n31198) );
  AO22X1 U34734 ( .IN1(\s5/msel/gnt_p0 [1]), .IN2(n31200), .IN3(n31199), .IN4(
        n31198), .Q(n17886) );
  OA21X1 U34735 ( .IN1(n31202), .IN2(n31217), .IN3(n31201), .Q(n31222) );
  OA21X1 U34736 ( .IN1(n31227), .IN2(n31222), .IN3(n31203), .Q(n31228) );
  OR3X1 U34737 ( .IN1(n34415), .IN2(n31204), .IN3(n31228), .Q(n31209) );
  NOR2X0 U34738 ( .IN1(n31204), .IN2(n31203), .QN(n31206) );
  INVX0 U34739 ( .INP(n31205), .ZN(n31220) );
  NOR2X0 U34740 ( .IN1(n31206), .IN2(n31220), .QN(n31211) );
  NAND2X0 U34741 ( .IN1(n31236), .IN2(n31237), .QN(n31210) );
  AO221X1 U34742 ( .IN1(n31222), .IN2(n31217), .IN3(n31222), .IN4(n34398), 
        .IN5(n31210), .Q(n31207) );
  AO21X1 U34743 ( .IN1(n31211), .IN2(n31207), .IN3(n31218), .Q(n31208) );
  NAND3X0 U34744 ( .IN1(\s5/msel/gnt_p0 [2]), .IN2(n31209), .IN3(n31208), .QN(
        n31235) );
  NOR2X0 U34745 ( .IN1(n34398), .IN2(n31210), .QN(n31214) );
  INVX0 U34746 ( .INP(n31211), .ZN(n31213) );
  AO221X1 U34747 ( .IN1(n31216), .IN2(n31214), .IN3(n31216), .IN4(n31213), 
        .IN5(n31212), .Q(n31233) );
  NAND3X0 U34748 ( .IN1(\s5/msel/gnt_p0 [1]), .IN2(n31215), .IN3(n31233), .QN(
        n31231) );
  NAND4X0 U34749 ( .IN1(\s5/msel/gnt_p0 [0]), .IN2(n31216), .IN3(n31237), 
        .IN4(n31215), .QN(n31221) );
  NOR2X0 U34750 ( .IN1(n31218), .IN2(n31217), .QN(n31219) );
  NAND2X0 U34751 ( .IN1(n31220), .IN2(n31219), .QN(n31226) );
  NAND3X0 U34752 ( .IN1(n31222), .IN2(n31221), .IN3(n31226), .QN(n31223) );
  NAND2X0 U34753 ( .IN1(n31224), .IN2(n31223), .QN(n31230) );
  AO221X1 U34754 ( .IN1(n31228), .IN2(n31227), .IN3(n31228), .IN4(n31226), 
        .IN5(n31225), .Q(n31229) );
  NAND4X0 U34755 ( .IN1(n34258), .IN2(n31231), .IN3(n31230), .IN4(n31229), 
        .QN(n31232) );
  OA221X1 U34756 ( .IN1(n31235), .IN2(n31234), .IN3(n31235), .IN4(n31233), 
        .IN5(n31232), .Q(n31242) );
  OA221X1 U34757 ( .IN1(\s5/msel/gnt_p0 [1]), .IN2(n31237), .IN3(n34415), 
        .IN4(n31236), .IN5(n31242), .Q(n31239) );
  NOR2X0 U34758 ( .IN1(n31239), .IN2(n31238), .QN(n31241) );
  AO221X1 U34759 ( .IN1(n31241), .IN2(\s5/msel/gnt_p0 [1]), .IN3(n31241), 
        .IN4(n31240), .IN5(\s5/msel/gnt_p0 [2]), .Q(n31247) );
  INVX0 U34760 ( .INP(n31242), .ZN(n31243) );
  AO221X1 U34761 ( .IN1(n34398), .IN2(n31244), .IN3(n34398), .IN4(n34258), 
        .IN5(n31243), .Q(n31245) );
  NAND3X0 U34762 ( .IN1(n31247), .IN2(n31246), .IN3(n31245), .QN(n17885) );
  INVX0 U34763 ( .INP(n31297), .ZN(n31306) );
  INVX0 U34764 ( .INP(n31273), .ZN(n31308) );
  MUX21X1 U34765 ( .IN1(n31306), .IN2(n31308), .S(\s5/msel/gnt_p2 [1]), .Q(
        n31328) );
  NAND2X0 U34766 ( .IN1(\s5/msel/gnt_p2 [1]), .IN2(n31287), .QN(n31326) );
  INVX0 U34767 ( .INP(n31248), .ZN(n31261) );
  NAND2X0 U34768 ( .IN1(n31324), .IN2(n31261), .QN(n31249) );
  AO22X1 U34769 ( .IN1(n34256), .IN2(n31328), .IN3(n31326), .IN4(n31249), .Q(
        n31255) );
  NOR2X0 U34770 ( .IN1(n34256), .IN2(n34396), .QN(n31296) );
  NAND2X0 U34771 ( .IN1(n31251), .IN2(n31296), .QN(n31320) );
  NAND3X0 U34772 ( .IN1(\s5/msel/gnt_p2 [1]), .IN2(n31285), .IN3(n34256), .QN(
        n31250) );
  NAND3X0 U34773 ( .IN1(n34426), .IN2(n31320), .IN3(n31250), .QN(n31277) );
  INVX0 U34774 ( .INP(n31294), .ZN(n31316) );
  INVX0 U34775 ( .INP(n31288), .ZN(n31283) );
  MUX21X1 U34776 ( .IN1(n31316), .IN2(n31283), .S(\s5/msel/gnt_p2 [0]), .Q(
        n31275) );
  NAND2X0 U34777 ( .IN1(n31256), .IN2(n31288), .QN(n31252) );
  AO221X1 U34778 ( .IN1(n34396), .IN2(n31275), .IN3(n34396), .IN4(n31252), 
        .IN5(n31251), .Q(n31253) );
  NOR3X0 U34779 ( .IN1(n34106), .IN2(n31277), .IN3(n31253), .QN(n31254) );
  AO221X1 U34780 ( .IN1(\s5/msel/gnt_p2 [2]), .IN2(n34105), .IN3(
        \s5/msel/gnt_p2 [2]), .IN4(n31255), .IN5(n31254), .Q(n17884) );
  NOR2X0 U34781 ( .IN1(n31256), .IN2(n31257), .QN(n31259) );
  NOR2X0 U34782 ( .IN1(n31257), .IN2(n31260), .QN(n31263) );
  NOR2X0 U34783 ( .IN1(\s5/msel/gnt_p2 [1]), .IN2(n31285), .QN(n31291) );
  OAI21X1 U34784 ( .IN1(n31291), .IN2(n31257), .IN3(n31261), .QN(n31267) );
  OA21X1 U34785 ( .IN1(n31263), .IN2(n31326), .IN3(n31267), .Q(n31258) );
  NOR2X0 U34786 ( .IN1(\s5/msel/gnt_p2 [0]), .IN2(\s5/msel/gnt_p2 [1]), .QN(
        n31304) );
  INVX0 U34787 ( .INP(n31304), .ZN(n31300) );
  OA22X1 U34788 ( .IN1(n31259), .IN2(n31258), .IN3(n31324), .IN4(n31300), .Q(
        n31272) );
  OA21X1 U34789 ( .IN1(n31261), .IN2(n31260), .IN3(n31284), .Q(n31265) );
  NAND2X0 U34790 ( .IN1(n31265), .IN2(n31318), .QN(n31262) );
  NAND3X0 U34791 ( .IN1(n31288), .IN2(n31262), .IN3(n34396), .QN(n31270) );
  INVX0 U34792 ( .INP(n31263), .ZN(n31264) );
  NAND2X0 U34793 ( .IN1(n31265), .IN2(n31264), .QN(n31266) );
  NAND2X0 U34794 ( .IN1(\s5/msel/gnt_p2 [1]), .IN2(n31266), .QN(n31269) );
  NAND4X0 U34795 ( .IN1(n31296), .IN2(n31297), .IN3(n31324), .IN4(n31267), 
        .QN(n31268) );
  NAND4X0 U34796 ( .IN1(n31270), .IN2(n34426), .IN3(n31269), .IN4(n31268), 
        .QN(n31271) );
  OA21X1 U34797 ( .IN1(n31272), .IN2(n34426), .IN3(n31271), .Q(n31282) );
  AND3X1 U34798 ( .IN1(\s5/msel/gnt_p2 [2]), .IN2(\s5/msel/gnt_p2 [0]), .IN3(
        n31324), .Q(n31281) );
  INVX0 U34799 ( .INP(n31282), .ZN(n31276) );
  OA22X1 U34800 ( .IN1(n31306), .IN2(n31276), .IN3(n34396), .IN4(n31273), .Q(
        n31274) );
  NOR2X0 U34801 ( .IN1(\s5/msel/gnt_p2 [0]), .IN2(n31274), .QN(n31279) );
  NOR2X0 U34802 ( .IN1(n31276), .IN2(n31275), .QN(n31278) );
  OA22X1 U34803 ( .IN1(n31279), .IN2(n34426), .IN3(n31278), .IN4(n31277), .Q(
        n31280) );
  AO221X1 U34804 ( .IN1(n31282), .IN2(\s5/msel/gnt_p2 [1]), .IN3(n31282), 
        .IN4(n31281), .IN5(n31280), .Q(n17883) );
  NAND2X0 U34805 ( .IN1(\s5/msel/gnt_p2 [0]), .IN2(n31283), .QN(n31317) );
  OA21X1 U34806 ( .IN1(n31306), .IN2(n31324), .IN3(n31284), .Q(n31307) );
  OA21X1 U34807 ( .IN1(n31285), .IN2(n31307), .IN3(n31288), .Q(n31302) );
  OR4X1 U34808 ( .IN1(n31287), .IN2(n31285), .IN3(n31308), .IN4(n31306), .Q(
        n31286) );
  NAND2X0 U34809 ( .IN1(n31302), .IN2(n31286), .QN(n31301) );
  OA21X1 U34810 ( .IN1(n31288), .IN2(n31316), .IN3(n31287), .Q(n31310) );
  INVX0 U34811 ( .INP(n31310), .ZN(n31290) );
  NOR2X0 U34812 ( .IN1(n31308), .IN2(n31306), .QN(n31289) );
  OA221X1 U34813 ( .IN1(n31290), .IN2(\s5/msel/gnt_p2 [0]), .IN3(n31290), 
        .IN4(n31294), .IN5(n31289), .Q(n31293) );
  INVX0 U34814 ( .INP(n31307), .ZN(n31292) );
  OA22X1 U34815 ( .IN1(n31293), .IN2(n31292), .IN3(n31291), .IN4(n34256), .Q(
        n31299) );
  NAND2X0 U34816 ( .IN1(n31318), .IN2(n31294), .QN(n31305) );
  OR2X1 U34817 ( .IN1(n34256), .IN2(n31305), .Q(n31295) );
  OAI221X1 U34818 ( .IN1(n31308), .IN2(n31310), .IN3(n31308), .IN4(n31295), 
        .IN5(n31324), .QN(n31303) );
  AND3X1 U34819 ( .IN1(n31303), .IN2(n31297), .IN3(n31296), .Q(n31298) );
  AO221X1 U34820 ( .IN1(n31304), .IN2(n31301), .IN3(n31300), .IN4(n31299), 
        .IN5(n31298), .Q(n31315) );
  OR3X1 U34821 ( .IN1(n34396), .IN2(n31316), .IN3(n31302), .Q(n31313) );
  NAND2X0 U34822 ( .IN1(n31304), .IN2(n31303), .QN(n31312) );
  AO221X1 U34823 ( .IN1(n31307), .IN2(n31306), .IN3(n31307), .IN4(n34256), 
        .IN5(n31305), .Q(n31309) );
  AO21X1 U34824 ( .IN1(n31310), .IN2(n31309), .IN3(n31308), .Q(n31311) );
  NAND4X0 U34825 ( .IN1(\s5/msel/gnt_p2 [2]), .IN2(n31313), .IN3(n31312), 
        .IN4(n31311), .QN(n31314) );
  OA21X1 U34826 ( .IN1(\s5/msel/gnt_p2 [2]), .IN2(n31315), .IN3(n31314), .Q(
        n31319) );
  INVX0 U34827 ( .INP(n31319), .ZN(n31327) );
  AO221X1 U34828 ( .IN1(n31317), .IN2(n31316), .IN3(n31317), .IN4(n31327), 
        .IN5(\s5/msel/gnt_p2 [1]), .Q(n31322) );
  NAND3X0 U34829 ( .IN1(\s5/msel/gnt_p2 [1]), .IN2(n31319), .IN3(n31318), .QN(
        n31321) );
  NAND3X0 U34830 ( .IN1(n31322), .IN2(n31321), .IN3(n31320), .QN(n31323) );
  NAND2X0 U34831 ( .IN1(n31323), .IN2(n34426), .QN(n31331) );
  NAND2X0 U34832 ( .IN1(n34396), .IN2(n31324), .QN(n31325) );
  NAND4X0 U34833 ( .IN1(\s5/msel/gnt_p2 [2]), .IN2(\s5/msel/gnt_p2 [0]), .IN3(
        n31326), .IN4(n31325), .QN(n31330) );
  AO221X1 U34834 ( .IN1(n34256), .IN2(n34426), .IN3(n34256), .IN4(n31328), 
        .IN5(n31327), .Q(n31329) );
  NAND3X0 U34835 ( .IN1(n31331), .IN2(n31330), .IN3(n31329), .QN(n17882) );
  NOR2X0 U34836 ( .IN1(n31332), .IN2(n34379), .QN(n31333) );
  MUX21X1 U34837 ( .IN1(n34629), .IN2(s15_data_o[0]), .S(n31333), .Q(n17881)
         );
  MUX21X1 U34838 ( .IN1(n34579), .IN2(s15_data_o[1]), .S(n31333), .Q(n17880)
         );
  MUX21X1 U34839 ( .IN1(n34237), .IN2(s15_data_o[2]), .S(n31333), .Q(n17879)
         );
  MUX21X1 U34840 ( .IN1(n34368), .IN2(s15_data_o[3]), .S(n31333), .Q(n17878)
         );
  MUX21X1 U34841 ( .IN1(n34362), .IN2(s15_data_o[4]), .S(n31333), .Q(n17877)
         );
  MUX21X1 U34842 ( .IN1(n34552), .IN2(s15_data_o[5]), .S(n31333), .Q(n17876)
         );
  MUX21X1 U34843 ( .IN1(n34346), .IN2(s15_data_o[6]), .S(n31333), .Q(n17875)
         );
  MUX21X1 U34844 ( .IN1(n34532), .IN2(s15_data_o[7]), .S(n31333), .Q(n17874)
         );
  MUX21X1 U34845 ( .IN1(n34630), .IN2(s15_data_o[8]), .S(n31333), .Q(n17873)
         );
  MUX21X1 U34846 ( .IN1(n34566), .IN2(s15_data_o[9]), .S(n31333), .Q(n17872)
         );
  MUX21X1 U34847 ( .IN1(n34345), .IN2(s15_data_o[10]), .S(n31333), .Q(n17871)
         );
  MUX21X1 U34848 ( .IN1(n34531), .IN2(s15_data_o[11]), .S(n31333), .Q(n17870)
         );
  MUX21X1 U34849 ( .IN1(n34366), .IN2(s15_data_o[12]), .S(n31333), .Q(n17869)
         );
  MUX21X1 U34850 ( .IN1(n34599), .IN2(s15_data_o[13]), .S(n31333), .Q(n17868)
         );
  MUX21X1 U34851 ( .IN1(n34628), .IN2(s15_data_o[14]), .S(n31333), .Q(n17867)
         );
  MUX21X1 U34852 ( .IN1(n34565), .IN2(s15_data_o[15]), .S(n31333), .Q(n17866)
         );
  NAND2X0 U34853 ( .IN1(m4s6_cyc), .IN2(n34566), .QN(n31334) );
  NOR2X0 U34854 ( .IN1(n13681), .IN2(n31334), .QN(n31405) );
  INVX0 U34855 ( .INP(n31405), .ZN(n31391) );
  NAND3X0 U34856 ( .IN1(m6s6_cyc), .IN2(n34366), .IN3(n34599), .QN(n31390) );
  OA221X1 U34857 ( .IN1(\s6/msel/gnt_p3 [1]), .IN2(n31391), .IN3(n34270), 
        .IN4(n31390), .IN5(\s6/msel/gnt_p3 [2]), .Q(n31422) );
  INVX0 U34858 ( .INP(n31390), .ZN(n31386) );
  NAND2X0 U34859 ( .IN1(m7s6_cyc), .IN2(n34565), .QN(n31335) );
  NOR2X0 U34860 ( .IN1(n13525), .IN2(n31335), .QN(n31358) );
  NOR2X0 U34861 ( .IN1(n31386), .IN2(n31358), .QN(n31367) );
  NOR2X0 U34862 ( .IN1(\s6/msel/gnt_p3 [1]), .IN2(n31367), .QN(n31337) );
  NAND2X0 U34863 ( .IN1(\s6/msel/gnt_p3 [0]), .IN2(\s6/msel/gnt_p3 [2]), .QN(
        n31435) );
  NOR2X0 U34864 ( .IN1(n31337), .IN2(n31435), .QN(n31350) );
  NOR2X0 U34865 ( .IN1(n31422), .IN2(n31350), .QN(n31341) );
  NAND2X0 U34866 ( .IN1(m0s6_cyc), .IN2(n34579), .QN(n31336) );
  NOR2X0 U34867 ( .IN1(n13892), .IN2(n31336), .QN(n31425) );
  NAND3X0 U34868 ( .IN1(m1s6_cyc), .IN2(n34237), .IN3(n34368), .QN(n31394) );
  INVX0 U34869 ( .INP(n31394), .ZN(n31423) );
  NOR2X0 U34870 ( .IN1(n31425), .IN2(n31423), .QN(n34115) );
  NAND3X0 U34871 ( .IN1(m2s6_cyc), .IN2(n34362), .IN3(n34552), .QN(n31409) );
  NAND3X0 U34872 ( .IN1(m3s6_cyc), .IN2(n34346), .IN3(n34532), .QN(n31392) );
  NAND2X0 U34873 ( .IN1(n31409), .IN2(n31392), .QN(n31351) );
  INVX0 U34874 ( .INP(n31351), .ZN(n34114) );
  NAND2X0 U34875 ( .IN1(n34115), .IN2(n34114), .QN(n31339) );
  INVX0 U34876 ( .INP(n31337), .ZN(n31338) );
  NAND2X0 U34877 ( .IN1(n31339), .IN2(n31338), .QN(n31340) );
  NOR2X0 U34878 ( .IN1(n31341), .IN2(n31340), .QN(n31349) );
  NAND3X0 U34879 ( .IN1(m5s6_cyc), .IN2(n34345), .IN3(n34531), .QN(n31393) );
  NAND2X0 U34880 ( .IN1(\s6/msel/gnt_p3 [1]), .IN2(n31358), .QN(n31376) );
  OA21X1 U34881 ( .IN1(\s6/msel/gnt_p3 [1]), .IN2(n31393), .IN3(n31376), .Q(
        n31434) );
  NOR2X0 U34882 ( .IN1(n34449), .IN2(n34270), .QN(n31372) );
  INVX0 U34883 ( .INP(n31372), .ZN(n31403) );
  INVX0 U34884 ( .INP(n31392), .ZN(n31384) );
  MUX21X1 U34885 ( .IN1(n31425), .IN2(n31423), .S(\s6/msel/gnt_p3 [0]), .Q(
        n31373) );
  NOR2X0 U34886 ( .IN1(\s6/msel/gnt_p3 [0]), .IN2(n34270), .QN(n31400) );
  INVX0 U34887 ( .INP(n31400), .ZN(n31342) );
  INVX0 U34888 ( .INP(n31409), .ZN(n31426) );
  OA222X1 U34889 ( .IN1(n31403), .IN2(n31384), .IN3(n31373), .IN4(
        \s6/msel/gnt_p3 [1]), .IN5(n31342), .IN6(n31426), .Q(n31343) );
  INVX0 U34890 ( .INP(n31393), .ZN(n31375) );
  NOR2X0 U34891 ( .IN1(n31405), .IN2(n31375), .QN(n31361) );
  AND2X1 U34892 ( .IN1(n31361), .IN2(n31367), .Q(n34113) );
  NOR2X0 U34893 ( .IN1(n31343), .IN2(n34113), .QN(n31347) );
  NOR2X0 U34894 ( .IN1(n31426), .IN2(n34449), .QN(n31414) );
  NOR2X0 U34895 ( .IN1(n31400), .IN2(n31414), .QN(n31344) );
  OA22X1 U34896 ( .IN1(n31384), .IN2(n31344), .IN3(n31423), .IN4(n31351), .Q(
        n31345) );
  NAND2X0 U34897 ( .IN1(n31345), .IN2(n31403), .QN(n31346) );
  NAND2X0 U34898 ( .IN1(n31347), .IN2(n31346), .QN(n31348) );
  AOI22X1 U34899 ( .IN1(n31349), .IN2(n31434), .IN3(n34640), .IN4(n31348), 
        .QN(n17865) );
  NOR2X0 U34900 ( .IN1(\s6/msel/gnt_p3 [0]), .IN2(n34640), .QN(n31369) );
  NOR2X0 U34901 ( .IN1(n31369), .IN2(n31350), .QN(n31355) );
  INVX0 U34902 ( .INP(n31425), .ZN(n31396) );
  NAND2X0 U34903 ( .IN1(n34270), .IN2(n31390), .QN(n31382) );
  AO21X1 U34904 ( .IN1(n31361), .IN2(n31382), .IN3(n31351), .Q(n31357) );
  NAND2X0 U34905 ( .IN1(n34449), .IN2(n31393), .QN(n31380) );
  NOR2X0 U34906 ( .IN1(\s6/msel/gnt_p3 [0]), .IN2(\s6/msel/gnt_p3 [1]), .QN(
        n31408) );
  INVX0 U34907 ( .INP(n31408), .ZN(n31388) );
  NAND3X0 U34908 ( .IN1(n31403), .IN2(n31388), .IN3(n31351), .QN(n31356) );
  NAND3X0 U34909 ( .IN1(n31403), .IN2(n31380), .IN3(n31356), .QN(n31352) );
  NAND4X0 U34910 ( .IN1(n31396), .IN2(n31394), .IN3(n31357), .IN4(n31352), 
        .QN(n31353) );
  NAND2X0 U34911 ( .IN1(n31353), .IN2(n31376), .QN(n31354) );
  NOR2X0 U34912 ( .IN1(n31355), .IN2(n31354), .QN(n31368) );
  INVX0 U34913 ( .INP(n31356), .ZN(n31365) );
  AND3X1 U34914 ( .IN1(n31408), .IN2(n31394), .IN3(n31357), .Q(n31364) );
  NAND2X0 U34915 ( .IN1(n31372), .IN2(n31396), .QN(n31419) );
  INVX0 U34916 ( .INP(n31358), .ZN(n31406) );
  NAND2X0 U34917 ( .IN1(n31419), .IN2(n31406), .QN(n31360) );
  INVX0 U34918 ( .INP(n31367), .ZN(n31359) );
  AO22X1 U34919 ( .IN1(n31394), .IN2(n31360), .IN3(n31388), .IN4(n31359), .Q(
        n31362) );
  OA221X1 U34920 ( .IN1(n31362), .IN2(n34115), .IN3(n31362), .IN4(n31400), 
        .IN5(n31361), .Q(n31363) );
  NOR4X0 U34921 ( .IN1(\s6/msel/gnt_p3 [2]), .IN2(n31365), .IN3(n31364), .IN4(
        n31363), .QN(n31366) );
  AO221X1 U34922 ( .IN1(n31368), .IN2(n31367), .IN3(n31368), .IN4(n31380), 
        .IN5(n31366), .Q(n31374) );
  OA22X1 U34923 ( .IN1(n31405), .IN2(n31374), .IN3(n34270), .IN4(n31390), .Q(
        n31371) );
  INVX0 U34924 ( .INP(n31369), .ZN(n31370) );
  OA22X1 U34925 ( .IN1(n31371), .IN2(n31370), .IN3(n34270), .IN4(n31374), .Q(
        n31379) );
  NAND2X0 U34926 ( .IN1(n31384), .IN2(n31372), .QN(n31427) );
  AO221X1 U34927 ( .IN1(n31427), .IN2(n31373), .IN3(n31427), .IN4(n31374), 
        .IN5(\s6/msel/gnt_p3 [2]), .Q(n31378) );
  NAND3X0 U34928 ( .IN1(n31379), .IN2(n31378), .IN3(n31377), .QN(n17864) );
  OA21X1 U34929 ( .IN1(n31425), .IN2(n31394), .IN3(n31406), .Q(n31399) );
  NOR2X0 U34930 ( .IN1(n31426), .IN2(n31425), .QN(n31383) );
  OAI221X1 U34931 ( .IN1(n31384), .IN2(n31391), .IN3(n31384), .IN4(n31380), 
        .IN5(n31383), .QN(n31381) );
  AO22X1 U34932 ( .IN1(\s6/msel/gnt_p3 [0]), .IN2(n31382), .IN3(n31399), .IN4(
        n31381), .Q(n31389) );
  NAND2X0 U34933 ( .IN1(n31384), .IN2(n31383), .QN(n31385) );
  OA21X1 U34934 ( .IN1(n31386), .IN2(n31399), .IN3(n31393), .Q(n31404) );
  OA21X1 U34935 ( .IN1(n31386), .IN2(n31385), .IN3(n31404), .Q(n31387) );
  OA221X1 U34936 ( .IN1(n31408), .IN2(n31389), .IN3(n31388), .IN4(n31387), 
        .IN5(\s6/msel/gnt_p3 [2]), .Q(n31421) );
  NAND2X0 U34937 ( .IN1(n31391), .IN2(n31390), .QN(n31407) );
  OA21X1 U34938 ( .IN1(n31405), .IN2(n31393), .IN3(n31392), .Q(n31397) );
  OA21X1 U34939 ( .IN1(n34449), .IN2(n31407), .IN3(n31397), .Q(n31395) );
  OA21X1 U34940 ( .IN1(n31426), .IN2(n31395), .IN3(n31394), .Q(n31420) );
  INVX0 U34941 ( .INP(n31407), .ZN(n31402) );
  NAND3X0 U34942 ( .IN1(n31402), .IN2(\s6/msel/gnt_p3 [0]), .IN3(n31396), .QN(
        n31398) );
  NAND2X0 U34943 ( .IN1(n31398), .IN2(n31397), .QN(n31413) );
  INVX0 U34944 ( .INP(n31399), .ZN(n31401) );
  OA221X1 U34945 ( .IN1(n31413), .IN2(n31402), .IN3(n31413), .IN4(n31401), 
        .IN5(n31400), .Q(n31417) );
  NOR3X0 U34946 ( .IN1(n31405), .IN2(n31404), .IN3(n31403), .QN(n31416) );
  NOR2X0 U34947 ( .IN1(n31407), .IN2(n31406), .QN(n31412) );
  INVX0 U34948 ( .INP(n31420), .ZN(n31410) );
  OA221X1 U34949 ( .IN1(n31410), .IN2(n31412), .IN3(n31410), .IN4(n31409), 
        .IN5(n31408), .Q(n31411) );
  AO221X1 U34950 ( .IN1(n31414), .IN2(n31413), .IN3(n31414), .IN4(n31412), 
        .IN5(n31411), .Q(n31415) );
  NOR4X0 U34951 ( .IN1(\s6/msel/gnt_p3 [2]), .IN2(n31417), .IN3(n31416), .IN4(
        n31415), .QN(n31418) );
  AO221X1 U34952 ( .IN1(n31421), .IN2(n31420), .IN3(n31421), .IN4(n31419), 
        .IN5(n31418), .Q(n31433) );
  NOR2X0 U34953 ( .IN1(\s6/msel/gnt_p3 [0]), .IN2(n31422), .QN(n31432) );
  NAND2X0 U34954 ( .IN1(\s6/msel/gnt_p3 [0]), .IN2(n31423), .QN(n31424) );
  NOR2X0 U34955 ( .IN1(n31424), .IN2(\s6/msel/gnt_p3 [1]), .QN(n31430) );
  AO221X1 U34956 ( .IN1(\s6/msel/gnt_p3 [1]), .IN2(n31426), .IN3(n34270), 
        .IN4(n31425), .IN5(n31433), .Q(n31428) );
  NAND2X0 U34957 ( .IN1(n31428), .IN2(n31427), .QN(n31429) );
  NOR2X0 U34958 ( .IN1(n31430), .IN2(n31429), .QN(n31431) );
  OAI222X1 U34959 ( .IN1(n31435), .IN2(n31434), .IN3(n31433), .IN4(n31432), 
        .IN5(n31431), .IN6(\s6/msel/gnt_p3 [2]), .QN(n17863) );
  NAND3X0 U34960 ( .IN1(n13469), .IN2(m7s6_cyc), .IN3(n34628), .QN(n31468) );
  NAND2X0 U34961 ( .IN1(\s6/msel/gnt_p1 [1]), .IN2(n31468), .QN(n31493) );
  NAND3X0 U34962 ( .IN1(n13603), .IN2(m5s6_cyc), .IN3(n34345), .QN(n31469) );
  NAND2X0 U34963 ( .IN1(n34666), .IN2(n31469), .QN(n31494) );
  NAND3X0 U34964 ( .IN1(n13551), .IN2(m6s6_cyc), .IN3(n34366), .QN(n31436) );
  NAND2X0 U34965 ( .IN1(n31436), .IN2(n31468), .QN(n31448) );
  NAND3X0 U34966 ( .IN1(n13759), .IN2(m2s6_cyc), .IN3(n34362), .QN(n31467) );
  INVX0 U34967 ( .INP(n31467), .ZN(n31483) );
  NAND3X0 U34968 ( .IN1(n13707), .IN2(m3s6_cyc), .IN3(n34346), .QN(n31496) );
  INVX0 U34969 ( .INP(n31496), .ZN(n31439) );
  NOR2X0 U34970 ( .IN1(n31483), .IN2(n31439), .QN(n34120) );
  NAND3X0 U34971 ( .IN1(n13863), .IN2(m0s6_cyc), .IN3(n34629), .QN(n31497) );
  NAND3X0 U34972 ( .IN1(n13811), .IN2(m1s6_cyc), .IN3(n34237), .QN(n31495) );
  NAND2X0 U34973 ( .IN1(n31497), .IN2(n31495), .QN(n31453) );
  INVX0 U34974 ( .INP(n31453), .ZN(n34121) );
  NAND3X0 U34975 ( .IN1(n13655), .IN2(m4s6_cyc), .IN3(n34630), .QN(n31449) );
  INVX0 U34976 ( .INP(n31449), .ZN(n31485) );
  INVX0 U34977 ( .INP(n31436), .ZN(n31480) );
  MUX21X1 U34978 ( .IN1(n31485), .IN2(n31480), .S(\s6/msel/gnt_p1 [1]), .Q(
        n31492) );
  AO22X1 U34979 ( .IN1(n34120), .IN2(n34121), .IN3(n34243), .IN4(n31492), .Q(
        n31437) );
  AO221X1 U34980 ( .IN1(n31493), .IN2(n31494), .IN3(n31493), .IN4(n31448), 
        .IN5(n31437), .Q(n31444) );
  MUX21X1 U34981 ( .IN1(n31497), .IN2(n31495), .S(\s6/msel/gnt_p1 [0]), .Q(
        n31460) );
  NAND2X0 U34982 ( .IN1(n34666), .IN2(n31495), .QN(n31446) );
  INVX0 U34983 ( .INP(n34120), .ZN(n31438) );
  OAI22X1 U34984 ( .IN1(n31439), .IN2(n34666), .IN3(n31446), .IN4(n31438), 
        .QN(n31440) );
  OA21X1 U34985 ( .IN1(n31460), .IN2(\s6/msel/gnt_p1 [1]), .IN3(n31440), .Q(
        n31443) );
  NAND2X0 U34986 ( .IN1(n31449), .IN2(n31469), .QN(n31452) );
  NOR2X0 U34987 ( .IN1(n31448), .IN2(n31452), .QN(n34119) );
  AO221X1 U34988 ( .IN1(\s6/msel/gnt_p1 [0]), .IN2(n31496), .IN3(n34243), 
        .IN4(n31467), .IN5(n34666), .Q(n31441) );
  NAND2X0 U34989 ( .IN1(n31441), .IN2(n34597), .QN(n31459) );
  NOR2X0 U34990 ( .IN1(n34119), .IN2(n31459), .QN(n31442) );
  AO22X1 U34991 ( .IN1(\s6/msel/gnt_p1 [2]), .IN2(n31444), .IN3(n31443), .IN4(
        n31442), .Q(n17862) );
  INVX0 U34992 ( .INP(n31448), .ZN(n31445) );
  OA21X1 U34993 ( .IN1(n31445), .IN2(n31452), .IN3(n34120), .Q(n31447) );
  OA22X1 U34994 ( .IN1(n31447), .IN2(n31446), .IN3(n31496), .IN4(n34666), .Q(
        n31451) );
  AO21X1 U34995 ( .IN1(\s6/msel/gnt_p1 [1]), .IN2(n34121), .IN3(n31448), .Q(
        n31456) );
  NAND4X0 U34996 ( .IN1(\s6/msel/gnt_p1 [1]), .IN2(n31469), .IN3(n31449), 
        .IN4(n31456), .QN(n31450) );
  NAND2X0 U34997 ( .IN1(n31451), .IN2(n31450), .QN(n31458) );
  NOR2X0 U34998 ( .IN1(n31453), .IN2(n31452), .QN(n31455) );
  NOR2X0 U34999 ( .IN1(n34120), .IN2(n31453), .QN(n31454) );
  AO221X1 U35000 ( .IN1(n31456), .IN2(n31455), .IN3(n31456), .IN4(n31493), 
        .IN5(n31454), .Q(n31457) );
  MUX21X1 U35001 ( .IN1(n31458), .IN2(n31457), .S(\s6/msel/gnt_p1 [2]), .Q(
        n31466) );
  AO21X1 U35002 ( .IN1(n31460), .IN2(n31466), .IN3(n31459), .Q(n31465) );
  NAND2X0 U35003 ( .IN1(n31485), .IN2(n34243), .QN(n31461) );
  NAND3X0 U35004 ( .IN1(n31461), .IN2(n31466), .IN3(n31469), .QN(n31463) );
  NAND3X0 U35005 ( .IN1(\s6/msel/gnt_p1 [1]), .IN2(n31480), .IN3(n34243), .QN(
        n31462) );
  NAND3X0 U35006 ( .IN1(\s6/msel/gnt_p1 [2]), .IN2(n31463), .IN3(n31462), .QN(
        n31464) );
  AO22X1 U35007 ( .IN1(\s6/msel/gnt_p1 [1]), .IN2(n31466), .IN3(n31465), .IN4(
        n31464), .Q(n17861) );
  OA21X1 U35008 ( .IN1(n31485), .IN2(n31469), .IN3(n31496), .Q(n31486) );
  OAI21X1 U35009 ( .IN1(n31483), .IN2(n31486), .IN3(n31495), .QN(n31478) );
  NAND3X0 U35010 ( .IN1(\s6/msel/gnt_p1 [1]), .IN2(n31478), .IN3(n31497), .QN(
        n31475) );
  NAND2X0 U35011 ( .IN1(n31467), .IN2(n31497), .QN(n31470) );
  INVX0 U35012 ( .INP(n31497), .ZN(n31481) );
  OA21X1 U35013 ( .IN1(n31481), .IN2(n31495), .IN3(n31468), .Q(n31482) );
  OA21X1 U35014 ( .IN1(n34243), .IN2(n31470), .IN3(n31482), .Q(n31472) );
  OA21X1 U35015 ( .IN1(n31480), .IN2(n31472), .IN3(n31469), .Q(n31476) );
  NAND2X0 U35016 ( .IN1(n34243), .IN2(n34666), .QN(n31477) );
  AND2X1 U35017 ( .IN1(n31485), .IN2(n31482), .Q(n31471) );
  OA22X1 U35018 ( .IN1(n31472), .IN2(n31471), .IN3(n31486), .IN4(n31470), .Q(
        n31473) );
  OA22X1 U35019 ( .IN1(n31476), .IN2(n31477), .IN3(n31480), .IN4(n31473), .Q(
        n31474) );
  NAND3X0 U35020 ( .IN1(n31475), .IN2(n31474), .IN3(\s6/msel/gnt_p1 [2]), .QN(
        n31491) );
  OR4X1 U35021 ( .IN1(n34666), .IN2(n34243), .IN3(n31485), .IN4(n31476), .Q(
        n31489) );
  INVX0 U35022 ( .INP(n31477), .ZN(n31479) );
  NAND2X0 U35023 ( .IN1(n31479), .IN2(n31478), .QN(n31488) );
  AO221X1 U35024 ( .IN1(n31482), .IN2(n31481), .IN3(n31482), .IN4(n34243), 
        .IN5(n31480), .Q(n31484) );
  AO221X1 U35025 ( .IN1(n31486), .IN2(n31485), .IN3(n31486), .IN4(n31484), 
        .IN5(n31483), .Q(n31487) );
  NAND4X0 U35026 ( .IN1(n34597), .IN2(n31489), .IN3(n31488), .IN4(n31487), 
        .QN(n31490) );
  NAND2X0 U35027 ( .IN1(n31491), .IN2(n31490), .QN(n31498) );
  AO221X1 U35028 ( .IN1(n34243), .IN2(n34597), .IN3(n34243), .IN4(n31492), 
        .IN5(n31498), .Q(n31503) );
  NAND4X0 U35029 ( .IN1(\s6/msel/gnt_p1 [2]), .IN2(\s6/msel/gnt_p1 [0]), .IN3(
        n31494), .IN4(n31493), .QN(n31502) );
  AO221X1 U35030 ( .IN1(\s6/msel/gnt_p1 [1]), .IN2(n31496), .IN3(n34666), 
        .IN4(n31495), .IN5(n34243), .Q(n31500) );
  NOR2X0 U35031 ( .IN1(\s6/msel/gnt_p1 [1]), .IN2(n31497), .QN(n31499) );
  AO221X1 U35032 ( .IN1(n31500), .IN2(n31499), .IN3(n31500), .IN4(n31498), 
        .IN5(\s6/msel/gnt_p1 [2]), .Q(n31501) );
  NAND3X0 U35033 ( .IN1(n31503), .IN2(n31502), .IN3(n31501), .QN(n17860) );
  NAND4X0 U35034 ( .IN1(n31507), .IN2(n34675), .IN3(n31505), .IN4(n31504), 
        .QN(n31517) );
  NAND2X0 U35035 ( .IN1(n31507), .IN2(n31506), .QN(n31518) );
  NAND3X0 U35036 ( .IN1(n31517), .IN2(n31518), .IN3(n31508), .QN(n31515) );
  NAND2X0 U35037 ( .IN1(n31509), .IN2(n31534), .QN(n31514) );
  NAND2X0 U35038 ( .IN1(n31511), .IN2(n31510), .QN(n31521) );
  NAND4X0 U35039 ( .IN1(\s6/msel/gnt_p0 [1]), .IN2(n31512), .IN3(n31530), 
        .IN4(n31521), .QN(n31513) );
  NAND3X0 U35040 ( .IN1(n31515), .IN2(n31514), .IN3(n31513), .QN(n31526) );
  NOR2X0 U35041 ( .IN1(n31530), .IN2(n31516), .QN(n31524) );
  OA221X1 U35042 ( .IN1(n31520), .IN2(n31519), .IN3(n31520), .IN4(n31518), 
        .IN5(n31517), .Q(n31522) );
  NAND2X0 U35043 ( .IN1(n31522), .IN2(n31521), .QN(n31523) );
  NOR2X0 U35044 ( .IN1(n31524), .IN2(n31523), .QN(n31525) );
  MUX21X1 U35045 ( .IN1(n31526), .IN2(n31525), .S(\s6/msel/gnt_p0 [2]), .Q(
        n31540) );
  AO21X1 U35046 ( .IN1(n31528), .IN2(n31540), .IN3(n31527), .Q(n31539) );
  NOR2X0 U35047 ( .IN1(\s6/msel/gnt_p0 [0]), .IN2(n31529), .QN(n31532) );
  NAND2X0 U35048 ( .IN1(n31540), .IN2(n31530), .QN(n31531) );
  NOR2X0 U35049 ( .IN1(n31532), .IN2(n31531), .QN(n31533) );
  NOR2X0 U35050 ( .IN1(n31533), .IN2(n34402), .QN(n31537) );
  NAND2X0 U35051 ( .IN1(n31535), .IN2(n31534), .QN(n31536) );
  NAND2X0 U35052 ( .IN1(n31537), .IN2(n31536), .QN(n31538) );
  AO22X1 U35053 ( .IN1(\s6/msel/gnt_p0 [1]), .IN2(n31540), .IN3(n31539), .IN4(
        n31538), .Q(n17858) );
  NAND3X0 U35054 ( .IN1(n13629), .IN2(m5s6_cyc), .IN3(n34531), .QN(n31588) );
  NAND2X0 U35055 ( .IN1(n34254), .IN2(n31588), .QN(n31620) );
  AND3X1 U35056 ( .IN1(n13577), .IN2(m6s6_cyc), .IN3(n34599), .Q(n31583) );
  NAND3X0 U35057 ( .IN1(n13525), .IN2(m7s6_cyc), .IN3(n34565), .QN(n31577) );
  INVX0 U35058 ( .INP(n31577), .ZN(n31603) );
  NOR2X0 U35059 ( .IN1(n31583), .IN2(n31603), .QN(n31548) );
  INVX0 U35060 ( .INP(n31548), .ZN(n31562) );
  NAND2X0 U35061 ( .IN1(\s6/msel/gnt_p2 [1]), .IN2(n31577), .QN(n31621) );
  OA21X1 U35062 ( .IN1(n31620), .IN2(n31562), .IN3(n31621), .Q(n31547) );
  NAND3X0 U35063 ( .IN1(n13785), .IN2(m2s6_cyc), .IN3(n34552), .QN(n31602) );
  NAND3X0 U35064 ( .IN1(n13733), .IN2(m3s6_cyc), .IN3(n34532), .QN(n31578) );
  NAND2X0 U35065 ( .IN1(n31602), .IN2(n31578), .QN(n31549) );
  INVX0 U35066 ( .INP(n31549), .ZN(n34117) );
  NAND3X0 U35067 ( .IN1(n13892), .IN2(m0s6_cyc), .IN3(n34579), .QN(n31579) );
  NAND3X0 U35068 ( .IN1(n13837), .IN2(m1s6_cyc), .IN3(n34368), .QN(n31582) );
  NAND2X0 U35069 ( .IN1(n31579), .IN2(n31582), .QN(n31561) );
  INVX0 U35070 ( .INP(n31561), .ZN(n34118) );
  NAND3X0 U35071 ( .IN1(n13681), .IN2(m4s6_cyc), .IN3(n34566), .QN(n31593) );
  INVX0 U35072 ( .INP(n31593), .ZN(n31581) );
  MUX21X1 U35073 ( .IN1(n31581), .IN2(n31583), .S(\s6/msel/gnt_p2 [1]), .Q(
        n31623) );
  AO22X1 U35074 ( .IN1(n34117), .IN2(n34118), .IN3(n34224), .IN4(n31623), .Q(
        n31546) );
  INVX0 U35075 ( .INP(n31582), .ZN(n31541) );
  NAND2X0 U35076 ( .IN1(n31541), .IN2(\s6/msel/gnt_p2 [0]), .QN(n31614) );
  OA21X1 U35077 ( .IN1(\s6/msel/gnt_p2 [0]), .IN2(n31579), .IN3(n31614), .Q(
        n31572) );
  NOR2X0 U35078 ( .IN1(\s6/msel/gnt_p2 [1]), .IN2(n31572), .QN(n31544) );
  NAND2X0 U35079 ( .IN1(n31593), .IN2(n31588), .QN(n31550) );
  NOR2X0 U35080 ( .IN1(n31550), .IN2(n31562), .QN(n34116) );
  INVX0 U35081 ( .INP(n31578), .ZN(n31552) );
  OR2X1 U35082 ( .IN1(\s6/msel/gnt_p2 [1]), .IN2(n31541), .Q(n31556) );
  OA22X1 U35083 ( .IN1(n31552), .IN2(n34254), .IN3(n31556), .IN4(n31549), .Q(
        n31543) );
  NAND2X0 U35084 ( .IN1(\s6/msel/gnt_p2 [1]), .IN2(n34224), .QN(n31553) );
  INVX0 U35085 ( .INP(n31553), .ZN(n31566) );
  INVX0 U35086 ( .INP(n31602), .ZN(n31615) );
  NAND2X0 U35087 ( .IN1(n31566), .IN2(n31615), .QN(n31542) );
  NOR2X0 U35088 ( .IN1(n34254), .IN2(n34224), .QN(n31558) );
  NAND2X0 U35089 ( .IN1(n31552), .IN2(n31558), .QN(n31618) );
  NAND3X0 U35090 ( .IN1(n31542), .IN2(n31618), .IN3(n34461), .QN(n31573) );
  NOR4X0 U35091 ( .IN1(n31544), .IN2(n34116), .IN3(n31543), .IN4(n31573), .QN(
        n31545) );
  AO221X1 U35092 ( .IN1(\s6/msel/gnt_p2 [2]), .IN2(n31547), .IN3(
        \s6/msel/gnt_p2 [2]), .IN4(n31546), .IN5(n31545), .Q(n17856) );
  NOR2X0 U35093 ( .IN1(n31548), .IN2(n31550), .QN(n31551) );
  NOR2X0 U35094 ( .IN1(n31551), .IN2(n31549), .QN(n31555) );
  NOR2X0 U35095 ( .IN1(n31550), .IN2(n31561), .QN(n31563) );
  NOR3X0 U35096 ( .IN1(n31552), .IN2(n31563), .IN3(n31551), .QN(n31554) );
  OA22X1 U35097 ( .IN1(n31556), .IN2(n31555), .IN3(n31554), .IN4(n31553), .Q(
        n31560) );
  OR2X1 U35098 ( .IN1(n31562), .IN2(n34118), .Q(n31557) );
  NAND4X0 U35099 ( .IN1(n31558), .IN2(n31593), .IN3(n31588), .IN4(n31557), 
        .QN(n31559) );
  NAND2X0 U35100 ( .IN1(n31560), .IN2(n31559), .QN(n31571) );
  NOR2X0 U35101 ( .IN1(n34117), .IN2(n31561), .QN(n31565) );
  OA22X1 U35102 ( .IN1(n31563), .IN2(n31621), .IN3(n31562), .IN4(
        \s6/msel/gnt_p2 [1]), .Q(n31564) );
  NOR2X0 U35103 ( .IN1(\s6/msel/gnt_p2 [1]), .IN2(\s6/msel/gnt_p2 [0]), .QN(
        n31589) );
  INVX0 U35104 ( .INP(n31589), .ZN(n31605) );
  OA22X1 U35105 ( .IN1(n31565), .IN2(n31564), .IN3(n31588), .IN4(n31605), .Q(
        n31567) );
  MUX21X1 U35106 ( .IN1(n31571), .IN2(n31567), .S(\s6/msel/gnt_p2 [2]), .Q(
        n31576) );
  AND3X1 U35107 ( .IN1(\s6/msel/gnt_p2 [0]), .IN2(\s6/msel/gnt_p2 [2]), .IN3(
        n31588), .Q(n31575) );
  NAND2X0 U35108 ( .IN1(n31566), .IN2(n31583), .QN(n31569) );
  NAND3X0 U35109 ( .IN1(n31567), .IN2(n34224), .IN3(n31593), .QN(n31568) );
  NAND3X0 U35110 ( .IN1(n31569), .IN2(n31568), .IN3(\s6/msel/gnt_p2 [2]), .QN(
        n31570) );
  OA221X1 U35111 ( .IN1(n31573), .IN2(n31572), .IN3(n31573), .IN4(n31571), 
        .IN5(n31570), .Q(n31574) );
  AO221X1 U35112 ( .IN1(n31576), .IN2(\s6/msel/gnt_p2 [1]), .IN3(n31576), 
        .IN4(n31575), .IN5(n31574), .Q(n17855) );
  INVX0 U35113 ( .INP(n31579), .ZN(n31613) );
  OA21X1 U35114 ( .IN1(n31613), .IN2(n31582), .IN3(n31577), .Q(n31597) );
  OA21X1 U35115 ( .IN1(n31581), .IN2(n31588), .IN3(n31578), .Q(n31595) );
  OA21X1 U35116 ( .IN1(n31581), .IN2(n34224), .IN3(n31595), .Q(n31580) );
  NAND2X0 U35117 ( .IN1(n31602), .IN2(n31579), .QN(n31584) );
  AO221X1 U35118 ( .IN1(n31597), .IN2(n31580), .IN3(n31597), .IN4(n31584), 
        .IN5(n31583), .Q(n31592) );
  NOR2X0 U35119 ( .IN1(n31583), .IN2(n31581), .QN(n31604) );
  INVX0 U35120 ( .INP(n31604), .ZN(n31596) );
  OA21X1 U35121 ( .IN1(n34224), .IN2(n31596), .IN3(n31595), .Q(n31599) );
  OA21X1 U35122 ( .IN1(n31615), .IN2(n31599), .IN3(n31582), .Q(n31607) );
  OR3X1 U35123 ( .IN1(n34254), .IN2(n31613), .IN3(n31607), .Q(n31591) );
  NOR2X0 U35124 ( .IN1(n34224), .IN2(n31583), .QN(n31586) );
  NAND2X0 U35125 ( .IN1(n31597), .IN2(n31584), .QN(n31585) );
  NAND2X0 U35126 ( .IN1(n31586), .IN2(n31585), .QN(n31587) );
  NAND2X0 U35127 ( .IN1(n31588), .IN2(n31587), .QN(n31594) );
  NAND2X0 U35128 ( .IN1(n31589), .IN2(n31594), .QN(n31590) );
  NAND4X0 U35129 ( .IN1(\s6/msel/gnt_p2 [2]), .IN2(n31592), .IN3(n31591), 
        .IN4(n31590), .QN(n31612) );
  NAND3X0 U35130 ( .IN1(\s6/msel/gnt_p2 [1]), .IN2(n31594), .IN3(n31593), .QN(
        n31610) );
  NAND2X0 U35131 ( .IN1(n31602), .IN2(n34254), .QN(n31601) );
  AND2X1 U35132 ( .IN1(n31613), .IN2(n31595), .Q(n31598) );
  OA22X1 U35133 ( .IN1(n31599), .IN2(n31598), .IN3(n31597), .IN4(n31596), .Q(
        n31600) );
  AO221X1 U35134 ( .IN1(\s6/msel/gnt_p2 [0]), .IN2(n31601), .IN3(n34224), 
        .IN4(n34254), .IN5(n31600), .Q(n31609) );
  NAND3X0 U35135 ( .IN1(n31604), .IN2(n31603), .IN3(n31602), .QN(n31606) );
  AO21X1 U35136 ( .IN1(n31607), .IN2(n31606), .IN3(n31605), .Q(n31608) );
  NAND4X0 U35137 ( .IN1(n34461), .IN2(n31610), .IN3(n31609), .IN4(n31608), 
        .QN(n31611) );
  NAND2X0 U35138 ( .IN1(n31612), .IN2(n31611), .QN(n31622) );
  AO221X1 U35139 ( .IN1(n31614), .IN2(n31613), .IN3(n31614), .IN4(n31622), 
        .IN5(\s6/msel/gnt_p2 [1]), .Q(n31617) );
  OR3X1 U35140 ( .IN1(n34254), .IN2(n31622), .IN3(n31615), .Q(n31616) );
  NAND3X0 U35141 ( .IN1(n31618), .IN2(n31617), .IN3(n31616), .QN(n31619) );
  NAND2X0 U35142 ( .IN1(n31619), .IN2(n34461), .QN(n31626) );
  NAND4X0 U35143 ( .IN1(\s6/msel/gnt_p2 [0]), .IN2(\s6/msel/gnt_p2 [2]), .IN3(
        n31621), .IN4(n31620), .QN(n31625) );
  AO221X1 U35144 ( .IN1(n34224), .IN2(n34461), .IN3(n34224), .IN4(n31623), 
        .IN5(n31622), .Q(n31624) );
  NAND3X0 U35145 ( .IN1(n31626), .IN2(n31625), .IN3(n31624), .QN(n17854) );
  NOR2X0 U35146 ( .IN1(n31627), .IN2(n34379), .QN(n31628) );
  MUX21X1 U35147 ( .IN1(n34349), .IN2(s15_data_o[0]), .S(n31628), .Q(n17853)
         );
  MUX21X1 U35148 ( .IN1(n34497), .IN2(s15_data_o[1]), .S(n31628), .Q(n17852)
         );
  MUX21X1 U35149 ( .IN1(n34348), .IN2(s15_data_o[2]), .S(n31628), .Q(n17851)
         );
  MUX21X1 U35150 ( .IN1(n34533), .IN2(s15_data_o[3]), .S(n31628), .Q(n17850)
         );
  MUX21X1 U35151 ( .IN1(n34363), .IN2(s15_data_o[4]), .S(n31628), .Q(n17849)
         );
  MUX21X1 U35152 ( .IN1(n34600), .IN2(s15_data_o[5]), .S(n31628), .Q(n17848)
         );
  MUX21X1 U35153 ( .IN1(n34318), .IN2(s15_data_o[6]), .S(n31628), .Q(n17847)
         );
  MUX21X1 U35154 ( .IN1(n34498), .IN2(s15_data_o[7]), .S(n31628), .Q(n17846)
         );
  MUX21X1 U35155 ( .IN1(n34649), .IN2(s15_data_o[8]), .S(n31628), .Q(n17845)
         );
  MUX21X1 U35156 ( .IN1(n34594), .IN2(s15_data_o[9]), .S(n31628), .Q(n17844)
         );
  MUX21X1 U35157 ( .IN1(n34350), .IN2(s15_data_o[10]), .S(n31628), .Q(n17843)
         );
  MUX21X1 U35158 ( .IN1(n34534), .IN2(s15_data_o[11]), .S(n31628), .Q(n17842)
         );
  MUX21X1 U35159 ( .IN1(n34374), .IN2(s15_data_o[12]), .S(n31628), .Q(n17841)
         );
  MUX21X1 U35160 ( .IN1(n34567), .IN2(s15_data_o[13]), .S(n31628), .Q(n17840)
         );
  MUX21X1 U35161 ( .IN1(n34347), .IN2(s15_data_o[14]), .S(n31628), .Q(n17839)
         );
  MUX21X1 U35162 ( .IN1(n34499), .IN2(s15_data_o[15]), .S(n31628), .Q(n17838)
         );
  NOR2X0 U35163 ( .IN1(n31683), .IN2(n31629), .QN(n31632) );
  AND2X1 U35164 ( .IN1(n31644), .IN2(\s7/msel/gnt_p3 [1]), .Q(n31631) );
  OA22X1 U35165 ( .IN1(n31632), .IN2(n31631), .IN3(n31630), .IN4(n31635), .Q(
        n31641) );
  INVX0 U35166 ( .INP(n31680), .ZN(n31660) );
  OAI221X1 U35167 ( .IN1(n31660), .IN2(n31652), .IN3(\s7/msel/gnt_p3 [1]), 
        .IN4(n31633), .IN5(n31671), .QN(n31640) );
  OA21X1 U35168 ( .IN1(\s7/msel/gnt_p3 [1]), .IN2(n31642), .IN3(n31634), .Q(
        n31685) );
  MUX21X1 U35169 ( .IN1(n31645), .IN2(n31643), .S(\s7/msel/gnt_p3 [1]), .Q(
        n31684) );
  NAND2X0 U35170 ( .IN1(n34410), .IN2(n31684), .QN(n31638) );
  NAND2X0 U35171 ( .IN1(n34262), .IN2(n31635), .QN(n31636) );
  NAND4X0 U35172 ( .IN1(n31685), .IN2(n31638), .IN3(n31637), .IN4(n31636), 
        .QN(n31639) );
  OA222X1 U35173 ( .IN1(\s7/msel/gnt_p3 [2]), .IN2(n31641), .IN3(
        \s7/msel/gnt_p3 [2]), .IN4(n31640), .IN5(n34380), .IN6(n31639), .Q(
        n17837) );
  INVX0 U35174 ( .INP(n31644), .ZN(n31682) );
  NOR3X0 U35175 ( .IN1(n31661), .IN2(n31681), .IN3(n31682), .QN(n31646) );
  OA21X1 U35176 ( .IN1(n31643), .IN2(n34410), .IN3(n31642), .Q(n31659) );
  OA21X1 U35177 ( .IN1(n31645), .IN2(n31659), .IN3(n31644), .Q(n31653) );
  NOR2X0 U35178 ( .IN1(n31646), .IN2(n31653), .QN(n31650) );
  NAND2X0 U35179 ( .IN1(n31670), .IN2(n31676), .QN(n31647) );
  NOR2X0 U35180 ( .IN1(n31657), .IN2(n31647), .QN(n31654) );
  NOR2X0 U35181 ( .IN1(n31660), .IN2(n31648), .QN(n31649) );
  OA21X1 U35182 ( .IN1(n31650), .IN2(n31654), .IN3(n31649), .Q(n31679) );
  INVX0 U35183 ( .INP(n31650), .ZN(n31651) );
  OR2X1 U35184 ( .IN1(n31652), .IN2(n31651), .Q(n31667) );
  OA21X1 U35185 ( .IN1(n31660), .IN2(n31653), .IN3(n31658), .Q(n31672) );
  INVX0 U35186 ( .INP(n31654), .ZN(n31656) );
  AO221X1 U35187 ( .IN1(n31672), .IN2(n31660), .IN3(n31672), .IN4(n31656), 
        .IN5(n31655), .Q(n31666) );
  INVX0 U35188 ( .INP(n31659), .ZN(n31663) );
  NOR2X0 U35189 ( .IN1(n31660), .IN2(n31673), .QN(n31668) );
  OR2X1 U35190 ( .IN1(n31661), .IN2(n31668), .Q(n31662) );
  AO22X1 U35191 ( .IN1(n31676), .IN2(n18195), .IN3(n31663), .IN4(n31662), .Q(
        n31664) );
  NAND3X0 U35192 ( .IN1(\s7/msel/gnt_p3 [1]), .IN2(n31664), .IN3(n31670), .QN(
        n31665) );
  NAND4X0 U35193 ( .IN1(n34380), .IN2(n31667), .IN3(n31666), .IN4(n31665), 
        .QN(n31678) );
  OA221X1 U35194 ( .IN1(n31682), .IN2(n31670), .IN3(n31682), .IN4(n31669), 
        .IN5(n31668), .Q(n31675) );
  NOR3X0 U35195 ( .IN1(n31673), .IN2(n31672), .IN3(n31671), .QN(n31674) );
  AO221X1 U35196 ( .IN1(n31676), .IN2(n18195), .IN3(n31676), .IN4(n31675), 
        .IN5(n31674), .Q(n31677) );
  OA22X1 U35197 ( .IN1(n31679), .IN2(n31678), .IN3(n34380), .IN4(n31677), .Q(
        n31687) );
  OA221X1 U35198 ( .IN1(\s7/msel/gnt_p3 [1]), .IN2(n31681), .IN3(n34262), 
        .IN4(n31680), .IN5(n31687), .Q(n31691) );
  OA221X1 U35199 ( .IN1(\s7/msel/gnt_p3 [1]), .IN2(n31683), .IN3(n34262), 
        .IN4(n31682), .IN5(\s7/msel/gnt_p3 [0]), .Q(n31690) );
  NOR2X0 U35200 ( .IN1(n34380), .IN2(n31684), .QN(n31688) );
  NOR2X0 U35201 ( .IN1(n31685), .IN2(n34380), .QN(n31686) );
  OA22X1 U35202 ( .IN1(\s7/msel/gnt_p3 [0]), .IN2(n31688), .IN3(n31687), .IN4(
        n31686), .Q(n31689) );
  AO221X1 U35203 ( .IN1(n34380), .IN2(n31691), .IN3(n34380), .IN4(n31690), 
        .IN5(n31689), .Q(n17835) );
  NAND2X0 U35204 ( .IN1(n34129), .IN2(n31696), .QN(n31692) );
  AND3X1 U35205 ( .IN1(n34130), .IN2(\s7/msel/gnt_p1 [1]), .IN3(n31692), .Q(
        n31707) );
  INVX0 U35206 ( .INP(n31737), .ZN(n31695) );
  AO221X1 U35207 ( .IN1(n34130), .IN2(\s7/msel/gnt_p1 [1]), .IN3(n34130), 
        .IN4(n31701), .IN5(n31699), .Q(n31698) );
  AO22X1 U35208 ( .IN1(n31695), .IN2(n31694), .IN3(n31693), .IN4(n31698), .Q(
        n31706) );
  INVX0 U35209 ( .INP(n31696), .ZN(n31700) );
  AO22X1 U35210 ( .IN1(n31700), .IN2(n31698), .IN3(n34245), .IN4(n31697), .Q(
        n31703) );
  OA221X1 U35211 ( .IN1(n31701), .IN2(n31700), .IN3(n31701), .IN4(n31699), 
        .IN5(n31734), .Q(n31702) );
  NAND2X0 U35212 ( .IN1(n34245), .IN2(n34439), .QN(n31739) );
  OA22X1 U35213 ( .IN1(n31704), .IN2(n31703), .IN3(n31702), .IN4(n31739), .Q(
        n31705) );
  AO222X1 U35214 ( .IN1(n34424), .IN2(n31707), .IN3(n34424), .IN4(n31706), 
        .IN5(\s7/msel/gnt_p1 [2]), .IN6(n31705), .Q(n31719) );
  AO21X1 U35215 ( .IN1(n31719), .IN2(n31709), .IN3(n31708), .Q(n31718) );
  AO221X1 U35216 ( .IN1(\s7/msel/gnt_p1 [0]), .IN2(n31720), .IN3(n34245), 
        .IN4(n31710), .IN5(n34439), .Q(n31716) );
  INVX0 U35217 ( .INP(n31719), .ZN(n31711) );
  NOR2X0 U35218 ( .IN1(n31712), .IN2(n31711), .QN(n31714) );
  NAND2X0 U35219 ( .IN1(n34245), .IN2(n31733), .QN(n31713) );
  NAND2X0 U35220 ( .IN1(n31714), .IN2(n31713), .QN(n31715) );
  NAND3X0 U35221 ( .IN1(\s7/msel/gnt_p1 [2]), .IN2(n31716), .IN3(n31715), .QN(
        n31717) );
  AO22X1 U35222 ( .IN1(\s7/msel/gnt_p1 [1]), .IN2(n31719), .IN3(n31718), .IN4(
        n31717), .Q(n17833) );
  INVX0 U35223 ( .INP(n31750), .ZN(n31731) );
  OA21X1 U35224 ( .IN1(n31731), .IN2(n31748), .IN3(n31720), .Q(n31735) );
  OA21X1 U35225 ( .IN1(n31742), .IN2(n31735), .IN3(n31734), .Q(n31740) );
  NOR3X0 U35226 ( .IN1(n31733), .IN2(n31740), .IN3(n31729), .QN(n31747) );
  NOR2X0 U35227 ( .IN1(n31733), .IN2(n31742), .QN(n31721) );
  NAND3X0 U35228 ( .IN1(n31721), .IN2(\s7/msel/gnt_p1 [0]), .IN3(n31750), .QN(
        n31722) );
  OA21X1 U35229 ( .IN1(n31733), .IN2(n31734), .IN3(n31737), .Q(n31725) );
  NAND2X0 U35230 ( .IN1(n31722), .IN2(n31725), .QN(n31724) );
  NOR3X0 U35231 ( .IN1(n31742), .IN2(n31733), .IN3(n31735), .QN(n31723) );
  NOR2X0 U35232 ( .IN1(n31724), .IN2(n31723), .QN(n31726) );
  OA21X1 U35233 ( .IN1(n31727), .IN2(n31725), .IN3(n31748), .Q(n31730) );
  OA22X1 U35234 ( .IN1(n31727), .IN2(n31726), .IN3(n31730), .IN4(n31739), .Q(
        n31728) );
  NAND2X0 U35235 ( .IN1(n31728), .IN2(n34424), .QN(n31746) );
  NOR3X0 U35236 ( .IN1(n31731), .IN2(n31730), .IN3(n31729), .QN(n31745) );
  NAND2X0 U35237 ( .IN1(n31750), .IN2(n31732), .QN(n31738) );
  AO21X1 U35238 ( .IN1(n34245), .IN2(n31734), .IN3(n31733), .Q(n31736) );
  OA221X1 U35239 ( .IN1(n31738), .IN2(n31737), .IN3(n31738), .IN4(n31736), 
        .IN5(n31735), .Q(n31741) );
  OA22X1 U35240 ( .IN1(n31742), .IN2(n31741), .IN3(n31740), .IN4(n31739), .Q(
        n31743) );
  NAND2X0 U35241 ( .IN1(\s7/msel/gnt_p1 [2]), .IN2(n31743), .QN(n31744) );
  OA22X1 U35242 ( .IN1(n31747), .IN2(n31746), .IN3(n31745), .IN4(n31744), .Q(
        n31753) );
  NOR2X0 U35243 ( .IN1(n34245), .IN2(n31748), .QN(n31749) );
  AO222X1 U35244 ( .IN1(n31753), .IN2(\s7/msel/gnt_p1 [1]), .IN3(n31753), 
        .IN4(n31750), .IN5(n34439), .IN6(n31749), .Q(n31751) );
  OAI21X1 U35245 ( .IN1(n31752), .IN2(n31751), .IN3(n34424), .QN(n31758) );
  INVX0 U35246 ( .INP(n31753), .ZN(n31754) );
  AO221X1 U35247 ( .IN1(n34245), .IN2(n31755), .IN3(n34245), .IN4(n34424), 
        .IN5(n31754), .Q(n31756) );
  NAND3X0 U35248 ( .IN1(n31758), .IN2(n31757), .IN3(n31756), .QN(n17832) );
  NAND3X0 U35249 ( .IN1(n13630), .IN2(n13604), .IN3(m5s7_cyc), .QN(n31806) );
  NAND2X0 U35250 ( .IN1(n34414), .IN2(n31806), .QN(n31761) );
  NAND3X0 U35251 ( .IN1(n13526), .IN2(n13470), .IN3(m7s7_cyc), .QN(n31759) );
  NAND2X0 U35252 ( .IN1(\s7/msel/gnt_p0 [1]), .IN2(n31759), .QN(n31760) );
  NAND4X0 U35253 ( .IN1(\s7/msel/gnt_p0 [2]), .IN2(\s7/msel/gnt_p0 [0]), .IN3(
        n31761), .IN4(n31760), .QN(n31853) );
  NAND3X0 U35254 ( .IN1(n13894), .IN2(n13864), .IN3(m0s7_cyc), .QN(n31844) );
  INVX0 U35255 ( .INP(n31844), .ZN(n31835) );
  NAND3X0 U35256 ( .IN1(n13838), .IN2(n13812), .IN3(m1s7_cyc), .QN(n31807) );
  INVX0 U35257 ( .INP(n31807), .ZN(n31814) );
  NOR2X0 U35258 ( .IN1(n31835), .IN2(n31814), .QN(n31789) );
  NAND3X0 U35259 ( .IN1(n13786), .IN2(n13760), .IN3(m2s7_cyc), .QN(n31843) );
  NAND3X0 U35260 ( .IN1(n13734), .IN2(n13708), .IN3(m3s7_cyc), .QN(n31831) );
  NAND2X0 U35261 ( .IN1(n31843), .IN2(n31831), .QN(n31788) );
  INVX0 U35262 ( .INP(n31788), .ZN(n31776) );
  NAND2X0 U35263 ( .IN1(n31789), .IN2(n31776), .QN(n31763) );
  NAND3X0 U35264 ( .IN1(n13578), .IN2(n13552), .IN3(m6s7_cyc), .QN(n31818) );
  NAND3X0 U35265 ( .IN1(n13682), .IN2(n13656), .IN3(m4s7_cyc), .QN(n31821) );
  AO221X1 U35266 ( .IN1(\s7/msel/gnt_p0 [1]), .IN2(n31818), .IN3(n34414), 
        .IN4(n31821), .IN5(\s7/msel/gnt_p0 [0]), .Q(n31850) );
  NAND2X0 U35267 ( .IN1(n31818), .IN2(n31759), .QN(n31787) );
  INVX0 U35268 ( .INP(n31759), .ZN(n31812) );
  NOR2X0 U35269 ( .IN1(\s7/msel/gnt_p0 [1]), .IN2(n34289), .QN(n31775) );
  NAND2X0 U35270 ( .IN1(n31775), .IN2(n31818), .QN(n31825) );
  OA21X1 U35271 ( .IN1(n31812), .IN2(n31825), .IN3(n31760), .Q(n31785) );
  OAI21X1 U35272 ( .IN1(n31761), .IN2(n31787), .IN3(n31785), .QN(n31762) );
  NAND3X0 U35273 ( .IN1(n31763), .IN2(n31850), .IN3(n31762), .QN(n31764) );
  NAND2X0 U35274 ( .IN1(n31764), .IN2(\s7/msel/gnt_p0 [2]), .QN(n31773) );
  NAND2X0 U35275 ( .IN1(\s7/msel/gnt_p0 [0]), .IN2(\s7/msel/gnt_p0 [1]), .QN(
        n31768) );
  NOR2X0 U35276 ( .IN1(n31831), .IN2(n31768), .QN(n31845) );
  NOR2X0 U35277 ( .IN1(\s7/msel/gnt_p0 [2]), .IN2(n31845), .QN(n31766) );
  INVX0 U35278 ( .INP(n31843), .ZN(n31813) );
  NOR2X0 U35279 ( .IN1(\s7/msel/gnt_p0 [0]), .IN2(n34414), .QN(n31797) );
  NAND2X0 U35280 ( .IN1(n31813), .IN2(n31797), .QN(n31765) );
  NAND2X0 U35281 ( .IN1(n31766), .IN2(n31765), .QN(n31795) );
  NAND2X0 U35282 ( .IN1(\s7/msel/gnt_p0 [0]), .IN2(n31814), .QN(n31847) );
  OA21X1 U35283 ( .IN1(\s7/msel/gnt_p0 [0]), .IN2(n31844), .IN3(n31847), .Q(
        n31796) );
  NAND2X0 U35284 ( .IN1(n31806), .IN2(n31821), .QN(n31783) );
  OAI22X1 U35285 ( .IN1(\s7/msel/gnt_p0 [1]), .IN2(n31796), .IN3(n31783), 
        .IN4(n31787), .QN(n31767) );
  NOR2X0 U35286 ( .IN1(n31795), .IN2(n31767), .QN(n31771) );
  NAND2X0 U35287 ( .IN1(n34289), .IN2(n34414), .QN(n31830) );
  NOR2X0 U35288 ( .IN1(n31814), .IN2(n31830), .QN(n31774) );
  AO21X1 U35289 ( .IN1(n31775), .IN2(n31843), .IN3(n31797), .Q(n31841) );
  AOI22X1 U35290 ( .IN1(n31774), .IN2(n31776), .IN3(n31831), .IN4(n31841), 
        .QN(n31769) );
  NAND2X0 U35291 ( .IN1(n31769), .IN2(n31768), .QN(n31770) );
  NAND2X0 U35292 ( .IN1(n31771), .IN2(n31770), .QN(n31772) );
  NAND3X0 U35293 ( .IN1(n31853), .IN2(n31773), .IN3(n31772), .QN(n17831) );
  NOR2X0 U35294 ( .IN1(n31775), .IN2(n31774), .QN(n31779) );
  INVX0 U35295 ( .INP(n31787), .ZN(n31777) );
  OA21X1 U35296 ( .IN1(n31777), .IN2(n31783), .IN3(n31776), .Q(n31778) );
  INVX0 U35297 ( .INP(n31797), .ZN(n31826) );
  OA22X1 U35298 ( .IN1(n31779), .IN2(n31778), .IN3(n31831), .IN4(n31826), .Q(
        n31782) );
  OR2X1 U35299 ( .IN1(n31787), .IN2(n31789), .Q(n31780) );
  NAND4X0 U35300 ( .IN1(\s7/msel/gnt_p0 [1]), .IN2(n31821), .IN3(n31806), 
        .IN4(n31780), .QN(n31781) );
  NAND2X0 U35301 ( .IN1(n31782), .IN2(n31781), .QN(n31794) );
  INVX0 U35302 ( .INP(n31825), .ZN(n31784) );
  NOR2X0 U35303 ( .IN1(n31784), .IN2(n31783), .QN(n31786) );
  AO221X1 U35304 ( .IN1(n31789), .IN2(n31786), .IN3(n31789), .IN4(n31788), 
        .IN5(n31785), .Q(n31793) );
  NOR2X0 U35305 ( .IN1(n31787), .IN2(n31830), .QN(n31791) );
  NAND2X0 U35306 ( .IN1(n31789), .IN2(n31788), .QN(n31790) );
  NAND2X0 U35307 ( .IN1(n31791), .IN2(n31790), .QN(n31792) );
  OA221X1 U35308 ( .IN1(\s7/msel/gnt_p0 [2]), .IN2(n31794), .IN3(n34550), 
        .IN4(n31793), .IN5(n31792), .Q(n31803) );
  AO21X1 U35309 ( .IN1(n31796), .IN2(n31803), .IN3(n31795), .Q(n31802) );
  INVX0 U35310 ( .INP(n31818), .ZN(n31810) );
  NAND2X0 U35311 ( .IN1(n31810), .IN2(n31797), .QN(n31800) );
  INVX0 U35312 ( .INP(n31821), .ZN(n31809) );
  NAND2X0 U35313 ( .IN1(n31809), .IN2(n34289), .QN(n31798) );
  NAND3X0 U35314 ( .IN1(n31806), .IN2(n31803), .IN3(n31798), .QN(n31799) );
  NAND3X0 U35315 ( .IN1(\s7/msel/gnt_p0 [2]), .IN2(n31800), .IN3(n31799), .QN(
        n31801) );
  AO22X1 U35316 ( .IN1(\s7/msel/gnt_p0 [1]), .IN2(n31803), .IN3(n31802), .IN4(
        n31801), .Q(n17830) );
  NOR2X0 U35317 ( .IN1(n31835), .IN2(n31807), .QN(n31804) );
  NOR2X0 U35318 ( .IN1(n31812), .IN2(n31804), .QN(n31828) );
  NAND2X0 U35319 ( .IN1(n31843), .IN2(n31844), .QN(n31822) );
  OR2X1 U35320 ( .IN1(n31822), .IN2(n31810), .Q(n31832) );
  OA22X1 U35321 ( .IN1(n31810), .IN2(n31828), .IN3(n34289), .IN4(n31832), .Q(
        n31805) );
  NAND2X0 U35322 ( .IN1(n31805), .IN2(n31806), .QN(n31829) );
  NAND3X0 U35323 ( .IN1(\s7/msel/gnt_p0 [1]), .IN2(n31821), .IN3(n31829), .QN(
        n31817) );
  OA21X1 U35324 ( .IN1(n31809), .IN2(n31806), .IN3(n31831), .Q(n31824) );
  NAND3X0 U35325 ( .IN1(\s7/msel/gnt_p0 [0]), .IN2(n31818), .IN3(n31821), .QN(
        n31808) );
  OA221X1 U35326 ( .IN1(n31813), .IN2(n31824), .IN3(n31813), .IN4(n31808), 
        .IN5(n31807), .Q(n31834) );
  NOR2X0 U35327 ( .IN1(n31810), .IN2(n31809), .QN(n31811) );
  NAND2X0 U35328 ( .IN1(n31812), .IN2(n31811), .QN(n31819) );
  AO221X1 U35329 ( .IN1(n31834), .IN2(n31813), .IN3(n31834), .IN4(n31819), 
        .IN5(n31830), .Q(n31816) );
  NAND4X0 U35330 ( .IN1(n31814), .IN2(n31844), .IN3(n31818), .IN4(n31821), 
        .QN(n31815) );
  NAND4X0 U35331 ( .IN1(n34550), .IN2(n31817), .IN3(n31816), .IN4(n31815), 
        .QN(n31842) );
  NAND4X0 U35332 ( .IN1(\s7/msel/gnt_p0 [0]), .IN2(n31818), .IN3(n31844), 
        .IN4(n31821), .QN(n31820) );
  NAND3X0 U35333 ( .IN1(n31824), .IN2(n31820), .IN3(n31819), .QN(n31840) );
  NAND2X0 U35334 ( .IN1(\s7/msel/gnt_p0 [0]), .IN2(n31821), .QN(n31823) );
  AO21X1 U35335 ( .IN1(n31824), .IN2(n31823), .IN3(n31822), .Q(n31827) );
  AO22X1 U35336 ( .IN1(n31828), .IN2(n31827), .IN3(n31826), .IN4(n31825), .Q(
        n31838) );
  INVX0 U35337 ( .INP(n31829), .ZN(n31833) );
  AO221X1 U35338 ( .IN1(n31833), .IN2(n31832), .IN3(n31833), .IN4(n31831), 
        .IN5(n31830), .Q(n31837) );
  OR3X1 U35339 ( .IN1(n34414), .IN2(n31835), .IN3(n31834), .Q(n31836) );
  NAND4X0 U35340 ( .IN1(\s7/msel/gnt_p0 [2]), .IN2(n31838), .IN3(n31837), 
        .IN4(n31836), .QN(n31839) );
  OA221X1 U35341 ( .IN1(n31842), .IN2(n31841), .IN3(n31842), .IN4(n31840), 
        .IN5(n31839), .Q(n31849) );
  OA221X1 U35342 ( .IN1(\s7/msel/gnt_p0 [1]), .IN2(n31844), .IN3(n34414), 
        .IN4(n31843), .IN5(n31849), .Q(n31846) );
  NOR2X0 U35343 ( .IN1(n31846), .IN2(n31845), .QN(n31848) );
  AO221X1 U35344 ( .IN1(n31848), .IN2(\s7/msel/gnt_p0 [1]), .IN3(n31848), 
        .IN4(n31847), .IN5(\s7/msel/gnt_p0 [2]), .Q(n31854) );
  NAND2X0 U35345 ( .IN1(n34550), .IN2(n34289), .QN(n31851) );
  NAND3X0 U35346 ( .IN1(n31851), .IN2(n31850), .IN3(n31849), .QN(n31852) );
  NAND3X0 U35347 ( .IN1(n31854), .IN2(n31853), .IN3(n31852), .QN(n17829) );
  NAND2X0 U35348 ( .IN1(\s7/msel/gnt_p2 [1]), .IN2(n31892), .QN(n31874) );
  OA21X1 U35349 ( .IN1(\s7/msel/gnt_p2 [1]), .IN2(n31902), .IN3(n31874), .Q(
        n31855) );
  NAND3X0 U35350 ( .IN1(\s7/msel/gnt_p2 [0]), .IN2(\s7/msel/gnt_p2 [2]), .IN3(
        n31855), .QN(n31936) );
  NOR2X0 U35351 ( .IN1(\s7/msel/gnt_p2 [1]), .IN2(n31908), .QN(n31934) );
  NOR2X0 U35352 ( .IN1(n31855), .IN2(n31934), .QN(n31857) );
  INVX0 U35353 ( .INP(n31916), .ZN(n31894) );
  NAND2X0 U35354 ( .IN1(\s7/msel/gnt_p2 [1]), .IN2(n31894), .QN(n31882) );
  NAND2X0 U35355 ( .IN1(n34133), .IN2(n34134), .QN(n31856) );
  OA221X1 U35356 ( .IN1(\s7/msel/gnt_p2 [0]), .IN2(n31857), .IN3(
        \s7/msel/gnt_p2 [0]), .IN4(n31882), .IN5(n31856), .Q(n31859) );
  AO221X1 U35357 ( .IN1(n31859), .IN2(\s7/msel/gnt_p2 [1]), .IN3(n31859), 
        .IN4(n31858), .IN5(n34435), .Q(n31864) );
  OR2X1 U35358 ( .IN1(n34429), .IN2(n31898), .Q(n31928) );
  OA21X1 U35359 ( .IN1(\s7/msel/gnt_p2 [0]), .IN2(n31895), .IN3(n31928), .Q(
        n31885) );
  NOR2X0 U35360 ( .IN1(\s7/msel/gnt_p2 [1]), .IN2(n31885), .QN(n31862) );
  AND2X1 U35361 ( .IN1(n34274), .IN2(n31898), .Q(n31871) );
  AOI22X1 U35362 ( .IN1(\s7/msel/gnt_p2 [1]), .IN2(n31890), .IN3(n34134), 
        .IN4(n31871), .QN(n31861) );
  NOR2X0 U35363 ( .IN1(\s7/msel/gnt_p2 [0]), .IN2(n34274), .QN(n31914) );
  NAND2X0 U35364 ( .IN1(n31914), .IN2(n31906), .QN(n31860) );
  NOR2X0 U35365 ( .IN1(n34429), .IN2(n34274), .QN(n31866) );
  NAND2X0 U35366 ( .IN1(n31917), .IN2(n31866), .QN(n31930) );
  NAND3X0 U35367 ( .IN1(n31860), .IN2(n31930), .IN3(n34435), .QN(n31886) );
  OR4X1 U35368 ( .IN1(n31862), .IN2(n34132), .IN3(n31861), .IN4(n31886), .Q(
        n31863) );
  NAND3X0 U35369 ( .IN1(n31936), .IN2(n31864), .IN3(n31863), .QN(n17828) );
  AO21X1 U35370 ( .IN1(\s7/msel/gnt_p2 [1]), .IN2(n34133), .IN3(n31867), .Q(
        n31865) );
  AND3X1 U35371 ( .IN1(n31866), .IN2(n31868), .IN3(n31865), .Q(n31881) );
  NAND2X0 U35372 ( .IN1(n34133), .IN2(n31868), .QN(n31876) );
  NAND2X0 U35373 ( .IN1(n31868), .IN2(n31867), .QN(n31869) );
  NAND3X0 U35374 ( .IN1(n31890), .IN2(n31876), .IN3(n31869), .QN(n31872) );
  NAND2X0 U35375 ( .IN1(n34134), .IN2(n31869), .QN(n31870) );
  AO22X1 U35376 ( .IN1(n31914), .IN2(n31872), .IN3(n31871), .IN4(n31870), .Q(
        n31880) );
  NOR2X0 U35377 ( .IN1(n34134), .IN2(n31873), .QN(n31878) );
  NOR2X0 U35378 ( .IN1(n31894), .IN2(\s7/msel/gnt_p2 [1]), .QN(n31913) );
  INVX0 U35379 ( .INP(n31874), .ZN(n31875) );
  AOI22X1 U35380 ( .IN1(n31892), .IN2(n31913), .IN3(n31876), .IN4(n31875), 
        .QN(n31877) );
  NAND2X0 U35381 ( .IN1(n34429), .IN2(n34274), .QN(n31919) );
  OA22X1 U35382 ( .IN1(n31878), .IN2(n31877), .IN3(n31891), .IN4(n31919), .Q(
        n31879) );
  AO222X1 U35383 ( .IN1(n34435), .IN2(n31881), .IN3(n34435), .IN4(n31880), 
        .IN5(n31879), .IN6(\s7/msel/gnt_p2 [2]), .Q(n31889) );
  NAND2X0 U35384 ( .IN1(\s7/msel/gnt_p2 [0]), .IN2(\s7/msel/gnt_p2 [2]), .QN(
        n31883) );
  NOR2X0 U35385 ( .IN1(n31902), .IN2(n31883), .QN(n31888) );
  NAND2X0 U35386 ( .IN1(\s7/msel/gnt_p2 [2]), .IN2(n31882), .QN(n31933) );
  OA221X1 U35387 ( .IN1(n31933), .IN2(n31908), .IN3(n31933), .IN4(n31889), 
        .IN5(n31883), .Q(n31884) );
  OA221X1 U35388 ( .IN1(n31886), .IN2(n31885), .IN3(n31886), .IN4(n31889), 
        .IN5(n31884), .Q(n31887) );
  AO221X1 U35389 ( .IN1(n31889), .IN2(\s7/msel/gnt_p2 [1]), .IN3(n31889), 
        .IN4(n31888), .IN5(n31887), .Q(n17827) );
  OA21X1 U35390 ( .IN1(n31891), .IN2(n31893), .IN3(n31890), .Q(n31900) );
  INVX0 U35391 ( .INP(n31900), .ZN(n31907) );
  INVX0 U35392 ( .INP(n31895), .ZN(n31929) );
  OA21X1 U35393 ( .IN1(n31898), .IN2(n31929), .IN3(n31892), .Q(n31909) );
  INVX0 U35394 ( .INP(n31909), .ZN(n31903) );
  NOR2X0 U35395 ( .IN1(n31894), .IN2(n31893), .QN(n31897) );
  OA221X1 U35396 ( .IN1(n31903), .IN2(\s7/msel/gnt_p2 [0]), .IN3(n31903), 
        .IN4(n31895), .IN5(n31897), .Q(n31896) );
  NOR2X0 U35397 ( .IN1(n31907), .IN2(n31896), .QN(n31901) );
  NAND2X0 U35398 ( .IN1(\s7/msel/gnt_p2 [0]), .IN2(n31897), .QN(n31899) );
  OA221X1 U35399 ( .IN1(n31906), .IN2(n31900), .IN3(n31906), .IN4(n31899), 
        .IN5(n31898), .Q(n31922) );
  OA22X1 U35400 ( .IN1(n31906), .IN2(n31901), .IN3(n31922), .IN4(n31919), .Q(
        n31905) );
  AO21X1 U35401 ( .IN1(n31916), .IN2(n31903), .IN3(n31902), .Q(n31915) );
  NAND4X0 U35402 ( .IN1(\s7/msel/gnt_p2 [1]), .IN2(\s7/msel/gnt_p2 [0]), .IN3(
        n31915), .IN4(n31908), .QN(n31904) );
  NAND3X0 U35403 ( .IN1(n34435), .IN2(n31905), .IN3(n31904), .QN(n31927) );
  NOR2X0 U35404 ( .IN1(n31929), .IN2(n31906), .QN(n31918) );
  AND2X1 U35405 ( .IN1(n31907), .IN2(n31918), .Q(n31912) );
  NAND3X0 U35406 ( .IN1(\s7/msel/gnt_p2 [0]), .IN2(n31918), .IN3(n31908), .QN(
        n31910) );
  NAND2X0 U35407 ( .IN1(n31910), .IN2(n31909), .QN(n31911) );
  OAI22X1 U35408 ( .IN1(n31914), .IN2(n31913), .IN3(n31912), .IN4(n31911), 
        .QN(n31925) );
  INVX0 U35409 ( .INP(n31915), .ZN(n31921) );
  NAND3X0 U35410 ( .IN1(n31918), .IN2(n31917), .IN3(n31916), .QN(n31920) );
  AO21X1 U35411 ( .IN1(n31921), .IN2(n31920), .IN3(n31919), .Q(n31924) );
  OR3X1 U35412 ( .IN1(n34274), .IN2(n31929), .IN3(n31922), .Q(n31923) );
  NAND4X0 U35413 ( .IN1(\s7/msel/gnt_p2 [2]), .IN2(n31925), .IN3(n31924), 
        .IN4(n31923), .QN(n31926) );
  NAND2X0 U35414 ( .IN1(n31927), .IN2(n31926), .QN(n31932) );
  OA222X1 U35415 ( .IN1(n31932), .IN2(n31929), .IN3(n31932), .IN4(n34274), 
        .IN5(\s7/msel/gnt_p2 [1]), .IN6(n31928), .Q(n31931) );
  AO21X1 U35416 ( .IN1(n31931), .IN2(n31930), .IN3(\s7/msel/gnt_p2 [2]), .Q(
        n31937) );
  AO221X1 U35417 ( .IN1(n34429), .IN2(n31934), .IN3(n34429), .IN4(n31933), 
        .IN5(n31932), .Q(n31935) );
  NAND3X0 U35418 ( .IN1(n31937), .IN2(n31936), .IN3(n31935), .QN(n17826) );
  NOR2X0 U35419 ( .IN1(n31938), .IN2(n34379), .QN(n31939) );
  MUX21X1 U35420 ( .IN1(n34659), .IN2(s15_data_o[0]), .S(n31939), .Q(n17825)
         );
  MUX21X1 U35421 ( .IN1(n34589), .IN2(s15_data_o[1]), .S(n31939), .Q(n17824)
         );
  MUX21X1 U35422 ( .IN1(n34660), .IN2(s15_data_o[2]), .S(n31939), .Q(n17823)
         );
  MUX21X1 U35423 ( .IN1(n34593), .IN2(s15_data_o[3]), .S(n31939), .Q(n17822)
         );
  MUX21X1 U35424 ( .IN1(n34662), .IN2(s15_data_o[4]), .S(n31939), .Q(n17821)
         );
  MUX21X1 U35425 ( .IN1(n34591), .IN2(s15_data_o[5]), .S(n31939), .Q(n17820)
         );
  MUX21X1 U35426 ( .IN1(n34663), .IN2(s15_data_o[6]), .S(n31939), .Q(n17819)
         );
  MUX21X1 U35427 ( .IN1(n34590), .IN2(s15_data_o[7]), .S(n31939), .Q(n17818)
         );
  MUX21X1 U35428 ( .IN1(n34238), .IN2(s15_data_o[8]), .S(n31939), .Q(n17817)
         );
  MUX21X1 U35429 ( .IN1(n34369), .IN2(s15_data_o[9]), .S(n31939), .Q(n17816)
         );
  MUX21X1 U35430 ( .IN1(n34588), .IN2(s15_data_o[10]), .S(n31939), .Q(n17815)
         );
  MUX21X1 U35431 ( .IN1(n34239), .IN2(s15_data_o[11]), .S(n31939), .Q(n17814)
         );
  MUX21X1 U35432 ( .IN1(n34631), .IN2(s15_data_o[12]), .S(n31939), .Q(n17813)
         );
  MUX21X1 U35433 ( .IN1(n34580), .IN2(s15_data_o[13]), .S(n31939), .Q(n17812)
         );
  MUX21X1 U35434 ( .IN1(n34661), .IN2(s15_data_o[14]), .S(n31939), .Q(n17811)
         );
  MUX21X1 U35435 ( .IN1(n34592), .IN2(s15_data_o[15]), .S(n31939), .Q(n17810)
         );
  OR2X1 U35436 ( .IN1(n31973), .IN2(n31958), .Q(n31954) );
  NAND2X0 U35437 ( .IN1(n34223), .IN2(n31954), .QN(n31942) );
  NOR2X0 U35438 ( .IN1(n31945), .IN2(n31946), .QN(n31960) );
  NOR2X0 U35439 ( .IN1(n31962), .IN2(n31955), .QN(n31959) );
  NAND2X0 U35440 ( .IN1(n31960), .IN2(n31959), .QN(n34142) );
  NAND2X0 U35441 ( .IN1(n34228), .IN2(n31940), .QN(n31941) );
  NAND4X0 U35442 ( .IN1(n31943), .IN2(n31942), .IN3(n34142), .IN4(n31941), 
        .QN(n31953) );
  OA21X1 U35443 ( .IN1(n31944), .IN2(n31959), .IN3(n34456), .Q(n31970) );
  AO21X1 U35444 ( .IN1(n31946), .IN2(n34228), .IN3(n31945), .Q(n31972) );
  INVX0 U35445 ( .INP(n31972), .ZN(n31947) );
  NOR2X0 U35446 ( .IN1(n31947), .IN2(\s8/msel/gnt_p3 [1]), .QN(n31951) );
  NAND2X0 U35447 ( .IN1(n31948), .IN2(n31961), .QN(n31968) );
  OR2X1 U35448 ( .IN1(n31968), .IN2(n31954), .Q(n34143) );
  NAND2X0 U35449 ( .IN1(n34143), .IN2(n31949), .QN(n31950) );
  NOR2X0 U35450 ( .IN1(n31951), .IN2(n31950), .QN(n31952) );
  AO22X1 U35451 ( .IN1(\s8/msel/gnt_p3 [2]), .IN2(n31953), .IN3(n31970), .IN4(
        n31952), .Q(n17809) );
  AOI21X1 U35452 ( .IN1(\s8/msel/gnt_p3 [1]), .IN2(n31960), .IN3(n31954), .QN(
        n31969) );
  AO21X1 U35453 ( .IN1(n31960), .IN2(n31955), .IN3(n31954), .Q(n31956) );
  NAND2X0 U35454 ( .IN1(n34223), .IN2(n31956), .QN(n31957) );
  NOR2X0 U35455 ( .IN1(n31977), .IN2(n31957), .QN(n31966) );
  AND2X1 U35456 ( .IN1(n31958), .IN2(\s8/msel/gnt_p3 [1]), .Q(n31965) );
  OAI222X1 U35457 ( .IN1(n34223), .IN2(n31959), .IN3(n34223), .IN4(n31968), 
        .IN5(n31959), .IN6(n34228), .QN(n31963) );
  OA221X1 U35458 ( .IN1(n31963), .IN2(n31962), .IN3(n31963), .IN4(n31961), 
        .IN5(n31960), .Q(n31964) );
  NOR4X0 U35459 ( .IN1(n31966), .IN2(n31965), .IN3(n31964), .IN4(n34456), .QN(
        n31967) );
  AO221X1 U35460 ( .IN1(n31970), .IN2(n31969), .IN3(n31970), .IN4(n31968), 
        .IN5(n31967), .Q(n31980) );
  OA21X1 U35461 ( .IN1(n31972), .IN2(n31980), .IN3(n31971), .Q(n31982) );
  NAND2X0 U35462 ( .IN1(\s8/msel/gnt_p3 [1]), .IN2(n31973), .QN(n31974) );
  OA21X1 U35463 ( .IN1(n31975), .IN2(n31980), .IN3(n31974), .Q(n31979) );
  OA21X1 U35464 ( .IN1(n31977), .IN2(n31980), .IN3(n31976), .Q(n31978) );
  OA221X1 U35465 ( .IN1(\s8/msel/gnt_p3 [0]), .IN2(n31979), .IN3(n34228), 
        .IN4(n31978), .IN5(\s8/msel/gnt_p3 [2]), .Q(n31981) );
  OAI22X1 U35466 ( .IN1(n31982), .IN2(n31981), .IN3(n34223), .IN4(n31980), 
        .QN(n17808) );
  NOR2X0 U35467 ( .IN1(n31994), .IN2(n31985), .QN(n31983) );
  NOR4X0 U35468 ( .IN1(n32009), .IN2(n32011), .IN3(n31983), .IN4(n34276), .QN(
        n32001) );
  NOR2X0 U35469 ( .IN1(n31984), .IN2(n31986), .QN(n31990) );
  NAND3X0 U35470 ( .IN1(n31987), .IN2(n18196), .IN3(n34276), .QN(n31989) );
  OAI22X1 U35471 ( .IN1(n31990), .IN2(n31989), .IN3(n31988), .IN4(n32007), 
        .QN(n32000) );
  INVX0 U35472 ( .INP(n31990), .ZN(n31991) );
  OA21X1 U35473 ( .IN1(n18196), .IN2(n31992), .IN3(n31991), .Q(n31995) );
  AO22X1 U35474 ( .IN1(n31995), .IN2(n31994), .IN3(n34229), .IN4(n31993), .Q(
        n31996) );
  OA22X1 U35475 ( .IN1(n18196), .IN2(n31998), .IN3(n31997), .IN4(n31996), .Q(
        n31999) );
  AO222X1 U35476 ( .IN1(n34420), .IN2(n32001), .IN3(n34420), .IN4(n32000), 
        .IN5(n31999), .IN6(\s8/msel/gnt_p1 [2]), .Q(n32018) );
  AO21X1 U35477 ( .IN1(n32003), .IN2(n32018), .IN3(n32002), .Q(n32017) );
  INVX0 U35478 ( .INP(n32004), .ZN(n32006) );
  OA22X1 U35479 ( .IN1(n32008), .IN2(n32007), .IN3(n32006), .IN4(n32005), .Q(
        n32015) );
  INVX0 U35480 ( .INP(n32018), .ZN(n32010) );
  NOR2X0 U35481 ( .IN1(n32010), .IN2(n32009), .QN(n32013) );
  NAND2X0 U35482 ( .IN1(n32011), .IN2(n34229), .QN(n32012) );
  NAND2X0 U35483 ( .IN1(n32013), .IN2(n32012), .QN(n32014) );
  NAND3X0 U35484 ( .IN1(\s8/msel/gnt_p1 [2]), .IN2(n32015), .IN3(n32014), .QN(
        n32016) );
  AO22X1 U35485 ( .IN1(\s8/msel/gnt_p1 [1]), .IN2(n32018), .IN3(n32017), .IN4(
        n32016), .Q(n17805) );
  OA21X1 U35486 ( .IN1(n32027), .IN2(n32030), .IN3(n32025), .Q(n32021) );
  AO21X1 U35487 ( .IN1(n32025), .IN2(n32030), .IN3(n32028), .Q(n32020) );
  AO221X1 U35488 ( .IN1(\s8/msel/gnt_p0 [1]), .IN2(n32021), .IN3(n34654), 
        .IN4(n32020), .IN5(n32019), .Q(n32033) );
  NAND2X0 U35489 ( .IN1(n32023), .IN2(n32022), .QN(n32024) );
  OA221X1 U35490 ( .IN1(n32026), .IN2(n32027), .IN3(n32026), .IN4(n32025), 
        .IN5(n32024), .Q(n32032) );
  AND2X1 U35491 ( .IN1(n32028), .IN2(n32027), .Q(n32029) );
  AO221X1 U35492 ( .IN1(n32032), .IN2(n32031), .IN3(n32032), .IN4(n32030), 
        .IN5(n32029), .Q(n32037) );
  MUX21X1 U35493 ( .IN1(n32033), .IN2(n32037), .S(\s8/msel/gnt_p0 [2]), .Q(
        n32048) );
  AO21X1 U35494 ( .IN1(n32035), .IN2(n32048), .IN3(n32034), .Q(n32047) );
  NOR2X0 U35495 ( .IN1(n32036), .IN2(\s8/msel/gnt_p0 [0]), .QN(n32040) );
  NAND2X0 U35496 ( .IN1(n32038), .IN2(n32037), .QN(n32039) );
  NOR2X0 U35497 ( .IN1(n32040), .IN2(n32039), .QN(n32041) );
  NOR2X0 U35498 ( .IN1(n32041), .IN2(n34403), .QN(n32045) );
  NAND2X0 U35499 ( .IN1(n32043), .IN2(n32042), .QN(n32044) );
  NAND2X0 U35500 ( .IN1(n32045), .IN2(n32044), .QN(n32046) );
  AO22X1 U35501 ( .IN1(\s8/msel/gnt_p0 [1]), .IN2(n32048), .IN3(n32047), .IN4(
        n32046), .Q(n17802) );
  NAND3X0 U35502 ( .IN1(n13695), .IN2(m4s8_cyc), .IN3(n34369), .QN(n32091) );
  NAND3X0 U35503 ( .IN1(n13591), .IN2(m6s8_cyc), .IN3(n34580), .QN(n32100) );
  OA221X1 U35504 ( .IN1(\s8/msel/gnt_p2 [1]), .IN2(n32091), .IN3(n34273), 
        .IN4(n32100), .IN5(\s8/msel/gnt_p2 [2]), .Q(n32049) );
  NOR2X0 U35505 ( .IN1(\s8/msel/gnt_p2 [0]), .IN2(n32049), .QN(n32133) );
  NAND3X0 U35506 ( .IN1(n13539), .IN2(m7s8_cyc), .IN3(n34592), .QN(n32092) );
  NAND2X0 U35507 ( .IN1(n32100), .IN2(n32092), .QN(n32067) );
  NAND2X0 U35508 ( .IN1(n32067), .IN2(n34273), .QN(n32051) );
  NAND3X0 U35509 ( .IN1(n13916), .IN2(m0s8_cyc), .IN3(n34589), .QN(n32129) );
  INVX0 U35510 ( .INP(n32129), .ZN(n32093) );
  NAND3X0 U35511 ( .IN1(n13851), .IN2(m1s8_cyc), .IN3(n34593), .QN(n32127) );
  INVX0 U35512 ( .INP(n32127), .ZN(n32107) );
  NOR2X0 U35513 ( .IN1(n32093), .IN2(n32107), .QN(n34140) );
  NAND3X0 U35514 ( .IN1(n13747), .IN2(m3s8_cyc), .IN3(n34590), .QN(n32089) );
  INVX0 U35515 ( .INP(n32089), .ZN(n32102) );
  NAND3X0 U35516 ( .IN1(n13799), .IN2(m2s8_cyc), .IN3(n34591), .QN(n32123) );
  INVX0 U35517 ( .INP(n32123), .ZN(n32053) );
  NOR2X0 U35518 ( .IN1(n32102), .IN2(n32053), .QN(n34139) );
  NAND2X0 U35519 ( .IN1(n34140), .IN2(n34139), .QN(n32050) );
  NAND3X0 U35520 ( .IN1(n13643), .IN2(m5s8_cyc), .IN3(n34239), .QN(n32099) );
  MUX21X1 U35521 ( .IN1(n32099), .IN2(n32092), .S(\s8/msel/gnt_p2 [1]), .Q(
        n32137) );
  NAND3X0 U35522 ( .IN1(n32051), .IN2(n32050), .IN3(n32137), .QN(n32059) );
  MUX21X1 U35523 ( .IN1(n32129), .IN2(n32127), .S(\s8/msel/gnt_p2 [0]), .Q(
        n32084) );
  NOR2X0 U35524 ( .IN1(\s8/msel/gnt_p2 [1]), .IN2(n32084), .QN(n32057) );
  NAND2X0 U35525 ( .IN1(n32099), .IN2(n32091), .QN(n32052) );
  NOR2X0 U35526 ( .IN1(n32052), .IN2(n32067), .QN(n34138) );
  NAND2X0 U35527 ( .IN1(n34467), .IN2(n34273), .QN(n32114) );
  NAND2X0 U35528 ( .IN1(\s8/msel/gnt_p2 [0]), .IN2(n34273), .QN(n32061) );
  OA21X1 U35529 ( .IN1(n32107), .IN2(n32114), .IN3(n32061), .Q(n32068) );
  INVX0 U35530 ( .INP(n34139), .ZN(n32060) );
  OA22X1 U35531 ( .IN1(n32102), .IN2(n34273), .IN3(n32068), .IN4(n32060), .Q(
        n32056) );
  NAND2X0 U35532 ( .IN1(\s8/msel/gnt_p2 [0]), .IN2(\s8/msel/gnt_p2 [1]), .QN(
        n32066) );
  NOR2X0 U35533 ( .IN1(n32089), .IN2(n32066), .QN(n32131) );
  NOR2X0 U35534 ( .IN1(\s8/msel/gnt_p2 [2]), .IN2(n32131), .QN(n32055) );
  NOR2X0 U35535 ( .IN1(\s8/msel/gnt_p2 [0]), .IN2(n34273), .QN(n32096) );
  NAND2X0 U35536 ( .IN1(n32053), .IN2(n32096), .QN(n32054) );
  NAND2X0 U35537 ( .IN1(n32055), .IN2(n32054), .QN(n32085) );
  NOR4X0 U35538 ( .IN1(n32057), .IN2(n34138), .IN3(n32056), .IN4(n32085), .QN(
        n32058) );
  AO221X1 U35539 ( .IN1(\s8/msel/gnt_p2 [2]), .IN2(n32133), .IN3(
        \s8/msel/gnt_p2 [2]), .IN4(n32059), .IN5(n32058), .Q(n17800) );
  NAND2X0 U35540 ( .IN1(n32060), .IN2(n34140), .QN(n32073) );
  INVX0 U35541 ( .INP(n32100), .ZN(n32105) );
  NOR2X0 U35542 ( .IN1(n32105), .IN2(n32061), .QN(n32095) );
  NAND4X0 U35543 ( .IN1(n32099), .IN2(n32129), .IN3(n32127), .IN4(n32091), 
        .QN(n32064) );
  OA221X1 U35544 ( .IN1(n32095), .IN2(\s8/msel/gnt_p2 [1]), .IN3(n32095), 
        .IN4(n32064), .IN5(n32092), .Q(n32062) );
  NAND2X0 U35545 ( .IN1(n32073), .IN2(n32062), .QN(n32063) );
  NOR2X0 U35546 ( .IN1(n32063), .IN2(n34430), .QN(n32078) );
  NAND3X0 U35547 ( .IN1(n32099), .IN2(n32091), .IN3(n32067), .QN(n32069) );
  NAND3X0 U35548 ( .IN1(n32069), .IN2(n32064), .IN3(n32089), .QN(n32065) );
  NAND2X0 U35549 ( .IN1(n32065), .IN2(n32096), .QN(n32072) );
  INVX0 U35550 ( .INP(n32091), .ZN(n32104) );
  NOR2X0 U35551 ( .IN1(n32104), .IN2(n32066), .QN(n32117) );
  AO21X1 U35552 ( .IN1(\s8/msel/gnt_p2 [1]), .IN2(n34140), .IN3(n32067), .Q(
        n32074) );
  NAND3X0 U35553 ( .IN1(n32117), .IN2(n32099), .IN3(n32074), .QN(n32071) );
  AO21X1 U35554 ( .IN1(n34139), .IN2(n32069), .IN3(n32068), .Q(n32070) );
  NAND4X0 U35555 ( .IN1(n34430), .IN2(n32072), .IN3(n32071), .IN4(n32070), 
        .QN(n32083) );
  INVX0 U35556 ( .INP(n32073), .ZN(n32075) );
  AO221X1 U35557 ( .IN1(n32099), .IN2(n32075), .IN3(n32099), .IN4(n32074), 
        .IN5(n32114), .Q(n32076) );
  NAND2X0 U35558 ( .IN1(n32083), .IN2(n32076), .QN(n32077) );
  NOR2X0 U35559 ( .IN1(n32078), .IN2(n32077), .QN(n32088) );
  INVX0 U35560 ( .INP(n32099), .ZN(n32079) );
  NAND2X0 U35561 ( .IN1(\s8/msel/gnt_p2 [2]), .IN2(\s8/msel/gnt_p2 [0]), .QN(
        n32136) );
  NOR2X0 U35562 ( .IN1(n32079), .IN2(n32136), .QN(n32087) );
  NAND2X0 U35563 ( .IN1(n32096), .IN2(n32105), .QN(n32081) );
  NAND3X0 U35564 ( .IN1(n32088), .IN2(n34467), .IN3(n32091), .QN(n32080) );
  NAND3X0 U35565 ( .IN1(n32081), .IN2(n32080), .IN3(\s8/msel/gnt_p2 [2]), .QN(
        n32082) );
  OA221X1 U35566 ( .IN1(n32085), .IN2(n32084), .IN3(n32085), .IN4(n32083), 
        .IN5(n32082), .Q(n32086) );
  AO221X1 U35567 ( .IN1(n32088), .IN2(\s8/msel/gnt_p2 [1]), .IN3(n32088), 
        .IN4(n32087), .IN5(n32086), .Q(n17799) );
  OA21X1 U35568 ( .IN1(n32104), .IN2(n32099), .IN3(n32089), .Q(n32106) );
  NAND2X0 U35569 ( .IN1(n32129), .IN2(n32123), .QN(n32090) );
  NOR2X0 U35570 ( .IN1(n32106), .IN2(n32090), .QN(n32098) );
  INVX0 U35571 ( .INP(n32090), .ZN(n32101) );
  NAND3X0 U35572 ( .IN1(\s8/msel/gnt_p2 [0]), .IN2(n32101), .IN3(n32091), .QN(
        n32094) );
  OA21X1 U35573 ( .IN1(n32093), .IN2(n32127), .IN3(n32092), .Q(n32111) );
  NAND2X0 U35574 ( .IN1(n32094), .IN2(n32111), .QN(n32097) );
  OA22X1 U35575 ( .IN1(n32098), .IN2(n32097), .IN3(n32096), .IN4(n32095), .Q(
        n32126) );
  OA21X1 U35576 ( .IN1(n32105), .IN2(n32111), .IN3(n32099), .Q(n32115) );
  NAND3X0 U35577 ( .IN1(n32102), .IN2(n32101), .IN3(n32100), .QN(n32103) );
  AO21X1 U35578 ( .IN1(n32115), .IN2(n32103), .IN3(n32114), .Q(n32110) );
  NOR2X0 U35579 ( .IN1(n32105), .IN2(n32104), .QN(n32112) );
  AND2X1 U35580 ( .IN1(\s8/msel/gnt_p2 [0]), .IN2(n32112), .Q(n32108) );
  INVX0 U35581 ( .INP(n32106), .ZN(n32122) );
  AO221X1 U35582 ( .IN1(n32123), .IN2(n32108), .IN3(n32123), .IN4(n32122), 
        .IN5(n32107), .Q(n32118) );
  NAND3X0 U35583 ( .IN1(\s8/msel/gnt_p2 [1]), .IN2(n32118), .IN3(n32129), .QN(
        n32109) );
  NAND3X0 U35584 ( .IN1(\s8/msel/gnt_p2 [2]), .IN2(n32110), .IN3(n32109), .QN(
        n32125) );
  INVX0 U35585 ( .INP(n32111), .ZN(n32113) );
  OA221X1 U35586 ( .IN1(n32113), .IN2(\s8/msel/gnt_p2 [0]), .IN3(n32113), 
        .IN4(n32129), .IN5(n32112), .Q(n32121) );
  INVX0 U35587 ( .INP(n32114), .ZN(n32119) );
  INVX0 U35588 ( .INP(n32115), .ZN(n32116) );
  AO22X1 U35589 ( .IN1(n32119), .IN2(n32118), .IN3(n32117), .IN4(n32116), .Q(
        n32120) );
  AO221X1 U35590 ( .IN1(n32123), .IN2(n32122), .IN3(n32123), .IN4(n32121), 
        .IN5(n32120), .Q(n32124) );
  OA22X1 U35591 ( .IN1(n32126), .IN2(n32125), .IN3(\s8/msel/gnt_p2 [2]), .IN4(
        n32124), .Q(n32132) );
  NOR2X0 U35592 ( .IN1(n34467), .IN2(n32127), .QN(n32128) );
  AO222X1 U35593 ( .IN1(n32132), .IN2(\s8/msel/gnt_p2 [1]), .IN3(n32132), 
        .IN4(n32129), .IN5(n34273), .IN6(n32128), .Q(n32130) );
  NOR2X0 U35594 ( .IN1(n32131), .IN2(n32130), .QN(n32135) );
  INVX0 U35595 ( .INP(n32132), .ZN(n32134) );
  OAI222X1 U35596 ( .IN1(n32137), .IN2(n32136), .IN3(\s8/msel/gnt_p2 [2]), 
        .IN4(n32135), .IN5(n32134), .IN6(n32133), .QN(n17798) );
  NOR2X0 U35597 ( .IN1(n32138), .IN2(n34379), .QN(n32139) );
  MUX21X1 U35598 ( .IN1(n34321), .IN2(s15_data_o[0]), .S(n32139), .Q(n17797)
         );
  MUX21X1 U35599 ( .IN1(n34502), .IN2(s15_data_o[1]), .S(n32139), .Q(n17796)
         );
  MUX21X1 U35600 ( .IN1(n34618), .IN2(s15_data_o[2]), .S(n32139), .Q(n17795)
         );
  MUX21X1 U35601 ( .IN1(n34581), .IN2(s15_data_o[3]), .S(n32139), .Q(n17794)
         );
  MUX21X1 U35602 ( .IN1(n34352), .IN2(s15_data_o[4]), .S(n32139), .Q(n17793)
         );
  MUX21X1 U35603 ( .IN1(n34535), .IN2(s15_data_o[5]), .S(n32139), .Q(n17792)
         );
  MUX21X1 U35604 ( .IN1(n34636), .IN2(s15_data_o[6]), .S(n32139), .Q(n17791)
         );
  MUX21X1 U35605 ( .IN1(n34596), .IN2(s15_data_o[7]), .S(n32139), .Q(n17790)
         );
  MUX21X1 U35606 ( .IN1(n34319), .IN2(s15_data_o[8]), .S(n32139), .Q(n17789)
         );
  MUX21X1 U35607 ( .IN1(n34536), .IN2(s15_data_o[9]), .S(n32139), .Q(n17788)
         );
  MUX21X1 U35608 ( .IN1(n34351), .IN2(s15_data_o[10]), .S(n32139), .Q(n17787)
         );
  MUX21X1 U35609 ( .IN1(n34501), .IN2(s15_data_o[11]), .S(n32139), .Q(n17786)
         );
  MUX21X1 U35610 ( .IN1(n34320), .IN2(s15_data_o[12]), .S(n32139), .Q(n17785)
         );
  MUX21X1 U35611 ( .IN1(n34500), .IN2(s15_data_o[13]), .S(n32139), .Q(n17784)
         );
  MUX21X1 U35612 ( .IN1(n34364), .IN2(s15_data_o[14]), .S(n32139), .Q(n17783)
         );
  MUX21X1 U35613 ( .IN1(n34603), .IN2(s15_data_o[15]), .S(n32139), .Q(n17782)
         );
  NAND3X0 U35614 ( .IN1(m0s9_cyc), .IN2(n34321), .IN3(n34502), .QN(n32196) );
  INVX0 U35615 ( .INP(n32196), .ZN(n32220) );
  NAND2X0 U35616 ( .IN1(m1s9_cyc), .IN2(n34581), .QN(n32140) );
  NOR2X0 U35617 ( .IN1(n13852), .IN2(n32140), .QN(n32177) );
  MUX21X1 U35618 ( .IN1(n32220), .IN2(n32177), .S(\s9/msel/gnt_p3 [0]), .Q(
        n32169) );
  NAND3X0 U35619 ( .IN1(m2s9_cyc), .IN2(n34352), .IN3(n34535), .QN(n32186) );
  NAND2X0 U35620 ( .IN1(\s9/msel/gnt_p3 [1]), .IN2(n32186), .QN(n32142) );
  NOR2X0 U35621 ( .IN1(n34282), .IN2(n34225), .QN(n32210) );
  INVX0 U35622 ( .INP(n32210), .ZN(n32141) );
  OA221X1 U35623 ( .IN1(n32169), .IN2(\s9/msel/gnt_p3 [1]), .IN3(n32142), 
        .IN4(\s9/msel/gnt_p3 [0]), .IN5(n32141), .Q(n32146) );
  NAND2X0 U35624 ( .IN1(m3s9_cyc), .IN2(n34596), .QN(n32143) );
  NOR2X0 U35625 ( .IN1(n13748), .IN2(n32143), .QN(n32195) );
  INVX0 U35626 ( .INP(n32195), .ZN(n32180) );
  NAND2X0 U35627 ( .IN1(n32186), .IN2(n32180), .QN(n32164) );
  NOR2X0 U35628 ( .IN1(\s9/msel/gnt_p3 [1]), .IN2(n34282), .QN(n32217) );
  NAND2X0 U35629 ( .IN1(n32217), .IN2(n32186), .QN(n32201) );
  AO21X1 U35630 ( .IN1(n34225), .IN2(n32201), .IN3(n32195), .Q(n32144) );
  OA21X1 U35631 ( .IN1(n32177), .IN2(n32164), .IN3(n32144), .Q(n32145) );
  NOR2X0 U35632 ( .IN1(n32146), .IN2(n32145), .QN(n32150) );
  NAND3X0 U35633 ( .IN1(m4s9_cyc), .IN2(n34319), .IN3(n34536), .QN(n32188) );
  INVX0 U35634 ( .INP(n32188), .ZN(n32179) );
  NAND3X0 U35635 ( .IN1(m5s9_cyc), .IN2(n34351), .IN3(n34501), .QN(n32174) );
  INVX0 U35636 ( .INP(n32174), .ZN(n32207) );
  NOR2X0 U35637 ( .IN1(n32179), .IN2(n32207), .QN(n32156) );
  NAND3X0 U35638 ( .IN1(m6s9_cyc), .IN2(n34320), .IN3(n34500), .QN(n32187) );
  NAND3X0 U35639 ( .IN1(m7s9_cyc), .IN2(n34364), .IN3(n34603), .QN(n32189) );
  AND2X1 U35640 ( .IN1(n32187), .IN2(n32189), .Q(n32151) );
  NAND2X0 U35641 ( .IN1(n32156), .IN2(n32151), .QN(n34158) );
  INVX0 U35642 ( .INP(n32187), .ZN(n32181) );
  MUX21X1 U35643 ( .IN1(n32179), .IN2(n32181), .S(\s9/msel/gnt_p3 [1]), .Q(
        n32216) );
  NAND2X0 U35644 ( .IN1(n32216), .IN2(n34282), .QN(n32148) );
  AO22X1 U35645 ( .IN1(\s9/msel/gnt_p3 [1]), .IN2(n32189), .IN3(n32151), .IN4(
        n32174), .Q(n32147) );
  INVX0 U35646 ( .INP(n32177), .ZN(n32219) );
  NAND2X0 U35647 ( .IN1(n32196), .IN2(n32219), .QN(n32152) );
  OR2X1 U35648 ( .IN1(n32152), .IN2(n32164), .Q(n34159) );
  NAND3X0 U35649 ( .IN1(n32148), .IN2(n32147), .IN3(n34159), .QN(n32149) );
  OA222X1 U35650 ( .IN1(\s9/msel/gnt_p3 [2]), .IN2(n32150), .IN3(
        \s9/msel/gnt_p3 [2]), .IN4(n34158), .IN5(n34560), .IN6(n32149), .Q(
        n17781) );
  NOR2X0 U35651 ( .IN1(n34225), .IN2(n32189), .QN(n32175) );
  NAND2X0 U35652 ( .IN1(n34225), .IN2(n32207), .QN(n32185) );
  AO21X1 U35653 ( .IN1(\s9/msel/gnt_p3 [1]), .IN2(n32156), .IN3(n32164), .Q(
        n32159) );
  NAND4X0 U35654 ( .IN1(n32196), .IN2(n32219), .IN3(n32185), .IN4(n32159), 
        .QN(n32155) );
  OA21X1 U35655 ( .IN1(n34225), .IN2(n32152), .IN3(n32151), .Q(n32158) );
  NOR2X0 U35656 ( .IN1(n32158), .IN2(\s9/msel/gnt_p3 [1]), .QN(n32153) );
  NAND2X0 U35657 ( .IN1(n32153), .IN2(n32174), .QN(n32154) );
  NAND3X0 U35658 ( .IN1(\s9/msel/gnt_p3 [2]), .IN2(n32155), .IN3(n32154), .QN(
        n32166) );
  NOR2X0 U35659 ( .IN1(\s9/msel/gnt_p3 [0]), .IN2(n34225), .QN(n32163) );
  INVX0 U35660 ( .INP(n32156), .ZN(n32157) );
  NOR2X0 U35661 ( .IN1(n32158), .IN2(n32157), .QN(n32161) );
  AND2X1 U35662 ( .IN1(n32159), .IN2(n34225), .Q(n32160) );
  OA22X1 U35663 ( .IN1(n32161), .IN2(n32160), .IN3(n32219), .IN4(
        \s9/msel/gnt_p3 [1]), .Q(n32162) );
  AO221X1 U35664 ( .IN1(n32164), .IN2(n32217), .IN3(n32164), .IN4(n32163), 
        .IN5(n32162), .Q(n32165) );
  OA22X1 U35665 ( .IN1(n32175), .IN2(n32166), .IN3(\s9/msel/gnt_p3 [2]), .IN4(
        n32165), .Q(n32168) );
  AO22X1 U35666 ( .IN1(\s9/msel/gnt_p3 [1]), .IN2(n32181), .IN3(n32168), .IN4(
        n32188), .Q(n32167) );
  NAND3X0 U35667 ( .IN1(\s9/msel/gnt_p3 [2]), .IN2(n34282), .IN3(n32167), .QN(
        n32173) );
  NAND2X0 U35668 ( .IN1(n32195), .IN2(n32210), .QN(n32223) );
  INVX0 U35669 ( .INP(n32168), .ZN(n32170) );
  AO221X1 U35670 ( .IN1(n32223), .IN2(n32170), .IN3(n32223), .IN4(n32169), 
        .IN5(\s9/msel/gnt_p3 [2]), .Q(n32172) );
  NAND2X0 U35671 ( .IN1(\s9/msel/gnt_p3 [0]), .IN2(\s9/msel/gnt_p3 [2]), .QN(
        n32230) );
  AO21X1 U35672 ( .IN1(n34225), .IN2(n32230), .IN3(n32170), .Q(n32171) );
  NAND3X0 U35673 ( .IN1(n32173), .IN2(n32172), .IN3(n32171), .QN(n17780) );
  NOR2X0 U35674 ( .IN1(\s9/msel/gnt_p3 [1]), .IN2(n32174), .QN(n32176) );
  NOR2X0 U35675 ( .IN1(n32176), .IN2(n32175), .QN(n32229) );
  OA221X1 U35676 ( .IN1(n32207), .IN2(\s9/msel/gnt_p3 [0]), .IN3(n32207), 
        .IN4(n32187), .IN5(n32188), .Q(n32208) );
  AO221X1 U35677 ( .IN1(n32186), .IN2(n32195), .IN3(n32186), .IN4(n32208), 
        .IN5(n32177), .Q(n32190) );
  NAND3X0 U35678 ( .IN1(\s9/msel/gnt_p3 [1]), .IN2(n32190), .IN3(n32196), .QN(
        n32184) );
  OA21X1 U35679 ( .IN1(n32220), .IN2(n32219), .IN3(n32189), .Q(n32194) );
  NOR2X0 U35680 ( .IN1(\s9/msel/gnt_p3 [0]), .IN2(n32207), .QN(n32178) );
  NAND2X0 U35681 ( .IN1(n32196), .IN2(n32186), .QN(n32204) );
  AO221X1 U35682 ( .IN1(n32180), .IN2(n32179), .IN3(n32180), .IN4(n32178), 
        .IN5(n32204), .Q(n32182) );
  AO21X1 U35683 ( .IN1(n32194), .IN2(n32182), .IN3(n32181), .Q(n32183) );
  NAND4X0 U35684 ( .IN1(\s9/msel/gnt_p3 [2]), .IN2(n32185), .IN3(n32184), 
        .IN4(n32183), .QN(n32215) );
  INVX0 U35685 ( .INP(n32186), .ZN(n32221) );
  NAND2X0 U35686 ( .IN1(n32188), .IN2(n32187), .QN(n32193) );
  OR2X1 U35687 ( .IN1(n32189), .IN2(n32193), .Q(n32202) );
  INVX0 U35688 ( .INP(n32190), .ZN(n32191) );
  OA21X1 U35689 ( .IN1(n32221), .IN2(n32202), .IN3(n32191), .Q(n32192) );
  NOR2X0 U35690 ( .IN1(n32192), .IN2(\s9/msel/gnt_p3 [0]), .QN(n32199) );
  NOR2X0 U35691 ( .IN1(n32194), .IN2(n32193), .QN(n32205) );
  AO221X1 U35692 ( .IN1(n32208), .IN2(n32207), .IN3(n32208), .IN4(n32196), 
        .IN5(n32195), .Q(n32200) );
  NOR2X0 U35693 ( .IN1(n32205), .IN2(n32200), .QN(n32197) );
  NAND2X0 U35694 ( .IN1(\s9/msel/gnt_p3 [1]), .IN2(n32197), .QN(n32198) );
  NAND2X0 U35695 ( .IN1(n32199), .IN2(n32198), .QN(n32213) );
  INVX0 U35696 ( .INP(n32200), .ZN(n32203) );
  AO21X1 U35697 ( .IN1(n32203), .IN2(n32202), .IN3(n32201), .Q(n32212) );
  INVX0 U35698 ( .INP(n32204), .ZN(n32206) );
  AO221X1 U35699 ( .IN1(n32208), .IN2(n32207), .IN3(n32208), .IN4(n32206), 
        .IN5(n32205), .Q(n32209) );
  NAND2X0 U35700 ( .IN1(n32210), .IN2(n32209), .QN(n32211) );
  NAND4X0 U35701 ( .IN1(n32213), .IN2(n34560), .IN3(n32212), .IN4(n32211), 
        .QN(n32214) );
  NAND2X0 U35702 ( .IN1(n32215), .IN2(n32214), .QN(n32228) );
  OA21X1 U35703 ( .IN1(n34560), .IN2(n32216), .IN3(n34282), .Q(n32227) );
  INVX0 U35704 ( .INP(n32217), .ZN(n32218) );
  NOR2X0 U35705 ( .IN1(n32219), .IN2(n32218), .QN(n32225) );
  AO221X1 U35706 ( .IN1(\s9/msel/gnt_p3 [1]), .IN2(n32221), .IN3(n34225), 
        .IN4(n32220), .IN5(n32228), .Q(n32222) );
  NAND2X0 U35707 ( .IN1(n32223), .IN2(n32222), .QN(n32224) );
  NOR2X0 U35708 ( .IN1(n32225), .IN2(n32224), .QN(n32226) );
  OAI222X1 U35709 ( .IN1(n32230), .IN2(n32229), .IN3(n32228), .IN4(n32227), 
        .IN5(n32226), .IN6(\s9/msel/gnt_p3 [2]), .QN(n17779) );
  NAND2X0 U35710 ( .IN1(n32231), .IN2(n34260), .QN(n32236) );
  NOR2X0 U35711 ( .IN1(n32233), .IN2(n32232), .QN(n32249) );
  AO21X1 U35712 ( .IN1(n32249), .IN2(n32234), .IN3(n32256), .Q(n32235) );
  NAND2X0 U35713 ( .IN1(n32237), .IN2(n32250), .QN(n32254) );
  INVX0 U35714 ( .INP(n32254), .ZN(n32248) );
  NAND2X0 U35715 ( .IN1(n32239), .IN2(n32238), .QN(n32257) );
  INVX0 U35716 ( .INP(n32257), .ZN(n32255) );
  NAND2X0 U35717 ( .IN1(n32248), .IN2(n32255), .QN(n34156) );
  NAND3X0 U35718 ( .IN1(n32236), .IN2(n32235), .IN3(n34156), .QN(n32247) );
  NAND2X0 U35719 ( .IN1(\s9/msel/gnt_p1 [1]), .IN2(n34260), .QN(n32266) );
  OA21X1 U35720 ( .IN1(n32237), .IN2(n32266), .IN3(n34442), .Q(n32263) );
  NOR2X0 U35721 ( .IN1(\s9/msel/gnt_p1 [0]), .IN2(n32238), .QN(n32264) );
  NAND2X0 U35722 ( .IN1(n34400), .IN2(n32239), .QN(n32252) );
  NOR3X0 U35723 ( .IN1(n32264), .IN2(n32252), .IN3(n32254), .QN(n32240) );
  NOR2X0 U35724 ( .IN1(\s9/msel/gnt_p1 [1]), .IN2(n32240), .QN(n32245) );
  NAND2X0 U35725 ( .IN1(n32242), .IN2(n32241), .QN(n32258) );
  INVX0 U35726 ( .INP(n32258), .ZN(n32243) );
  NAND2X0 U35727 ( .IN1(n32249), .IN2(n32243), .QN(n34157) );
  NAND2X0 U35728 ( .IN1(n34157), .IN2(n32250), .QN(n32244) );
  NOR2X0 U35729 ( .IN1(n32245), .IN2(n32244), .QN(n32246) );
  AO22X1 U35730 ( .IN1(\s9/msel/gnt_p1 [2]), .IN2(n32247), .IN3(n32263), .IN4(
        n32246), .Q(n17778) );
  OA21X1 U35731 ( .IN1(n32249), .IN2(n32258), .IN3(n32248), .Q(n32253) );
  OA21X1 U35732 ( .IN1(n34400), .IN2(n32257), .IN3(n32249), .Q(n32259) );
  OA21X1 U35733 ( .IN1(n32259), .IN2(n32258), .IN3(n32250), .Q(n32251) );
  OA22X1 U35734 ( .IN1(n32253), .IN2(n32252), .IN3(n32251), .IN4(n34400), .Q(
        n32262) );
  NAND2X0 U35735 ( .IN1(n32255), .IN2(n32254), .QN(n32261) );
  OA21X1 U35736 ( .IN1(n32258), .IN2(n32257), .IN3(n32256), .Q(n32260) );
  AO221X1 U35737 ( .IN1(n32261), .IN2(n32260), .IN3(n32261), .IN4(n32259), 
        .IN5(n34442), .Q(n32267) );
  OA21X1 U35738 ( .IN1(\s9/msel/gnt_p1 [2]), .IN2(n32262), .IN3(n32267), .Q(
        n32277) );
  OA21X1 U35739 ( .IN1(n32277), .IN2(n32264), .IN3(n32263), .Q(n32276) );
  NOR2X0 U35740 ( .IN1(n32266), .IN2(n32265), .QN(n32274) );
  NOR2X0 U35741 ( .IN1(n32268), .IN2(n32267), .QN(n32271) );
  NAND2X0 U35742 ( .IN1(n32269), .IN2(n34260), .QN(n32270) );
  NAND2X0 U35743 ( .IN1(n32271), .IN2(n32270), .QN(n32272) );
  NAND2X0 U35744 ( .IN1(n32272), .IN2(\s9/msel/gnt_p1 [2]), .QN(n32273) );
  NOR2X0 U35745 ( .IN1(n32274), .IN2(n32273), .QN(n32275) );
  OAI22X1 U35746 ( .IN1(n32277), .IN2(n34400), .IN3(n32276), .IN4(n32275), 
        .QN(n17777) );
  NAND3X0 U35747 ( .IN1(n13592), .IN2(n13566), .IN3(m6s9_cyc), .QN(n32346) );
  NAND3X0 U35748 ( .IN1(n13540), .IN2(n13490), .IN3(m7s9_cyc), .QN(n32318) );
  AND2X1 U35749 ( .IN1(n32346), .IN2(n32318), .Q(n32302) );
  NAND3X0 U35750 ( .IN1(n13644), .IN2(n13618), .IN3(m5s9_cyc), .QN(n32321) );
  NAND2X0 U35751 ( .IN1(n32302), .IN2(n32321), .QN(n32279) );
  NAND2X0 U35752 ( .IN1(\s9/msel/gnt_p0 [1]), .IN2(n32318), .QN(n32282) );
  NAND4X0 U35753 ( .IN1(\s9/msel/gnt_p0 [0]), .IN2(n32346), .IN3(n34266), 
        .IN4(n32318), .QN(n32292) );
  NAND2X0 U35754 ( .IN1(n32282), .IN2(n32292), .QN(n32295) );
  INVX0 U35755 ( .INP(n32295), .ZN(n32278) );
  NAND3X0 U35756 ( .IN1(n13696), .IN2(n13670), .IN3(m4s9_cyc), .QN(n32345) );
  INVX0 U35757 ( .INP(n32345), .ZN(n32341) );
  INVX0 U35758 ( .INP(n32346), .ZN(n32319) );
  MUX21X1 U35759 ( .IN1(n32341), .IN2(n32319), .S(\s9/msel/gnt_p0 [1]), .Q(
        n32362) );
  NAND3X0 U35760 ( .IN1(n13800), .IN2(n13774), .IN3(m2s9_cyc), .QN(n32325) );
  INVX0 U35761 ( .INP(n32325), .ZN(n32347) );
  AND3X1 U35762 ( .IN1(n13748), .IN2(n13722), .IN3(m3s9_cyc), .Q(n32331) );
  NOR2X0 U35763 ( .IN1(n32347), .IN2(n32331), .QN(n32300) );
  NAND3X0 U35764 ( .IN1(n13918), .IN2(n13878), .IN3(m0s9_cyc), .QN(n32326) );
  NAND3X0 U35765 ( .IN1(n13852), .IN2(n13826), .IN3(m1s9_cyc), .QN(n32359) );
  NAND2X0 U35766 ( .IN1(n32326), .IN2(n32359), .QN(n32301) );
  INVX0 U35767 ( .INP(n32301), .ZN(n32291) );
  AO222X1 U35768 ( .IN1(n32279), .IN2(n32278), .IN3(n34436), .IN4(n32362), 
        .IN5(n32300), .IN6(n32291), .Q(n32280) );
  NAND2X0 U35769 ( .IN1(\s9/msel/gnt_p0 [2]), .IN2(n32280), .QN(n32290) );
  NAND2X0 U35770 ( .IN1(n34266), .IN2(n32321), .QN(n32281) );
  NAND4X0 U35771 ( .IN1(\s9/msel/gnt_p0 [2]), .IN2(\s9/msel/gnt_p0 [0]), .IN3(
        n32282), .IN4(n32281), .QN(n32364) );
  NOR2X0 U35772 ( .IN1(\s9/msel/gnt_p0 [0]), .IN2(n34266), .QN(n32334) );
  INVX0 U35773 ( .INP(n32334), .ZN(n32312) );
  NOR2X0 U35774 ( .IN1(n32312), .IN2(n32325), .QN(n32284) );
  NOR2X0 U35775 ( .IN1(n34436), .IN2(n34266), .QN(n32327) );
  NAND2X0 U35776 ( .IN1(n32331), .IN2(n32327), .QN(n32356) );
  NAND2X0 U35777 ( .IN1(n32356), .IN2(n34284), .QN(n32283) );
  NOR2X0 U35778 ( .IN1(n32284), .IN2(n32283), .QN(n32309) );
  INVX0 U35779 ( .INP(n32326), .ZN(n32357) );
  INVX0 U35780 ( .INP(n32359), .ZN(n32323) );
  MUX21X1 U35781 ( .IN1(n32357), .IN2(n32323), .S(\s9/msel/gnt_p0 [0]), .Q(
        n32310) );
  NAND2X0 U35782 ( .IN1(n34266), .IN2(n32310), .QN(n32288) );
  NAND2X0 U35783 ( .IN1(n32321), .IN2(n32345), .QN(n32299) );
  INVX0 U35784 ( .INP(n32299), .ZN(n32304) );
  NAND2X0 U35785 ( .IN1(n32302), .IN2(n32304), .QN(n32287) );
  OR2X1 U35786 ( .IN1(\s9/msel/gnt_p0 [1]), .IN2(n32323), .Q(n32298) );
  INVX0 U35787 ( .INP(n32300), .ZN(n32293) );
  OA22X1 U35788 ( .IN1(n32331), .IN2(n32312), .IN3(n32298), .IN4(n32293), .Q(
        n32285) );
  INVX0 U35789 ( .INP(n32327), .ZN(n32342) );
  NAND2X0 U35790 ( .IN1(n32285), .IN2(n32342), .QN(n32286) );
  NAND4X0 U35791 ( .IN1(n32309), .IN2(n32288), .IN3(n32287), .IN4(n32286), 
        .QN(n32289) );
  NAND3X0 U35792 ( .IN1(n32290), .IN2(n32364), .IN3(n32289), .QN(n17775) );
  NOR2X0 U35793 ( .IN1(\s9/msel/gnt_p0 [0]), .IN2(\s9/msel/gnt_p0 [1]), .QN(
        n32339) );
  INVX0 U35794 ( .INP(n32321), .ZN(n32328) );
  AO221X1 U35795 ( .IN1(n32302), .IN2(n32300), .IN3(n32302), .IN4(n32301), 
        .IN5(n32328), .Q(n32296) );
  OAI221X1 U35796 ( .IN1(n32293), .IN2(n32292), .IN3(n32293), .IN4(n32304), 
        .IN5(n32291), .QN(n32294) );
  AO22X1 U35797 ( .IN1(n32339), .IN2(n32296), .IN3(n32295), .IN4(n32294), .Q(
        n32297) );
  NAND2X0 U35798 ( .IN1(\s9/msel/gnt_p0 [2]), .IN2(n32297), .QN(n32311) );
  AO221X1 U35799 ( .IN1(n32300), .IN2(n32302), .IN3(n32300), .IN4(n32299), 
        .IN5(n32298), .Q(n32307) );
  NAND2X0 U35800 ( .IN1(n32302), .IN2(n32301), .QN(n32303) );
  NAND3X0 U35801 ( .IN1(\s9/msel/gnt_p0 [1]), .IN2(n32304), .IN3(n32303), .QN(
        n32306) );
  NAND2X0 U35802 ( .IN1(n32331), .IN2(n32334), .QN(n32305) );
  NAND4X0 U35803 ( .IN1(n34284), .IN2(n32307), .IN3(n32306), .IN4(n32305), 
        .QN(n32308) );
  NAND2X0 U35804 ( .IN1(n32311), .IN2(n32308), .QN(n32315) );
  OA21X1 U35805 ( .IN1(n32315), .IN2(n32310), .IN3(n32309), .Q(n32317) );
  INVX0 U35806 ( .INP(n32311), .ZN(n32314) );
  OA221X1 U35807 ( .IN1(\s9/msel/gnt_p0 [0]), .IN2(n32341), .IN3(n34436), 
        .IN4(n32328), .IN5(\s9/msel/gnt_p0 [2]), .Q(n32313) );
  OA22X1 U35808 ( .IN1(n32314), .IN2(n32313), .IN3(n32346), .IN4(n32312), .Q(
        n32316) );
  OAI22X1 U35809 ( .IN1(n32317), .IN2(n32316), .IN3(n34266), .IN4(n32315), 
        .QN(n17774) );
  INVX0 U35810 ( .INP(n32339), .ZN(n32320) );
  OA21X1 U35811 ( .IN1(n32357), .IN2(n32359), .IN3(n32318), .Q(n32349) );
  OA21X1 U35812 ( .IN1(n32319), .IN2(n32349), .IN3(n32321), .Q(n32340) );
  OR2X1 U35813 ( .IN1(n32320), .IN2(n32340), .Q(n32337) );
  NOR2X0 U35814 ( .IN1(n32341), .IN2(n32321), .QN(n32322) );
  NOR2X0 U35815 ( .IN1(n32331), .IN2(n32322), .QN(n32343) );
  AO21X1 U35816 ( .IN1(n32325), .IN2(n32324), .IN3(n32323), .Q(n32338) );
  NAND3X0 U35817 ( .IN1(n32327), .IN2(n32326), .IN3(n32338), .QN(n32336) );
  OA21X1 U35818 ( .IN1(\s9/msel/gnt_p0 [0]), .IN2(n32328), .IN3(n32345), .Q(
        n32330) );
  NOR2X0 U35819 ( .IN1(n32357), .IN2(n32347), .QN(n32329) );
  OA21X1 U35820 ( .IN1(n32331), .IN2(n32330), .IN3(n32329), .Q(n32333) );
  INVX0 U35821 ( .INP(n32349), .ZN(n32332) );
  OAI22X1 U35822 ( .IN1(n32346), .IN2(n32334), .IN3(n32333), .IN4(n32332), 
        .QN(n32335) );
  NAND4X0 U35823 ( .IN1(\s9/msel/gnt_p0 [2]), .IN2(n32337), .IN3(n32336), 
        .IN4(n32335), .QN(n32355) );
  NAND2X0 U35824 ( .IN1(n32339), .IN2(n32338), .QN(n32353) );
  OR3X1 U35825 ( .IN1(n32342), .IN2(n32341), .IN3(n32340), .Q(n32352) );
  NAND3X0 U35826 ( .IN1(\s9/msel/gnt_p0 [0]), .IN2(n32346), .IN3(n32345), .QN(
        n32344) );
  OA21X1 U35827 ( .IN1(n32357), .IN2(n32344), .IN3(n32343), .Q(n32350) );
  NAND2X0 U35828 ( .IN1(n32346), .IN2(n32345), .QN(n32348) );
  AO221X1 U35829 ( .IN1(n32350), .IN2(n32349), .IN3(n32350), .IN4(n32348), 
        .IN5(n32347), .Q(n32351) );
  NAND4X0 U35830 ( .IN1(n34284), .IN2(n32353), .IN3(n32352), .IN4(n32351), 
        .QN(n32354) );
  NAND2X0 U35831 ( .IN1(n32355), .IN2(n32354), .QN(n32361) );
  OA221X1 U35832 ( .IN1(n32361), .IN2(n32357), .IN3(n32361), .IN4(n34266), 
        .IN5(n32356), .Q(n32360) );
  NAND2X0 U35833 ( .IN1(\s9/msel/gnt_p0 [0]), .IN2(n34266), .QN(n32358) );
  AO221X1 U35834 ( .IN1(n32360), .IN2(n32359), .IN3(n32360), .IN4(n32358), 
        .IN5(\s9/msel/gnt_p0 [2]), .Q(n32365) );
  AO221X1 U35835 ( .IN1(n34436), .IN2(n34284), .IN3(n34436), .IN4(n32362), 
        .IN5(n32361), .Q(n32363) );
  NAND3X0 U35836 ( .IN1(n32365), .IN2(n32364), .IN3(n32363), .QN(n17773) );
  NAND3X0 U35837 ( .IN1(n13592), .IN2(m6s9_cyc), .IN3(n34500), .QN(n32411) );
  INVX0 U35838 ( .INP(n32411), .ZN(n32435) );
  AND3X1 U35839 ( .IN1(n13540), .IN2(m7s9_cyc), .IN3(n34603), .Q(n32414) );
  NOR2X0 U35840 ( .IN1(n32435), .IN2(n32414), .QN(n34154) );
  INVX0 U35841 ( .INP(n34154), .ZN(n32382) );
  NAND3X0 U35842 ( .IN1(n13644), .IN2(m5s9_cyc), .IN3(n34501), .QN(n32421) );
  INVX0 U35843 ( .INP(n32421), .ZN(n32410) );
  NOR2X0 U35844 ( .IN1(n32382), .IN2(n32410), .QN(n32366) );
  NAND2X0 U35845 ( .IN1(\s9/msel/gnt_p2 [1]), .IN2(n34462), .QN(n32391) );
  NOR2X0 U35846 ( .IN1(n32414), .IN2(n32391), .QN(n32377) );
  NAND2X0 U35847 ( .IN1(\s9/msel/gnt_p2 [0]), .IN2(\s9/msel/gnt_p2 [1]), .QN(
        n32388) );
  INVX0 U35848 ( .INP(n32388), .ZN(n32428) );
  NOR3X0 U35849 ( .IN1(n32366), .IN2(n32377), .IN3(n32428), .QN(n32368) );
  NAND3X0 U35850 ( .IN1(n13918), .IN2(m0s9_cyc), .IN3(n34502), .QN(n32446) );
  NAND3X0 U35851 ( .IN1(n13852), .IN2(m1s9_cyc), .IN3(n34581), .QN(n32369) );
  NAND2X0 U35852 ( .IN1(n32446), .IN2(n32369), .QN(n32378) );
  NAND3X0 U35853 ( .IN1(n13800), .IN2(m2s9_cyc), .IN3(n34535), .QN(n32444) );
  NAND3X0 U35854 ( .IN1(n13748), .IN2(m3s9_cyc), .IN3(n34596), .QN(n32433) );
  NAND2X0 U35855 ( .IN1(n32444), .IN2(n32433), .QN(n32380) );
  NOR2X0 U35856 ( .IN1(n32378), .IN2(n32380), .QN(n34152) );
  NAND3X0 U35857 ( .IN1(n13696), .IN2(m4s9_cyc), .IN3(n34536), .QN(n32422) );
  MUX21X1 U35858 ( .IN1(n32422), .IN2(n32411), .S(\s9/msel/gnt_p2 [1]), .Q(
        n32452) );
  NOR2X0 U35859 ( .IN1(\s9/msel/gnt_p2 [0]), .IN2(n32452), .QN(n32367) );
  OA221X1 U35860 ( .IN1(\s9/msel/gnt_p2 [1]), .IN2(n32410), .IN3(n34466), 
        .IN4(n32414), .IN5(\s9/msel/gnt_p2 [0]), .Q(n32454) );
  OR4X1 U35861 ( .IN1(n32368), .IN2(n34152), .IN3(n32367), .IN4(n32454), .Q(
        n32376) );
  OA21X1 U35862 ( .IN1(n32433), .IN2(n32388), .IN3(n34469), .Q(n32450) );
  OA21X1 U35863 ( .IN1(n32444), .IN2(n32391), .IN3(n32450), .Q(n32401) );
  INVX0 U35864 ( .INP(n32369), .ZN(n32415) );
  NAND2X0 U35865 ( .IN1(\s9/msel/gnt_p2 [0]), .IN2(n32415), .QN(n32445) );
  OA21X1 U35866 ( .IN1(\s9/msel/gnt_p2 [0]), .IN2(n32446), .IN3(n32445), .Q(
        n32399) );
  NOR2X0 U35867 ( .IN1(n32399), .IN2(\s9/msel/gnt_p2 [1]), .QN(n32374) );
  INVX0 U35868 ( .INP(n32422), .ZN(n32437) );
  NOR2X0 U35869 ( .IN1(n32410), .IN2(n32437), .QN(n34153) );
  NAND2X0 U35870 ( .IN1(n34154), .IN2(n34153), .QN(n32372) );
  INVX0 U35871 ( .INP(n32380), .ZN(n32383) );
  NAND2X0 U35872 ( .IN1(\s9/msel/gnt_p2 [0]), .IN2(n34466), .QN(n32385) );
  NOR2X0 U35873 ( .IN1(\s9/msel/gnt_p2 [0]), .IN2(\s9/msel/gnt_p2 [1]), .QN(
        n32430) );
  NAND2X0 U35874 ( .IN1(n32430), .IN2(n32369), .QN(n32384) );
  NAND2X0 U35875 ( .IN1(n32385), .IN2(n32384), .QN(n32370) );
  AO22X1 U35876 ( .IN1(\s9/msel/gnt_p2 [1]), .IN2(n32433), .IN3(n32383), .IN4(
        n32370), .Q(n32371) );
  NAND2X0 U35877 ( .IN1(n32372), .IN2(n32371), .QN(n32373) );
  NOR2X0 U35878 ( .IN1(n32374), .IN2(n32373), .QN(n32375) );
  AO22X1 U35879 ( .IN1(\s9/msel/gnt_p2 [2]), .IN2(n32376), .IN3(n32401), .IN4(
        n32375), .Q(n17772) );
  AND2X1 U35880 ( .IN1(n34466), .IN2(n32444), .Q(n32417) );
  OA21X1 U35881 ( .IN1(n32417), .IN2(n32378), .IN3(n34154), .Q(n32387) );
  OA22X1 U35882 ( .IN1(n32387), .IN2(n32377), .IN3(n32383), .IN4(n32378), .Q(
        n32379) );
  INVX0 U35883 ( .INP(n32378), .ZN(n32381) );
  NAND4X0 U35884 ( .IN1(\s9/msel/gnt_p2 [1]), .IN2(n32381), .IN3(n32422), 
        .IN4(n32421), .QN(n32389) );
  NAND2X0 U35885 ( .IN1(n32379), .IN2(n32389), .QN(n32398) );
  AO221X1 U35886 ( .IN1(n32381), .IN2(n34153), .IN3(n32381), .IN4(n32380), 
        .IN5(n32388), .Q(n32397) );
  NAND2X0 U35887 ( .IN1(n32382), .IN2(n34153), .QN(n32390) );
  AND2X1 U35888 ( .IN1(n32390), .IN2(n32383), .Q(n32386) );
  OA221X1 U35889 ( .IN1(n32386), .IN2(n32385), .IN3(n32386), .IN4(n32384), 
        .IN5(n34469), .Q(n32395) );
  OR4X1 U35890 ( .IN1(n32388), .IN2(n32410), .IN3(n32437), .IN4(n32387), .Q(
        n32394) );
  NAND3X0 U35891 ( .IN1(n32390), .IN2(n32389), .IN3(n32433), .QN(n32392) );
  INVX0 U35892 ( .INP(n32391), .ZN(n32403) );
  NAND2X0 U35893 ( .IN1(n32392), .IN2(n32403), .QN(n32393) );
  NAND3X0 U35894 ( .IN1(n32395), .IN2(n32394), .IN3(n32393), .QN(n32396) );
  OA221X1 U35895 ( .IN1(n34469), .IN2(n32398), .IN3(n34469), .IN4(n32397), 
        .IN5(n32396), .Q(n32409) );
  NAND2X0 U35896 ( .IN1(n32409), .IN2(n32399), .QN(n32400) );
  NAND2X0 U35897 ( .IN1(n32401), .IN2(n32400), .QN(n32408) );
  NAND2X0 U35898 ( .IN1(n32437), .IN2(n34462), .QN(n32402) );
  NAND3X0 U35899 ( .IN1(n32402), .IN2(n32421), .IN3(n32409), .QN(n32406) );
  NAND2X0 U35900 ( .IN1(n32414), .IN2(n32428), .QN(n32405) );
  NAND2X0 U35901 ( .IN1(n32435), .IN2(n32403), .QN(n32404) );
  NAND4X0 U35902 ( .IN1(\s9/msel/gnt_p2 [2]), .IN2(n32406), .IN3(n32405), 
        .IN4(n32404), .QN(n32407) );
  AO22X1 U35903 ( .IN1(\s9/msel/gnt_p2 [1]), .IN2(n32409), .IN3(n32408), .IN4(
        n32407), .Q(n17771) );
  NAND2X0 U35904 ( .IN1(n32422), .IN2(n32410), .QN(n32432) );
  NAND2X0 U35905 ( .IN1(n32433), .IN2(n32432), .QN(n32418) );
  AO21X1 U35906 ( .IN1(n32444), .IN2(n32418), .IN3(n32415), .Q(n32427) );
  INVX0 U35907 ( .INP(n32427), .ZN(n32413) );
  NAND4X0 U35908 ( .IN1(n32414), .IN2(n32444), .IN3(n32411), .IN4(n32422), 
        .QN(n32412) );
  NAND2X0 U35909 ( .IN1(n32413), .IN2(n32412), .QN(n32426) );
  INVX0 U35910 ( .INP(n32430), .ZN(n32425) );
  AO21X1 U35911 ( .IN1(n32415), .IN2(n32446), .IN3(n32414), .Q(n32420) );
  NOR2X0 U35912 ( .IN1(n32435), .IN2(n32437), .QN(n32416) );
  OA221X1 U35913 ( .IN1(n32420), .IN2(\s9/msel/gnt_p2 [0]), .IN3(n32420), 
        .IN4(n32446), .IN5(n32416), .Q(n32419) );
  OA22X1 U35914 ( .IN1(n32419), .IN2(n32418), .IN3(n32417), .IN4(n34462), .Q(
        n32424) );
  INVX0 U35915 ( .INP(n32420), .ZN(n32431) );
  NAND2X0 U35916 ( .IN1(n32444), .IN2(n32446), .QN(n32434) );
  OR2X1 U35917 ( .IN1(n34462), .IN2(n32434), .Q(n32436) );
  OAI221X1 U35918 ( .IN1(n32435), .IN2(n32431), .IN3(n32435), .IN4(n32436), 
        .IN5(n32421), .QN(n32429) );
  AND3X1 U35919 ( .IN1(n32429), .IN2(n32422), .IN3(n32428), .Q(n32423) );
  AO221X1 U35920 ( .IN1(n32430), .IN2(n32426), .IN3(n32425), .IN4(n32424), 
        .IN5(n32423), .Q(n32443) );
  NAND3X0 U35921 ( .IN1(n32428), .IN2(n32446), .IN3(n32427), .QN(n32441) );
  NAND2X0 U35922 ( .IN1(n32430), .IN2(n32429), .QN(n32440) );
  OA221X1 U35923 ( .IN1(n32434), .IN2(n32433), .IN3(n32434), .IN4(n32432), 
        .IN5(n32431), .Q(n32438) );
  AO221X1 U35924 ( .IN1(n32438), .IN2(n32437), .IN3(n32438), .IN4(n32436), 
        .IN5(n32435), .Q(n32439) );
  NAND4X0 U35925 ( .IN1(\s9/msel/gnt_p2 [2]), .IN2(n32441), .IN3(n32440), 
        .IN4(n32439), .QN(n32442) );
  OA21X1 U35926 ( .IN1(\s9/msel/gnt_p2 [2]), .IN2(n32443), .IN3(n32442), .Q(
        n32451) );
  NAND3X0 U35927 ( .IN1(\s9/msel/gnt_p2 [1]), .IN2(n32451), .IN3(n32444), .QN(
        n32449) );
  INVX0 U35928 ( .INP(n32445), .ZN(n32447) );
  OAI221X1 U35929 ( .IN1(n32447), .IN2(n32446), .IN3(n32447), .IN4(n32451), 
        .IN5(n34466), .QN(n32448) );
  NAND3X0 U35930 ( .IN1(n32450), .IN2(n32449), .IN3(n32448), .QN(n32455) );
  OA221X1 U35931 ( .IN1(\s9/msel/gnt_p2 [0]), .IN2(\s9/msel/gnt_p2 [2]), .IN3(
        \s9/msel/gnt_p2 [0]), .IN4(n32452), .IN5(n32451), .Q(n32453) );
  AO221X1 U35932 ( .IN1(n32455), .IN2(n34469), .IN3(n32455), .IN4(n32454), 
        .IN5(n32453), .Q(n17770) );
  NOR2X0 U35933 ( .IN1(n32456), .IN2(n34379), .QN(n32457) );
  MUX21X1 U35934 ( .IN1(n34619), .IN2(s15_data_o[0]), .S(n32457), .Q(n17769)
         );
  MUX21X1 U35935 ( .IN1(n34582), .IN2(s15_data_o[1]), .S(n32457), .Q(n17768)
         );
  MUX21X1 U35936 ( .IN1(n34638), .IN2(s15_data_o[2]), .S(n32457), .Q(n17767)
         );
  MUX21X1 U35937 ( .IN1(n34611), .IN2(s15_data_o[3]), .S(n32457), .Q(n17766)
         );
  MUX21X1 U35938 ( .IN1(n34322), .IN2(s15_data_o[4]), .S(n32457), .Q(n17765)
         );
  MUX21X1 U35939 ( .IN1(n34503), .IN2(s15_data_o[5]), .S(n32457), .Q(n17764)
         );
  MUX21X1 U35940 ( .IN1(n34606), .IN2(s15_data_o[6]), .S(n32457), .Q(n17763)
         );
  MUX21X1 U35941 ( .IN1(n34372), .IN2(s15_data_o[7]), .S(n32457), .Q(n17762)
         );
  MUX21X1 U35942 ( .IN1(n34620), .IN2(s15_data_o[8]), .S(n32457), .Q(n17761)
         );
  MUX21X1 U35943 ( .IN1(n34583), .IN2(s15_data_o[9]), .S(n32457), .Q(n17760)
         );
  MUX21X1 U35944 ( .IN1(n34323), .IN2(s15_data_o[10]), .S(n32457), .Q(n17759)
         );
  MUX21X1 U35945 ( .IN1(n34504), .IN2(s15_data_o[11]), .S(n32457), .Q(n17758)
         );
  MUX21X1 U35946 ( .IN1(n34632), .IN2(s15_data_o[12]), .S(n32457), .Q(n17757)
         );
  MUX21X1 U35947 ( .IN1(n34568), .IN2(s15_data_o[13]), .S(n32457), .Q(n17756)
         );
  MUX21X1 U35948 ( .IN1(n34353), .IN2(s15_data_o[14]), .S(n32457), .Q(n17755)
         );
  MUX21X1 U35949 ( .IN1(n34505), .IN2(s15_data_o[15]), .S(n32457), .Q(n17754)
         );
  NOR2X0 U35950 ( .IN1(\s10/msel/gnt_p3 [1]), .IN2(n32509), .QN(n32503) );
  NAND2X0 U35951 ( .IN1(n32511), .IN2(n34251), .QN(n32520) );
  AO221X1 U35952 ( .IN1(n34251), .IN2(n32539), .IN3(\s10/msel/gnt_p3 [1]), 
        .IN4(n32511), .IN5(n34472), .Q(n32546) );
  NAND2X0 U35953 ( .IN1(\s10/msel/gnt_p3 [0]), .IN2(\s10/msel/gnt_p3 [2]), 
        .QN(n32559) );
  NAND2X0 U35954 ( .IN1(n32546), .IN2(n32559), .QN(n32458) );
  NAND4X0 U35955 ( .IN1(n32508), .IN2(n32520), .IN3(n32459), .IN4(n32458), 
        .QN(n32466) );
  NAND2X0 U35956 ( .IN1(\s10/msel/gnt_p3 [1]), .IN2(n34464), .QN(n32483) );
  NAND2X0 U35957 ( .IN1(\s10/msel/gnt_p3 [0]), .IN2(\s10/msel/gnt_p3 [1]), 
        .QN(n32521) );
  MUX21X1 U35958 ( .IN1(n32549), .IN2(n32505), .S(\s10/msel/gnt_p3 [0]), .Q(
        n32497) );
  OAI222X1 U35959 ( .IN1(n32483), .IN2(n32550), .IN3(n32521), .IN4(n32513), 
        .IN5(n32497), .IN6(\s10/msel/gnt_p3 [1]), .QN(n32464) );
  NAND2X0 U35960 ( .IN1(\s10/msel/gnt_p3 [0]), .IN2(n34251), .QN(n32547) );
  OA21X1 U35961 ( .IN1(n32550), .IN2(n32547), .IN3(n32483), .Q(n32535) );
  INVX0 U35962 ( .INP(n32460), .ZN(n32472) );
  OA22X1 U35963 ( .IN1(n32513), .IN2(n32535), .IN3(n32505), .IN4(n32472), .Q(
        n32461) );
  NAND2X0 U35964 ( .IN1(n32461), .IN2(n32521), .QN(n32462) );
  AND3X1 U35965 ( .IN1(n32464), .IN2(n32463), .IN3(n32462), .Q(n32465) );
  OA22X1 U35966 ( .IN1(n32503), .IN2(n32466), .IN3(\s10/msel/gnt_p3 [2]), 
        .IN4(n32465), .Q(n17753) );
  NAND2X0 U35967 ( .IN1(n34464), .IN2(n34251), .QN(n32528) );
  NAND3X0 U35968 ( .IN1(n32528), .IN2(n32521), .IN3(n32472), .QN(n32489) );
  INVX0 U35969 ( .INP(n32489), .ZN(n32468) );
  NOR2X0 U35970 ( .IN1(n32483), .IN2(n32482), .QN(n32467) );
  NOR2X0 U35971 ( .IN1(n32468), .IN2(n32467), .QN(n32470) );
  INVX0 U35972 ( .INP(n32509), .ZN(n32499) );
  NOR2X0 U35973 ( .IN1(n32499), .IN2(n32528), .QN(n32474) );
  NAND2X0 U35974 ( .IN1(n32513), .IN2(n32474), .QN(n32469) );
  NAND2X0 U35975 ( .IN1(n32470), .IN2(n32469), .QN(n32471) );
  OA221X1 U35976 ( .IN1(n32471), .IN2(n32550), .IN3(n32471), .IN4(n32474), 
        .IN5(n32481), .Q(n32493) );
  NOR2X0 U35977 ( .IN1(n32549), .IN2(n32521), .QN(n32507) );
  INVX0 U35978 ( .INP(n32505), .ZN(n32548) );
  AO221X1 U35979 ( .IN1(n32473), .IN2(\s10/msel/gnt_p3 [1]), .IN3(n32473), 
        .IN4(n32511), .IN5(n32472), .Q(n32486) );
  NAND3X0 U35980 ( .IN1(n32507), .IN2(n32548), .IN3(n32486), .QN(n32478) );
  NOR2X0 U35981 ( .IN1(n34251), .IN2(n32508), .QN(n32504) );
  INVX0 U35982 ( .INP(n32504), .ZN(n32477) );
  INVX0 U35983 ( .INP(n32474), .ZN(n32475) );
  AO21X1 U35984 ( .IN1(n32547), .IN2(n32475), .IN3(n32480), .Q(n32476) );
  NAND4X0 U35985 ( .IN1(\s10/msel/gnt_p3 [2]), .IN2(n32478), .IN3(n32477), 
        .IN4(n32476), .QN(n32492) );
  INVX0 U35986 ( .INP(n32528), .ZN(n32487) );
  NOR2X0 U35987 ( .IN1(n32527), .IN2(n32507), .QN(n32479) );
  OA22X1 U35988 ( .IN1(n32487), .IN2(n32480), .IN3(n32505), .IN4(n32479), .Q(
        n32485) );
  INVX0 U35989 ( .INP(n32481), .ZN(n32484) );
  AO221X1 U35990 ( .IN1(n32485), .IN2(n32484), .IN3(n32485), .IN4(n32483), 
        .IN5(n32482), .Q(n32490) );
  NAND3X0 U35991 ( .IN1(n32487), .IN2(n32548), .IN3(n32486), .QN(n32488) );
  NAND4X0 U35992 ( .IN1(n32490), .IN2(n34472), .IN3(n32489), .IN4(n32488), 
        .QN(n32491) );
  OA21X1 U35993 ( .IN1(n32493), .IN2(n32492), .IN3(n32491), .Q(n32496) );
  AO22X1 U35994 ( .IN1(\s10/msel/gnt_p3 [1]), .IN2(n32511), .IN3(n32496), 
        .IN4(n32512), .Q(n32494) );
  NAND3X0 U35995 ( .IN1(\s10/msel/gnt_p3 [2]), .IN2(n34464), .IN3(n32494), 
        .QN(n32502) );
  INVX0 U35996 ( .INP(n32521), .ZN(n32495) );
  NAND2X0 U35997 ( .IN1(n32513), .IN2(n32495), .QN(n32552) );
  INVX0 U35998 ( .INP(n32496), .ZN(n32498) );
  AO221X1 U35999 ( .IN1(n32552), .IN2(n32497), .IN3(n32552), .IN4(n32498), 
        .IN5(\s10/msel/gnt_p3 [2]), .Q(n32501) );
  AO221X1 U36000 ( .IN1(n34251), .IN2(n32499), .IN3(n34251), .IN4(n32559), 
        .IN5(n32498), .Q(n32500) );
  NAND3X0 U36001 ( .IN1(n32502), .IN2(n32501), .IN3(n32500), .QN(n17752) );
  NOR2X0 U36002 ( .IN1(n32504), .IN2(n32503), .QN(n32558) );
  NOR2X0 U36003 ( .IN1(n32511), .IN2(n32539), .QN(n32534) );
  NOR2X0 U36004 ( .IN1(n32509), .IN2(n32539), .QN(n32515) );
  OR2X1 U36005 ( .IN1(n32513), .IN2(n32515), .Q(n32532) );
  AO21X1 U36006 ( .IN1(\s10/msel/gnt_p3 [0]), .IN2(n32534), .IN3(n32532), .Q(
        n32506) );
  AO21X1 U36007 ( .IN1(n32526), .IN2(n32506), .IN3(n32505), .Q(n32525) );
  NAND2X0 U36008 ( .IN1(n32507), .IN2(n32525), .QN(n32524) );
  OA21X1 U36009 ( .IN1(n32549), .IN2(n32548), .IN3(n32508), .Q(n32537) );
  NOR2X0 U36010 ( .IN1(n32550), .IN2(n32549), .QN(n32514) );
  NAND2X0 U36011 ( .IN1(\s10/msel/gnt_p3 [0]), .IN2(n32514), .QN(n32510) );
  OA221X1 U36012 ( .IN1(n32511), .IN2(n32537), .IN3(n32511), .IN4(n32510), 
        .IN5(n32509), .Q(n32540) );
  OR2X1 U36013 ( .IN1(n32528), .IN2(n32540), .Q(n32523) );
  INVX0 U36014 ( .INP(n32549), .ZN(n32531) );
  NAND4X0 U36015 ( .IN1(\s10/msel/gnt_p3 [0]), .IN2(n32531), .IN3(n32526), 
        .IN4(n32512), .QN(n32518) );
  NAND2X0 U36016 ( .IN1(n32514), .IN2(n32513), .QN(n32517) );
  NAND3X0 U36017 ( .IN1(n32515), .IN2(n32531), .IN3(n32526), .QN(n32516) );
  NAND4X0 U36018 ( .IN1(n32537), .IN2(n32518), .IN3(n32517), .IN4(n32516), 
        .QN(n32519) );
  NAND3X0 U36019 ( .IN1(n32521), .IN2(n32520), .IN3(n32519), .QN(n32522) );
  NAND4X0 U36020 ( .IN1(\s10/msel/gnt_p3 [2]), .IN2(n32524), .IN3(n32523), 
        .IN4(n32522), .QN(n32545) );
  INVX0 U36021 ( .INP(n32525), .ZN(n32530) );
  NAND3X0 U36022 ( .IN1(n32527), .IN2(n32534), .IN3(n32526), .QN(n32529) );
  AO21X1 U36023 ( .IN1(n32530), .IN2(n32529), .IN3(n32528), .Q(n32543) );
  AND3X1 U36024 ( .IN1(n32531), .IN2(n32534), .IN3(\s10/msel/gnt_p3 [0]), .Q(
        n32533) );
  NOR2X0 U36025 ( .IN1(n32533), .IN2(n32532), .QN(n32538) );
  INVX0 U36026 ( .INP(n32534), .ZN(n32536) );
  AO221X1 U36027 ( .IN1(n32538), .IN2(n32537), .IN3(n32538), .IN4(n32536), 
        .IN5(n32535), .Q(n32542) );
  OR3X1 U36028 ( .IN1(n34251), .IN2(n32540), .IN3(n32539), .Q(n32541) );
  NAND4X0 U36029 ( .IN1(n34472), .IN2(n32543), .IN3(n32542), .IN4(n32541), 
        .QN(n32544) );
  NAND2X0 U36030 ( .IN1(n32545), .IN2(n32544), .QN(n32557) );
  AND2X1 U36031 ( .IN1(n34464), .IN2(n32546), .Q(n32556) );
  NOR2X0 U36032 ( .IN1(n32548), .IN2(n32547), .QN(n32554) );
  AO221X1 U36033 ( .IN1(\s10/msel/gnt_p3 [1]), .IN2(n32550), .IN3(n34251), 
        .IN4(n32549), .IN5(n32557), .Q(n32551) );
  NAND2X0 U36034 ( .IN1(n32552), .IN2(n32551), .QN(n32553) );
  NOR2X0 U36035 ( .IN1(n32554), .IN2(n32553), .QN(n32555) );
  OAI222X1 U36036 ( .IN1(n32559), .IN2(n32558), .IN3(n32557), .IN4(n32556), 
        .IN5(n32555), .IN6(\s10/msel/gnt_p3 [2]), .QN(n17751) );
  INVX0 U36037 ( .INP(n32560), .ZN(n32562) );
  NAND2X0 U36038 ( .IN1(n34253), .IN2(n32582), .QN(n32561) );
  NAND4X0 U36039 ( .IN1(\s10/msel/gnt_p1 [2]), .IN2(n32563), .IN3(n32562), 
        .IN4(n32561), .QN(n32575) );
  NOR2X0 U36040 ( .IN1(n32564), .IN2(n32580), .QN(n32572) );
  OA21X1 U36041 ( .IN1(\s10/msel/gnt_p1 [0]), .IN2(n32566), .IN3(n32565), .Q(
        n32601) );
  NOR2X0 U36042 ( .IN1(\s10/msel/gnt_p1 [1]), .IN2(n32601), .QN(n32571) );
  NAND3X0 U36043 ( .IN1(n34434), .IN2(n32567), .IN3(\s10/msel/gnt_p1 [1]), 
        .QN(n32569) );
  NAND2X0 U36044 ( .IN1(n32569), .IN2(n32568), .QN(n32599) );
  NOR4X0 U36045 ( .IN1(n32572), .IN2(n32571), .IN3(n32570), .IN4(n32599), .QN(
        n32573) );
  AO222X1 U36046 ( .IN1(\s10/msel/gnt_p1 [2]), .IN2(n32575), .IN3(
        \s10/msel/gnt_p1 [2]), .IN4(n32574), .IN5(n32575), .IN6(n32573), .Q(
        n17750) );
  NOR2X0 U36047 ( .IN1(\s10/msel/gnt_p1 [0]), .IN2(n34253), .QN(n32597) );
  NAND4X0 U36048 ( .IN1(n32578), .IN2(n32577), .IN3(n32586), .IN4(n32576), 
        .QN(n32588) );
  NAND2X0 U36049 ( .IN1(n32580), .IN2(n32579), .QN(n32590) );
  NAND3X0 U36050 ( .IN1(n34253), .IN2(n32588), .IN3(n32590), .QN(n32585) );
  OA21X1 U36051 ( .IN1(n32589), .IN2(n32582), .IN3(n32581), .Q(n32587) );
  NAND3X0 U36052 ( .IN1(\s10/msel/gnt_p1 [1]), .IN2(n32587), .IN3(n32583), 
        .QN(n32584) );
  NAND3X0 U36053 ( .IN1(n32586), .IN2(n32585), .IN3(n32584), .QN(n32600) );
  AND2X1 U36054 ( .IN1(n32588), .IN2(n32587), .Q(n32593) );
  AND2X1 U36055 ( .IN1(n32590), .IN2(n32589), .Q(n32592) );
  OA22X1 U36056 ( .IN1(\s10/msel/gnt_p1 [1]), .IN2(n32593), .IN3(n32592), 
        .IN4(n32591), .Q(n32594) );
  MUX21X1 U36057 ( .IN1(n32600), .IN2(n32594), .S(\s10/msel/gnt_p1 [2]), .Q(
        n32602) );
  NAND2X0 U36058 ( .IN1(n32595), .IN2(n34434), .QN(n32596) );
  AO22X1 U36059 ( .IN1(n32598), .IN2(n32597), .IN3(n32602), .IN4(n32596), .Q(
        n32605) );
  AO21X1 U36060 ( .IN1(n32601), .IN2(n32600), .IN3(n32599), .Q(n32604) );
  AND2X1 U36061 ( .IN1(\s10/msel/gnt_p1 [1]), .IN2(n32602), .Q(n32603) );
  AO221X1 U36062 ( .IN1(\s10/msel/gnt_p1 [2]), .IN2(n32605), .IN3(n34610), 
        .IN4(n32604), .IN5(n32603), .Q(n17749) );
  NAND3X0 U36063 ( .IN1(n13645), .IN2(n13619), .IN3(m5s10_cyc), .QN(n32650) );
  INVX0 U36064 ( .INP(n32650), .ZN(n32643) );
  NAND3X0 U36065 ( .IN1(n13541), .IN2(n13494), .IN3(m7s10_cyc), .QN(n32668) );
  INVX0 U36066 ( .INP(n32668), .ZN(n32606) );
  OA221X1 U36067 ( .IN1(\s10/msel/gnt_p0 [1]), .IN2(n32643), .IN3(n34257), 
        .IN4(n32606), .IN5(\s10/msel/gnt_p0 [0]), .Q(n32694) );
  NOR2X0 U36068 ( .IN1(\s10/msel/gnt_p0 [1]), .IN2(n34417), .QN(n32642) );
  NAND3X0 U36069 ( .IN1(n13593), .IN2(n13567), .IN3(m6s10_cyc), .QN(n32648) );
  NAND2X0 U36070 ( .IN1(n32642), .IN2(n32648), .QN(n32661) );
  AO21X1 U36071 ( .IN1(n34257), .IN2(n32661), .IN3(n32606), .Q(n32619) );
  NAND2X0 U36072 ( .IN1(n32648), .IN2(n32668), .QN(n32620) );
  NAND3X0 U36073 ( .IN1(n13697), .IN2(n13671), .IN3(m4s10_cyc), .QN(n32655) );
  MUX21X1 U36074 ( .IN1(n32655), .IN2(n32648), .S(\s10/msel/gnt_p0 [1]), .Q(
        n32692) );
  NOR2X0 U36075 ( .IN1(\s10/msel/gnt_p0 [0]), .IN2(n32692), .QN(n32607) );
  AO221X1 U36076 ( .IN1(n32619), .IN2(n32643), .IN3(n32619), .IN4(n32620), 
        .IN5(n32607), .Q(n32608) );
  NOR2X0 U36077 ( .IN1(n32694), .IN2(n32608), .QN(n32610) );
  NAND3X0 U36078 ( .IN1(n13920), .IN2(n13879), .IN3(m0s10_cyc), .QN(n32647) );
  INVX0 U36079 ( .INP(n32647), .ZN(n32685) );
  NAND3X0 U36080 ( .IN1(n13853), .IN2(n13827), .IN3(m1s10_cyc), .QN(n32649) );
  INVX0 U36081 ( .INP(n32649), .ZN(n32644) );
  NOR2X0 U36082 ( .IN1(n32685), .IN2(n32644), .QN(n32621) );
  NAND3X0 U36083 ( .IN1(n13801), .IN2(n13775), .IN3(m2s10_cyc), .QN(n32646) );
  INVX0 U36084 ( .INP(n32646), .ZN(n32686) );
  NAND3X0 U36085 ( .IN1(n13749), .IN2(n13723), .IN3(m3s10_cyc), .QN(n32656) );
  INVX0 U36086 ( .INP(n32656), .ZN(n32652) );
  NOR2X0 U36087 ( .IN1(n32686), .IN2(n32652), .QN(n32618) );
  NAND2X0 U36088 ( .IN1(n32621), .IN2(n32618), .QN(n32609) );
  NAND2X0 U36089 ( .IN1(n32610), .IN2(n32609), .QN(n32616) );
  NAND2X0 U36090 ( .IN1(\s10/msel/gnt_p0 [1]), .IN2(n34417), .QN(n32662) );
  NAND2X0 U36091 ( .IN1(\s10/msel/gnt_p0 [0]), .IN2(\s10/msel/gnt_p0 [1]), 
        .QN(n32612) );
  OA21X1 U36092 ( .IN1(n32656), .IN2(n32612), .IN3(n34451), .Q(n32687) );
  OA21X1 U36093 ( .IN1(n32646), .IN2(n32662), .IN3(n32687), .Q(n32634) );
  NAND2X0 U36094 ( .IN1(n32650), .IN2(n32655), .QN(n32617) );
  INVX0 U36095 ( .INP(n32642), .ZN(n32625) );
  OA21X1 U36096 ( .IN1(n32686), .IN2(n32625), .IN3(n32662), .Q(n32677) );
  NAND2X0 U36097 ( .IN1(n34417), .IN2(n34257), .QN(n32669) );
  OR2X1 U36098 ( .IN1(n32669), .IN2(n32644), .Q(n32626) );
  INVX0 U36099 ( .INP(n32618), .ZN(n32611) );
  OA22X1 U36100 ( .IN1(n32652), .IN2(n32677), .IN3(n32626), .IN4(n32611), .Q(
        n32613) );
  MUX21X1 U36101 ( .IN1(n32685), .IN2(n32644), .S(\s10/msel/gnt_p0 [0]), .Q(
        n32635) );
  AOI22X1 U36102 ( .IN1(n32613), .IN2(n32612), .IN3(n34257), .IN4(n32635), 
        .QN(n32614) );
  OA21X1 U36103 ( .IN1(n32620), .IN2(n32617), .IN3(n32614), .Q(n32615) );
  AO22X1 U36104 ( .IN1(\s10/msel/gnt_p0 [2]), .IN2(n32616), .IN3(n32634), 
        .IN4(n32615), .Q(n17747) );
  NAND2X0 U36105 ( .IN1(n32618), .IN2(n32617), .QN(n32628) );
  OR4X1 U36106 ( .IN1(n32620), .IN2(\s10/msel/gnt_p0 [1]), .IN3(n32686), .IN4(
        n32652), .Q(n32627) );
  OA221X1 U36107 ( .IN1(n32619), .IN2(n32621), .IN3(n32619), .IN4(n32628), 
        .IN5(n32627), .Q(n32623) );
  NOR2X0 U36108 ( .IN1(n32621), .IN2(n32620), .QN(n32624) );
  NOR2X0 U36109 ( .IN1(n32643), .IN2(n32624), .QN(n32622) );
  AO221X1 U36110 ( .IN1(n32623), .IN2(n32622), .IN3(n32623), .IN4(n32669), 
        .IN5(n34451), .Q(n32636) );
  INVX0 U36111 ( .INP(n32655), .ZN(n32672) );
  OR4X1 U36112 ( .IN1(n34257), .IN2(n32672), .IN3(n32643), .IN4(n32624), .Q(
        n32632) );
  OR2X1 U36113 ( .IN1(n32656), .IN2(n32662), .Q(n32631) );
  NAND2X0 U36114 ( .IN1(n32626), .IN2(n32625), .QN(n32629) );
  NAND3X0 U36115 ( .IN1(n32629), .IN2(n32628), .IN3(n32627), .QN(n32630) );
  NAND4X0 U36116 ( .IN1(n34451), .IN2(n32632), .IN3(n32631), .IN4(n32630), 
        .QN(n32633) );
  NAND2X0 U36117 ( .IN1(n32636), .IN2(n32633), .QN(n32639) );
  OA21X1 U36118 ( .IN1(n32639), .IN2(n32635), .IN3(n32634), .Q(n32641) );
  INVX0 U36119 ( .INP(n32636), .ZN(n32638) );
  OA221X1 U36120 ( .IN1(\s10/msel/gnt_p0 [0]), .IN2(n32672), .IN3(n34417), 
        .IN4(n32643), .IN5(\s10/msel/gnt_p0 [2]), .Q(n32637) );
  OA22X1 U36121 ( .IN1(n32638), .IN2(n32637), .IN3(n32648), .IN4(n32662), .Q(
        n32640) );
  OAI22X1 U36122 ( .IN1(n32641), .IN2(n32640), .IN3(n34257), .IN4(n32639), 
        .QN(n17746) );
  NAND2X0 U36123 ( .IN1(n32644), .IN2(n32642), .QN(n32689) );
  NAND2X0 U36124 ( .IN1(n32648), .IN2(n32655), .QN(n32675) );
  NOR2X0 U36125 ( .IN1(n34417), .IN2(n32675), .QN(n32645) );
  NAND2X0 U36126 ( .IN1(n32643), .IN2(n32655), .QN(n32657) );
  NAND2X0 U36127 ( .IN1(n32656), .IN2(n32657), .QN(n32674) );
  AO221X1 U36128 ( .IN1(n32646), .IN2(n32645), .IN3(n32646), .IN4(n32674), 
        .IN5(n32644), .Q(n32667) );
  NAND3X0 U36129 ( .IN1(\s10/msel/gnt_p0 [1]), .IN2(n32667), .IN3(n32647), 
        .QN(n32666) );
  INVX0 U36130 ( .INP(n32648), .ZN(n32654) );
  OA21X1 U36131 ( .IN1(n32685), .IN2(n32649), .IN3(n32668), .Q(n32676) );
  NOR2X0 U36132 ( .IN1(n32686), .IN2(n32685), .QN(n32659) );
  NAND2X0 U36133 ( .IN1(\s10/msel/gnt_p0 [0]), .IN2(n32659), .QN(n32651) );
  OA221X1 U36134 ( .IN1(n32654), .IN2(n32676), .IN3(n32654), .IN4(n32651), 
        .IN5(n32650), .Q(n32673) );
  NAND2X0 U36135 ( .IN1(n32659), .IN2(n32652), .QN(n32653) );
  AO221X1 U36136 ( .IN1(n32673), .IN2(n32654), .IN3(n32673), .IN4(n32653), 
        .IN5(n32669), .Q(n32665) );
  NAND2X0 U36137 ( .IN1(\s10/msel/gnt_p0 [0]), .IN2(n32655), .QN(n32658) );
  NAND3X0 U36138 ( .IN1(n32658), .IN2(n32657), .IN3(n32656), .QN(n32660) );
  NAND2X0 U36139 ( .IN1(n32660), .IN2(n32659), .QN(n32663) );
  AO22X1 U36140 ( .IN1(n32676), .IN2(n32663), .IN3(n32662), .IN4(n32661), .Q(
        n32664) );
  NAND4X0 U36141 ( .IN1(\s10/msel/gnt_p0 [2]), .IN2(n32666), .IN3(n32665), 
        .IN4(n32664), .QN(n32684) );
  INVX0 U36142 ( .INP(n32667), .ZN(n32671) );
  OR3X1 U36143 ( .IN1(n32668), .IN2(n32675), .IN3(n32686), .Q(n32670) );
  AO21X1 U36144 ( .IN1(n32671), .IN2(n32670), .IN3(n32669), .Q(n32682) );
  OR3X1 U36145 ( .IN1(n34257), .IN2(n32673), .IN3(n32672), .Q(n32681) );
  INVX0 U36146 ( .INP(n32674), .ZN(n32679) );
  AO221X1 U36147 ( .IN1(n32676), .IN2(n32685), .IN3(n32676), .IN4(n34417), 
        .IN5(n32675), .Q(n32678) );
  AO21X1 U36148 ( .IN1(n32679), .IN2(n32678), .IN3(n32677), .Q(n32680) );
  NAND4X0 U36149 ( .IN1(n34451), .IN2(n32682), .IN3(n32681), .IN4(n32680), 
        .QN(n32683) );
  NAND2X0 U36150 ( .IN1(n32684), .IN2(n32683), .QN(n32690) );
  AO221X1 U36151 ( .IN1(\s10/msel/gnt_p0 [1]), .IN2(n32686), .IN3(n34257), 
        .IN4(n32685), .IN5(n32690), .Q(n32688) );
  NAND3X0 U36152 ( .IN1(n32689), .IN2(n32688), .IN3(n32687), .QN(n32695) );
  INVX0 U36153 ( .INP(n32690), .ZN(n32691) );
  OA221X1 U36154 ( .IN1(\s10/msel/gnt_p0 [0]), .IN2(\s10/msel/gnt_p0 [2]), 
        .IN3(\s10/msel/gnt_p0 [0]), .IN4(n32692), .IN5(n32691), .Q(n32693) );
  AO221X1 U36155 ( .IN1(n32695), .IN2(n34451), .IN3(n32695), .IN4(n32694), 
        .IN5(n32693), .Q(n17745) );
  NOR2X0 U36156 ( .IN1(n32696), .IN2(n34255), .QN(n32703) );
  OA221X1 U36157 ( .IN1(\s10/msel/gnt_p2 [0]), .IN2(n32699), .IN3(
        \s10/msel/gnt_p2 [0]), .IN4(n32698), .IN5(n32697), .Q(n32700) );
  OA221X1 U36158 ( .IN1(n32703), .IN2(n32702), .IN3(n32703), .IN4(n32701), 
        .IN5(n32700), .Q(n32713) );
  OA22X1 U36159 ( .IN1(n32706), .IN2(n34255), .IN3(n32705), .IN4(n32704), .Q(
        n32712) );
  NAND2X0 U36160 ( .IN1(n32707), .IN2(n34255), .QN(n32710) );
  NAND3X0 U36161 ( .IN1(n32710), .IN2(n32709), .IN3(n32708), .QN(n32711) );
  OAI22X1 U36162 ( .IN1(n32713), .IN2(n34405), .IN3(n32712), .IN4(n32711), 
        .QN(n17744) );
  NOR2X0 U36163 ( .IN1(n32714), .IN2(n34379), .QN(n32715) );
  MUX21X1 U36164 ( .IN1(n34621), .IN2(s15_data_o[0]), .S(n32715), .Q(n17741)
         );
  MUX21X1 U36165 ( .IN1(n34584), .IN2(s15_data_o[1]), .S(n32715), .Q(n17740)
         );
  MUX21X1 U36166 ( .IN1(n34326), .IN2(s15_data_o[2]), .S(n32715), .Q(n17739)
         );
  MUX21X1 U36167 ( .IN1(n34537), .IN2(s15_data_o[3]), .S(n32715), .Q(n17738)
         );
  MUX21X1 U36168 ( .IN1(n34325), .IN2(s15_data_o[4]), .S(n32715), .Q(n17737)
         );
  MUX21X1 U36169 ( .IN1(n34538), .IN2(s15_data_o[5]), .S(n32715), .Q(n17736)
         );
  MUX21X1 U36170 ( .IN1(n34365), .IN2(s15_data_o[6]), .S(n32715), .Q(n17735)
         );
  MUX21X1 U36171 ( .IN1(n34601), .IN2(s15_data_o[7]), .S(n32715), .Q(n17734)
         );
  MUX21X1 U36172 ( .IN1(n34622), .IN2(s15_data_o[8]), .S(n32715), .Q(n17733)
         );
  MUX21X1 U36173 ( .IN1(n34569), .IN2(s15_data_o[9]), .S(n32715), .Q(n17732)
         );
  MUX21X1 U36174 ( .IN1(n34375), .IN2(s15_data_o[10]), .S(n32715), .Q(n17731)
         );
  MUX21X1 U36175 ( .IN1(n34585), .IN2(s15_data_o[11]), .S(n32715), .Q(n17730)
         );
  MUX21X1 U36176 ( .IN1(n34633), .IN2(s15_data_o[12]), .S(n32715), .Q(n17729)
         );
  MUX21X1 U36177 ( .IN1(n34570), .IN2(s15_data_o[13]), .S(n32715), .Q(n17728)
         );
  MUX21X1 U36178 ( .IN1(n34324), .IN2(s15_data_o[14]), .S(n32715), .Q(n17727)
         );
  MUX21X1 U36179 ( .IN1(n34539), .IN2(s15_data_o[15]), .S(n32715), .Q(n17726)
         );
  NOR2X0 U36180 ( .IN1(n32717), .IN2(n32716), .QN(n34168) );
  INVX0 U36181 ( .INP(n34168), .ZN(n32720) );
  NAND2X0 U36182 ( .IN1(n32778), .IN2(n34419), .QN(n32719) );
  MUX21X1 U36183 ( .IN1(n32736), .IN2(n32749), .S(\s11/msel/gnt_p3 [1]), .Q(
        n32776) );
  NAND2X0 U36184 ( .IN1(n34399), .IN2(n32776), .QN(n32718) );
  NAND4X0 U36185 ( .IN1(n32721), .IN2(n32720), .IN3(n32719), .IN4(n32718), 
        .QN(n32728) );
  AND2X1 U36186 ( .IN1(n32723), .IN2(n32722), .Q(n34169) );
  NOR2X0 U36187 ( .IN1(n34169), .IN2(n32724), .QN(n32727) );
  AO22X1 U36188 ( .IN1(n34419), .IN2(n32725), .IN3(n32739), .IN4(
        \s11/msel/gnt_p3 [1]), .Q(n32726) );
  AO22X1 U36189 ( .IN1(\s11/msel/gnt_p3 [2]), .IN2(n32728), .IN3(n32727), 
        .IN4(n32726), .Q(n17725) );
  INVX0 U36190 ( .INP(n32746), .ZN(n32775) );
  OA21X1 U36191 ( .IN1(n32749), .IN2(n32760), .IN3(n32741), .Q(n32731) );
  NAND3X0 U36192 ( .IN1(n32775), .IN2(n32730), .IN3(n32772), .QN(n32729) );
  NAND2X0 U36193 ( .IN1(n32731), .IN2(n32729), .QN(n32751) );
  NAND3X0 U36194 ( .IN1(\s11/msel/gnt_p3 [1]), .IN2(n32751), .IN3(n32756), 
        .QN(n32738) );
  NAND2X0 U36195 ( .IN1(\s11/msel/gnt_p3 [0]), .IN2(n32730), .QN(n32732) );
  OA21X1 U36196 ( .IN1(n32733), .IN2(n32732), .IN3(n32731), .Q(n32735) );
  INVX0 U36197 ( .INP(n32771), .ZN(n32734) );
  AO221X1 U36198 ( .IN1(n32739), .IN2(n32736), .IN3(n32739), .IN4(n32735), 
        .IN5(n32734), .Q(n32737) );
  NAND3X0 U36199 ( .IN1(n34444), .IN2(n32738), .IN3(n32737), .QN(n32770) );
  NOR2X0 U36200 ( .IN1(\s11/msel/gnt_p3 [0]), .IN2(\s11/msel/gnt_p3 [1]), .QN(
        n32769) );
  INVX0 U36201 ( .INP(n32739), .ZN(n32750) );
  NAND2X0 U36202 ( .IN1(n32750), .IN2(n32771), .QN(n32745) );
  NAND2X0 U36203 ( .IN1(n32756), .IN2(n32771), .QN(n32740) );
  NOR2X0 U36204 ( .IN1(n34399), .IN2(n32740), .QN(n32743) );
  NAND2X0 U36205 ( .IN1(n32741), .IN2(n32749), .QN(n32742) );
  NAND2X0 U36206 ( .IN1(n32743), .IN2(n32742), .QN(n32744) );
  NAND3X0 U36207 ( .IN1(n32746), .IN2(n32745), .IN3(n32744), .QN(n32768) );
  NAND2X0 U36208 ( .IN1(n32747), .IN2(n32768), .QN(n32766) );
  INVX0 U36209 ( .INP(n32769), .ZN(n32748) );
  NOR2X0 U36210 ( .IN1(n32749), .IN2(n32748), .QN(n32754) );
  NAND3X0 U36211 ( .IN1(n32750), .IN2(n32772), .IN3(n32771), .QN(n32758) );
  INVX0 U36212 ( .INP(n32751), .ZN(n32752) );
  NAND2X0 U36213 ( .IN1(n32758), .IN2(n32752), .QN(n32753) );
  NAND2X0 U36214 ( .IN1(n32754), .IN2(n32753), .QN(n32765) );
  NAND2X0 U36215 ( .IN1(n32775), .IN2(n32772), .QN(n32759) );
  NAND4X0 U36216 ( .IN1(n32756), .IN2(n32772), .IN3(n32771), .IN4(n32755), 
        .QN(n32757) );
  AND4X1 U36217 ( .IN1(n32760), .IN2(n32759), .IN3(n32758), .IN4(n32757), .Q(
        n32761) );
  OR3X1 U36218 ( .IN1(n32763), .IN2(n32762), .IN3(n32761), .Q(n32764) );
  NAND4X0 U36219 ( .IN1(\s11/msel/gnt_p3 [2]), .IN2(n32766), .IN3(n32765), 
        .IN4(n32764), .QN(n32767) );
  OA221X1 U36220 ( .IN1(n32770), .IN2(n32769), .IN3(n32770), .IN4(n32768), 
        .IN5(n32767), .Q(n32780) );
  MUX21X1 U36221 ( .IN1(n32772), .IN2(n32771), .S(\s11/msel/gnt_p3 [1]), .Q(
        n32773) );
  AO22X1 U36222 ( .IN1(n32775), .IN2(n32774), .IN3(n32780), .IN4(n32773), .Q(
        n32783) );
  NOR2X0 U36223 ( .IN1(n34444), .IN2(n32776), .QN(n32781) );
  OA221X1 U36224 ( .IN1(\s11/msel/gnt_p3 [1]), .IN2(n32778), .IN3(n34419), 
        .IN4(n32777), .IN5(\s11/msel/gnt_p3 [2]), .Q(n32779) );
  OA22X1 U36225 ( .IN1(\s11/msel/gnt_p3 [0]), .IN2(n32781), .IN3(n32780), 
        .IN4(n32779), .Q(n32782) );
  AO221X1 U36226 ( .IN1(n34444), .IN2(n32784), .IN3(n34444), .IN4(n32783), 
        .IN5(n32782), .Q(n17723) );
  NOR2X0 U36227 ( .IN1(n32786), .IN2(n32785), .QN(n32818) );
  NOR2X0 U36228 ( .IN1(n32787), .IN2(n32818), .QN(n32827) );
  NAND2X0 U36229 ( .IN1(n32789), .IN2(n32788), .QN(n32810) );
  OR2X1 U36230 ( .IN1(\s11/msel/gnt_p1 [1]), .IN2(n32810), .Q(n32822) );
  NOR2X0 U36231 ( .IN1(n32801), .IN2(n32796), .QN(n34174) );
  NOR2X0 U36232 ( .IN1(n32791), .IN2(n32790), .QN(n34175) );
  AO22X1 U36233 ( .IN1(n34174), .IN2(n34175), .IN3(n34655), .IN4(n32792), .Q(
        n32793) );
  AO221X1 U36234 ( .IN1(n32827), .IN2(n32835), .IN3(n32827), .IN4(n32822), 
        .IN5(n32793), .Q(n32794) );
  NAND2X0 U36235 ( .IN1(\s11/msel/gnt_p1 [2]), .IN2(n32794), .QN(n32808) );
  AND2X1 U36236 ( .IN1(n34390), .IN2(n32798), .Q(n32815) );
  NAND2X0 U36237 ( .IN1(n34174), .IN2(n32815), .QN(n32795) );
  OA21X1 U36238 ( .IN1(n32796), .IN2(n34390), .IN3(n32795), .Q(n32805) );
  NAND2X0 U36239 ( .IN1(n32836), .IN2(n32797), .QN(n32809) );
  NOR2X0 U36240 ( .IN1(n32809), .IN2(n32810), .QN(n34173) );
  MUX21X1 U36241 ( .IN1(n32799), .IN2(n32798), .S(\s11/msel/gnt_p1 [0]), .Q(
        n32831) );
  NOR2X0 U36242 ( .IN1(\s11/msel/gnt_p1 [1]), .IN2(n32831), .QN(n32804) );
  NOR2X0 U36243 ( .IN1(\s11/msel/gnt_p1 [2]), .IN2(n32800), .QN(n32803) );
  NAND2X0 U36244 ( .IN1(n32801), .IN2(n32833), .QN(n32802) );
  NAND2X0 U36245 ( .IN1(n32803), .IN2(n32802), .QN(n32830) );
  OR4X1 U36246 ( .IN1(n32805), .IN2(n34173), .IN3(n32804), .IN4(n32830), .Q(
        n32806) );
  NAND3X0 U36247 ( .IN1(n32808), .IN2(n32807), .IN3(n32806), .QN(n17722) );
  INVX0 U36248 ( .INP(n32809), .ZN(n32820) );
  NAND2X0 U36249 ( .IN1(n32822), .IN2(n32820), .QN(n32812) );
  NOR2X0 U36250 ( .IN1(n32810), .IN2(n34175), .QN(n32813) );
  OAI21X1 U36251 ( .IN1(n32812), .IN2(n32813), .IN3(n32811), .QN(n32817) );
  NAND2X0 U36252 ( .IN1(n34174), .IN2(n32812), .QN(n32816) );
  NOR2X0 U36253 ( .IN1(n32835), .IN2(n32813), .QN(n32821) );
  AO222X1 U36254 ( .IN1(n32817), .IN2(n32833), .IN3(n32816), .IN4(n32815), 
        .IN5(n32814), .IN6(n32821), .Q(n32829) );
  INVX0 U36255 ( .INP(n34174), .ZN(n32823) );
  INVX0 U36256 ( .INP(n32818), .ZN(n32819) );
  OA221X1 U36257 ( .IN1(n32823), .IN2(n32820), .IN3(n32823), .IN4(n32819), 
        .IN5(n34175), .Q(n32826) );
  OA21X1 U36258 ( .IN1(n32823), .IN2(n32822), .IN3(n32821), .Q(n32825) );
  OA22X1 U36259 ( .IN1(n32827), .IN2(n32826), .IN3(n32825), .IN4(n32824), .Q(
        n32828) );
  MUX21X1 U36260 ( .IN1(n32829), .IN2(n32828), .S(\s11/msel/gnt_p1 [2]), .Q(
        n32844) );
  AO21X1 U36261 ( .IN1(n32831), .IN2(n32844), .IN3(n32830), .Q(n32843) );
  NAND2X0 U36262 ( .IN1(n32833), .IN2(n32832), .QN(n32841) );
  INVX0 U36263 ( .INP(n32844), .ZN(n32834) );
  NOR2X0 U36264 ( .IN1(n32835), .IN2(n32834), .QN(n32839) );
  INVX0 U36265 ( .INP(n32836), .ZN(n32837) );
  NAND2X0 U36266 ( .IN1(n32837), .IN2(n34655), .QN(n32838) );
  NAND2X0 U36267 ( .IN1(n32839), .IN2(n32838), .QN(n32840) );
  NAND3X0 U36268 ( .IN1(n32841), .IN2(n32840), .IN3(\s11/msel/gnt_p1 [2]), 
        .QN(n32842) );
  AO22X1 U36269 ( .IN1(\s11/msel/gnt_p1 [1]), .IN2(n32844), .IN3(n32843), 
        .IN4(n32842), .Q(n17721) );
  NAND3X0 U36270 ( .IN1(n13802), .IN2(n13776), .IN3(m2s11_cyc), .QN(n32848) );
  NAND2X0 U36271 ( .IN1(\s11/msel/gnt_p0 [1]), .IN2(n34249), .QN(n32888) );
  NAND3X0 U36272 ( .IN1(n13750), .IN2(n13724), .IN3(m3s11_cyc), .QN(n32881) );
  OA22X1 U36273 ( .IN1(n32848), .IN2(n32888), .IN3(n32881), .IN4(n34668), .Q(
        n32845) );
  NAND2X0 U36274 ( .IN1(n32845), .IN2(n34452), .QN(n32868) );
  NAND3X0 U36275 ( .IN1(n13698), .IN2(n13672), .IN3(m4s11_cyc), .QN(n32880) );
  NAND3X0 U36276 ( .IN1(n13646), .IN2(n13620), .IN3(m5s11_cyc), .QN(n32882) );
  AND2X1 U36277 ( .IN1(n32880), .IN2(n32882), .Q(n32860) );
  NAND3X0 U36278 ( .IN1(n13594), .IN2(n13568), .IN3(m6s11_cyc), .QN(n32900) );
  NAND3X0 U36279 ( .IN1(n13542), .IN2(n13495), .IN3(m7s11_cyc), .QN(n32907) );
  NAND2X0 U36280 ( .IN1(n32900), .IN2(n32907), .QN(n32862) );
  INVX0 U36281 ( .INP(n32862), .ZN(n32846) );
  NAND2X0 U36282 ( .IN1(n32848), .IN2(n32881), .QN(n32857) );
  AO22X1 U36283 ( .IN1(n32860), .IN2(n32846), .IN3(n34668), .IN4(n32857), .Q(
        n32847) );
  NOR2X0 U36284 ( .IN1(n32868), .IN2(n32847), .QN(n32854) );
  NAND3X0 U36285 ( .IN1(n13922), .IN2(n13880), .IN3(m0s11_cyc), .QN(n32884) );
  NAND3X0 U36286 ( .IN1(n13854), .IN2(n13828), .IN3(m1s11_cyc), .QN(n32883) );
  OA21X1 U36287 ( .IN1(\s11/msel/gnt_p0 [0]), .IN2(n32884), .IN3(n32883), .Q(
        n32869) );
  INVX0 U36288 ( .INP(n32884), .ZN(n32897) );
  INVX0 U36289 ( .INP(n32848), .ZN(n32906) );
  NOR2X0 U36290 ( .IN1(n32897), .IN2(n32906), .QN(n32885) );
  NAND4X0 U36291 ( .IN1(\s11/msel/gnt_p0 [2]), .IN2(n32885), .IN3(n32881), 
        .IN4(n32883), .QN(n32852) );
  INVX0 U36292 ( .INP(n32880), .ZN(n32911) );
  INVX0 U36293 ( .INP(n32900), .ZN(n32877) );
  MUX21X1 U36294 ( .IN1(n32911), .IN2(n32877), .S(\s11/msel/gnt_p0 [1]), .Q(
        n32922) );
  NAND3X0 U36295 ( .IN1(\s11/msel/gnt_p0 [2]), .IN2(n32922), .IN3(n34249), 
        .QN(n32851) );
  NAND2X0 U36296 ( .IN1(n34668), .IN2(n32882), .QN(n32919) );
  OR2X1 U36297 ( .IN1(n32919), .IN2(n32862), .Q(n32849) );
  NAND2X0 U36298 ( .IN1(\s11/msel/gnt_p0 [1]), .IN2(n32907), .QN(n32920) );
  NAND3X0 U36299 ( .IN1(\s11/msel/gnt_p0 [2]), .IN2(n32849), .IN3(n32920), 
        .QN(n32850) );
  NAND3X0 U36300 ( .IN1(n32852), .IN2(n32851), .IN3(n32850), .QN(n32853) );
  AO221X1 U36301 ( .IN1(n32854), .IN2(\s11/msel/gnt_p0 [1]), .IN3(n32854), 
        .IN4(n32869), .IN5(n32853), .Q(n17719) );
  AND2X1 U36302 ( .IN1(n32884), .IN2(n32883), .Q(n32861) );
  OA21X1 U36303 ( .IN1(n32861), .IN2(n32862), .IN3(n32860), .Q(n32856) );
  AO21X1 U36304 ( .IN1(n32860), .IN2(n32862), .IN3(n32857), .Q(n32855) );
  INVX0 U36305 ( .INP(n32881), .ZN(n32878) );
  AO221X1 U36306 ( .IN1(\s11/msel/gnt_p0 [1]), .IN2(n32856), .IN3(n34668), 
        .IN4(n32855), .IN5(n32878), .Q(n32867) );
  AND2X1 U36307 ( .IN1(n32857), .IN2(n32861), .Q(n32865) );
  NAND3X0 U36308 ( .IN1(\s11/msel/gnt_p0 [0]), .IN2(n34668), .IN3(n32900), 
        .QN(n32887) );
  INVX0 U36309 ( .INP(n32887), .ZN(n32858) );
  NAND2X0 U36310 ( .IN1(n32858), .IN2(n32907), .QN(n32859) );
  OA221X1 U36311 ( .IN1(n32920), .IN2(n32861), .IN3(n32920), .IN4(n32860), 
        .IN5(n32859), .Q(n32864) );
  OA21X1 U36312 ( .IN1(n32865), .IN2(n32862), .IN3(n32882), .Q(n32863) );
  NAND2X0 U36313 ( .IN1(n34249), .IN2(n34668), .QN(n32893) );
  OA22X1 U36314 ( .IN1(n32865), .IN2(n32864), .IN3(n32863), .IN4(n32893), .Q(
        n32866) );
  MUX21X1 U36315 ( .IN1(n32867), .IN2(n32866), .S(\s11/msel/gnt_p0 [2]), .Q(
        n32876) );
  AO21X1 U36316 ( .IN1(n32869), .IN2(n32876), .IN3(n32868), .Q(n32875) );
  NOR2X0 U36317 ( .IN1(n32888), .IN2(n32900), .QN(n32873) );
  NOR2X0 U36318 ( .IN1(\s11/msel/gnt_p0 [0]), .IN2(n32911), .QN(n32901) );
  NOR2X0 U36319 ( .IN1(\s11/msel/gnt_p0 [0]), .IN2(n32901), .QN(n32871) );
  NAND2X0 U36320 ( .IN1(n32876), .IN2(n32882), .QN(n32870) );
  NOR2X0 U36321 ( .IN1(n32871), .IN2(n32870), .QN(n32872) );
  OR3X1 U36322 ( .IN1(n32873), .IN2(n32872), .IN3(n34452), .Q(n32874) );
  AO22X1 U36323 ( .IN1(\s11/msel/gnt_p0 [1]), .IN2(n32876), .IN3(n32875), 
        .IN4(n32874), .Q(n17718) );
  AO221X1 U36324 ( .IN1(\s11/msel/gnt_p0 [1]), .IN2(n32881), .IN3(n34668), 
        .IN4(n32883), .IN5(n34249), .Q(n32918) );
  NOR2X0 U36325 ( .IN1(\s11/msel/gnt_p0 [1]), .IN2(n32884), .QN(n32917) );
  OA21X1 U36326 ( .IN1(n32897), .IN2(n32883), .IN3(n32907), .Q(n32898) );
  OA21X1 U36327 ( .IN1(n32877), .IN2(n32898), .IN3(n32882), .Q(n32910) );
  NAND3X0 U36328 ( .IN1(n32878), .IN2(n32885), .IN3(n32900), .QN(n32879) );
  AO21X1 U36329 ( .IN1(n32910), .IN2(n32879), .IN3(n32893), .Q(n32892) );
  NAND2X0 U36330 ( .IN1(n32880), .IN2(n32900), .QN(n32908) );
  OA21X1 U36331 ( .IN1(n32882), .IN2(n32911), .IN3(n32881), .Q(n32902) );
  OA21X1 U36332 ( .IN1(n34249), .IN2(n32908), .IN3(n32902), .Q(n32896) );
  OAI21X1 U36333 ( .IN1(n32906), .IN2(n32896), .IN3(n32883), .QN(n32894) );
  NAND3X0 U36334 ( .IN1(\s11/msel/gnt_p0 [1]), .IN2(n32894), .IN3(n32884), 
        .QN(n32891) );
  INVX0 U36335 ( .INP(n32885), .ZN(n32886) );
  AO22X1 U36336 ( .IN1(n32898), .IN2(n32889), .IN3(n32888), .IN4(n32887), .Q(
        n32890) );
  NAND4X0 U36337 ( .IN1(\s11/msel/gnt_p0 [2]), .IN2(n32892), .IN3(n32891), 
        .IN4(n32890), .QN(n32916) );
  INVX0 U36338 ( .INP(n32893), .ZN(n32895) );
  NAND2X0 U36339 ( .IN1(n32895), .IN2(n32894), .QN(n32914) );
  NOR2X0 U36340 ( .IN1(n32897), .IN2(n32896), .QN(n32905) );
  INVX0 U36341 ( .INP(n32898), .ZN(n32899) );
  NAND3X0 U36342 ( .IN1(n32901), .IN2(n32900), .IN3(n32899), .QN(n32903) );
  NAND2X0 U36343 ( .IN1(n32903), .IN2(n32902), .QN(n32904) );
  NOR2X0 U36344 ( .IN1(n32905), .IN2(n32904), .QN(n32909) );
  AO221X1 U36345 ( .IN1(n32909), .IN2(n32908), .IN3(n32909), .IN4(n32907), 
        .IN5(n32906), .Q(n32913) );
  OR4X1 U36346 ( .IN1(n34668), .IN2(n34249), .IN3(n32911), .IN4(n32910), .Q(
        n32912) );
  NAND4X0 U36347 ( .IN1(n34452), .IN2(n32914), .IN3(n32913), .IN4(n32912), 
        .QN(n32915) );
  NAND2X0 U36348 ( .IN1(n32916), .IN2(n32915), .QN(n32921) );
  AO221X1 U36349 ( .IN1(n32918), .IN2(n32917), .IN3(n32918), .IN4(n32921), 
        .IN5(\s11/msel/gnt_p0 [2]), .Q(n32925) );
  NAND4X0 U36350 ( .IN1(\s11/msel/gnt_p0 [2]), .IN2(\s11/msel/gnt_p0 [0]), 
        .IN3(n32920), .IN4(n32919), .QN(n32924) );
  AO221X1 U36351 ( .IN1(n34249), .IN2(n32922), .IN3(n34249), .IN4(n34452), 
        .IN5(n32921), .Q(n32923) );
  NAND3X0 U36352 ( .IN1(n32925), .IN2(n32924), .IN3(n32923), .QN(n17717) );
  INVX0 U36353 ( .INP(n32926), .ZN(n32943) );
  OA22X1 U36354 ( .IN1(\s11/msel/gnt_p2 [1]), .IN2(n32935), .IN3(n34171), 
        .IN4(n34172), .Q(n32931) );
  AND3X1 U36355 ( .IN1(n32929), .IN2(n32928), .IN3(n32927), .Q(n32930) );
  AO221X1 U36356 ( .IN1(n32931), .IN2(\s11/msel/gnt_p2 [0]), .IN3(n32931), 
        .IN4(n32930), .IN5(n34401), .Q(n32942) );
  NAND2X0 U36357 ( .IN1(n34407), .IN2(n32932), .QN(n32939) );
  INVX0 U36358 ( .INP(n32933), .ZN(n32934) );
  NAND2X0 U36359 ( .IN1(n32935), .IN2(n32934), .QN(n34170) );
  OAI22X1 U36360 ( .IN1(n32937), .IN2(n34407), .IN3(n32936), .IN4(n34171), 
        .QN(n32938) );
  NAND4X0 U36361 ( .IN1(n32940), .IN2(n32939), .IN3(n34170), .IN4(n32938), 
        .QN(n32941) );
  NAND3X0 U36362 ( .IN1(n32943), .IN2(n32942), .IN3(n32941), .QN(n17716) );
  NOR2X0 U36363 ( .IN1(n32944), .IN2(n34379), .QN(n32945) );
  MUX21X1 U36364 ( .IN1(n34354), .IN2(s15_data_o[0]), .S(n32945), .Q(n17713)
         );
  MUX21X1 U36365 ( .IN1(n34509), .IN2(s15_data_o[1]), .S(n32945), .Q(n17712)
         );
  MUX21X1 U36366 ( .IN1(n34355), .IN2(s15_data_o[2]), .S(n32945), .Q(n17711)
         );
  MUX21X1 U36367 ( .IN1(n34508), .IN2(s15_data_o[3]), .S(n32945), .Q(n17710)
         );
  MUX21X1 U36368 ( .IN1(n34329), .IN2(s15_data_o[4]), .S(n32945), .Q(n17709)
         );
  MUX21X1 U36369 ( .IN1(n34541), .IN2(s15_data_o[5]), .S(n32945), .Q(n17708)
         );
  MUX21X1 U36370 ( .IN1(n34330), .IN2(s15_data_o[6]), .S(n32945), .Q(n17707)
         );
  MUX21X1 U36371 ( .IN1(n34507), .IN2(s15_data_o[7]), .S(n32945), .Q(n17706)
         );
  MUX21X1 U36372 ( .IN1(n34475), .IN2(s15_data_o[8]), .S(n32945), .Q(n17705)
         );
  MUX21X1 U36373 ( .IN1(n34642), .IN2(s15_data_o[9]), .S(n32945), .Q(n17704)
         );
  MUX21X1 U36374 ( .IN1(n34328), .IN2(s15_data_o[10]), .S(n32945), .Q(n17703)
         );
  MUX21X1 U36375 ( .IN1(n34506), .IN2(s15_data_o[11]), .S(n32945), .Q(n17702)
         );
  MUX21X1 U36376 ( .IN1(n34327), .IN2(s15_data_o[12]), .S(n32945), .Q(n17701)
         );
  MUX21X1 U36377 ( .IN1(n34540), .IN2(s15_data_o[13]), .S(n32945), .Q(n17700)
         );
  MUX21X1 U36378 ( .IN1(n34474), .IN2(s15_data_o[14]), .S(n32945), .Q(n17699)
         );
  MUX21X1 U36379 ( .IN1(n34643), .IN2(s15_data_o[15]), .S(n32945), .Q(n17698)
         );
  AO22X1 U36380 ( .IN1(n33003), .IN2(n34183), .IN3(n32980), .IN4(n32946), .Q(
        n32947) );
  NOR2X0 U36381 ( .IN1(n32947), .IN2(n32948), .QN(n32955) );
  INVX0 U36382 ( .INP(n32948), .ZN(n32951) );
  NAND2X0 U36383 ( .IN1(\s12/msel/gnt_p3 [1]), .IN2(n32968), .QN(n32950) );
  OA222X1 U36384 ( .IN1(n32951), .IN2(n32965), .IN3(n32950), .IN4(
        \s12/msel/gnt_p3 [0]), .IN5(n32949), .IN6(\s12/msel/gnt_p3 [1]), .Q(
        n32954) );
  NAND2X0 U36385 ( .IN1(n32994), .IN2(n32979), .QN(n32953) );
  NOR2X0 U36386 ( .IN1(n32953), .IN2(n32952), .QN(n34182) );
  NOR3X0 U36387 ( .IN1(n32955), .IN2(n32954), .IN3(n34182), .QN(n32961) );
  OA21X1 U36388 ( .IN1(\s12/msel/gnt_p3 [1]), .IN2(n32979), .IN3(n32956), .Q(
        n33013) );
  NAND2X0 U36389 ( .IN1(n34184), .IN2(n34183), .QN(n32959) );
  INVX0 U36390 ( .INP(n32976), .ZN(n32993) );
  AO221X1 U36391 ( .IN1(n34230), .IN2(n32962), .IN3(\s12/msel/gnt_p3 [1]), 
        .IN4(n32993), .IN5(n34450), .Q(n33001) );
  NAND2X0 U36392 ( .IN1(\s12/msel/gnt_p3 [0]), .IN2(\s12/msel/gnt_p3 [2]), 
        .QN(n33014) );
  NAND2X0 U36393 ( .IN1(n33001), .IN2(n33014), .QN(n32957) );
  NAND4X0 U36394 ( .IN1(n33013), .IN2(n32959), .IN3(n32958), .IN4(n32957), 
        .QN(n32960) );
  OA21X1 U36395 ( .IN1(\s12/msel/gnt_p3 [2]), .IN2(n32961), .IN3(n32960), .Q(
        n17697) );
  NAND2X0 U36396 ( .IN1(n32969), .IN2(n32968), .QN(n32970) );
  OA21X1 U36397 ( .IN1(n33004), .IN2(n33003), .IN3(n32978), .Q(n32992) );
  OA21X1 U36398 ( .IN1(n32980), .IN2(n32970), .IN3(n32992), .Q(n32972) );
  NOR2X0 U36399 ( .IN1(n32962), .IN2(n32970), .QN(n32963) );
  NAND2X0 U36400 ( .IN1(n32963), .IN2(\s12/msel/gnt_p3 [0]), .QN(n32964) );
  NAND2X0 U36401 ( .IN1(\s12/msel/gnt_p3 [0]), .IN2(n32976), .QN(n32971) );
  AO22X1 U36402 ( .IN1(n32972), .IN2(n32964), .IN3(n32971), .IN4(n32983), .Q(
        n32975) );
  NAND2X0 U36403 ( .IN1(n32979), .IN2(n32971), .QN(n32966) );
  AO21X1 U36404 ( .IN1(n32994), .IN2(n32966), .IN3(n32965), .Q(n32981) );
  AO21X1 U36405 ( .IN1(n32968), .IN2(n32981), .IN3(n32967), .Q(n32987) );
  NAND3X0 U36406 ( .IN1(\s12/msel/gnt_p3 [1]), .IN2(n32987), .IN3(n32969), 
        .QN(n32974) );
  OA21X1 U36407 ( .IN1(n32971), .IN2(n32970), .IN3(n32979), .Q(n32991) );
  AO221X1 U36408 ( .IN1(n32991), .IN2(n32993), .IN3(n32991), .IN4(n32972), 
        .IN5(n32988), .Q(n32973) );
  NAND4X0 U36409 ( .IN1(\s12/msel/gnt_p3 [2]), .IN2(n32975), .IN3(n32974), 
        .IN4(n32973), .QN(n33000) );
  OR2X1 U36410 ( .IN1(n33002), .IN2(n33005), .Q(n32986) );
  NAND2X0 U36411 ( .IN1(n32994), .IN2(n32976), .QN(n32977) );
  OR2X1 U36412 ( .IN1(n32978), .IN2(n32977), .Q(n32989) );
  NAND3X0 U36413 ( .IN1(n32980), .IN2(n33004), .IN3(n32979), .QN(n32982) );
  NAND2X0 U36414 ( .IN1(n32982), .IN2(n32981), .QN(n32985) );
  OR2X1 U36415 ( .IN1(n32983), .IN2(n32985), .Q(n32984) );
  OA221X1 U36416 ( .IN1(n32986), .IN2(n32989), .IN3(n32986), .IN4(n32985), 
        .IN5(n32984), .Q(n32998) );
  INVX0 U36417 ( .INP(n32987), .ZN(n32990) );
  AO221X1 U36418 ( .IN1(n32990), .IN2(n33005), .IN3(n32990), .IN4(n32989), 
        .IN5(n32988), .Q(n32997) );
  OAI21X1 U36419 ( .IN1(n32993), .IN2(n32992), .IN3(n32991), .QN(n32995) );
  NAND3X0 U36420 ( .IN1(\s12/msel/gnt_p3 [1]), .IN2(n32995), .IN3(n32994), 
        .QN(n32996) );
  NAND4X0 U36421 ( .IN1(n32998), .IN2(n34450), .IN3(n32997), .IN4(n32996), 
        .QN(n32999) );
  NAND2X0 U36422 ( .IN1(n33000), .IN2(n32999), .QN(n33012) );
  AND2X1 U36423 ( .IN1(n34269), .IN2(n33001), .Q(n33011) );
  NOR2X0 U36424 ( .IN1(n33003), .IN2(n33002), .QN(n33009) );
  AO221X1 U36425 ( .IN1(\s12/msel/gnt_p3 [1]), .IN2(n33005), .IN3(n34230), 
        .IN4(n33004), .IN5(n33012), .Q(n33006) );
  NAND2X0 U36426 ( .IN1(n33007), .IN2(n33006), .QN(n33008) );
  NOR2X0 U36427 ( .IN1(n33009), .IN2(n33008), .QN(n33010) );
  OAI222X1 U36428 ( .IN1(n33014), .IN2(n33013), .IN3(n33012), .IN4(n33011), 
        .IN5(n33010), .IN6(\s12/msel/gnt_p3 [2]), .QN(n17695) );
  NAND3X0 U36429 ( .IN1(n13561), .IN2(m6s12_cyc), .IN3(n34327), .QN(n33066) );
  NAND3X0 U36430 ( .IN1(n13613), .IN2(m5s12_cyc), .IN3(n34328), .QN(n33057) );
  NAND3X0 U36431 ( .IN1(n13481), .IN2(m7s12_cyc), .IN3(n34474), .QN(n33080) );
  OA221X1 U36432 ( .IN1(\s12/msel/gnt_p1 [1]), .IN2(n33066), .IN3(
        \s12/msel/gnt_p1 [1]), .IN4(n33057), .IN5(n33080), .Q(n33016) );
  NAND3X0 U36433 ( .IN1(n13665), .IN2(m4s12_cyc), .IN3(n34475), .QN(n33063) );
  MUX21X1 U36434 ( .IN1(n33063), .IN2(n33066), .S(\s12/msel/gnt_p1 [1]), .Q(
        n33082) );
  NAND3X0 U36435 ( .IN1(n13873), .IN2(m0s12_cyc), .IN3(n34354), .QN(n33078) );
  NAND3X0 U36436 ( .IN1(n13821), .IN2(m1s12_cyc), .IN3(n34355), .QN(n33054) );
  NAND2X0 U36437 ( .IN1(n33078), .IN2(n33054), .QN(n33032) );
  NAND3X0 U36438 ( .IN1(n13769), .IN2(m2s12_cyc), .IN3(n34329), .QN(n33065) );
  INVX0 U36439 ( .INP(n33065), .ZN(n33052) );
  NAND3X0 U36440 ( .IN1(n13717), .IN2(m3s12_cyc), .IN3(n34330), .QN(n33051) );
  INVX0 U36441 ( .INP(n33051), .ZN(n33035) );
  NOR2X0 U36442 ( .IN1(n33052), .IN2(n33035), .QN(n34189) );
  INVX0 U36443 ( .INP(n34189), .ZN(n33024) );
  OA22X1 U36444 ( .IN1(\s12/msel/gnt_p1 [0]), .IN2(n33082), .IN3(n33032), 
        .IN4(n33024), .Q(n33015) );
  NAND2X0 U36445 ( .IN1(n33016), .IN2(n33015), .QN(n33022) );
  NAND2X0 U36446 ( .IN1(\s12/msel/gnt_p1 [0]), .IN2(\s12/msel/gnt_p1 [1]), 
        .QN(n33079) );
  INVX0 U36447 ( .INP(n33079), .ZN(n33019) );
  NOR2X0 U36448 ( .IN1(\s12/msel/gnt_p1 [0]), .IN2(n34545), .QN(n33045) );
  AO22X1 U36449 ( .IN1(n33054), .IN2(n34189), .IN3(n33045), .IN4(n33051), .Q(
        n33018) );
  INVX0 U36450 ( .INP(n33078), .ZN(n33053) );
  NAND2X0 U36451 ( .IN1(n33053), .IN2(n34664), .QN(n33017) );
  OA22X1 U36452 ( .IN1(n33019), .IN2(n33018), .IN3(\s12/msel/gnt_p1 [1]), 
        .IN4(n33017), .Q(n33021) );
  NAND2X0 U36453 ( .IN1(n33066), .IN2(n33080), .QN(n33029) );
  NAND2X0 U36454 ( .IN1(n33063), .IN2(n33057), .QN(n33023) );
  NOR2X0 U36455 ( .IN1(n33029), .IN2(n33023), .QN(n34187) );
  AO21X1 U36456 ( .IN1(n33035), .IN2(n33019), .IN3(\s12/msel/gnt_p1 [2]), .Q(
        n33077) );
  AO21X1 U36457 ( .IN1(n33052), .IN2(n33045), .IN3(n33077), .Q(n33040) );
  NOR2X0 U36458 ( .IN1(n34187), .IN2(n33040), .QN(n33020) );
  AO22X1 U36459 ( .IN1(\s12/msel/gnt_p1 [2]), .IN2(n33022), .IN3(n33021), 
        .IN4(n33020), .Q(n17694) );
  NAND2X0 U36460 ( .IN1(\s12/msel/gnt_p1 [1]), .IN2(n33080), .QN(n33028) );
  INVX0 U36461 ( .INP(n33032), .ZN(n34188) );
  NAND2X0 U36462 ( .IN1(n34189), .IN2(n33023), .QN(n33030) );
  NOR2X0 U36463 ( .IN1(\s12/msel/gnt_p1 [1]), .IN2(n33029), .QN(n33026) );
  NAND2X0 U36464 ( .IN1(n34188), .IN2(n33024), .QN(n33025) );
  NAND2X0 U36465 ( .IN1(n33026), .IN2(n33025), .QN(n33027) );
  OA221X1 U36466 ( .IN1(n33028), .IN2(n34188), .IN3(n33028), .IN4(n33030), 
        .IN5(n33027), .Q(n33039) );
  INVX0 U36467 ( .INP(n33029), .ZN(n33033) );
  NAND2X0 U36468 ( .IN1(n34189), .IN2(n33033), .QN(n33031) );
  NAND4X0 U36469 ( .IN1(n34545), .IN2(n33054), .IN3(n33031), .IN4(n33030), 
        .QN(n33038) );
  NAND2X0 U36470 ( .IN1(n33033), .IN2(n33032), .QN(n33034) );
  NAND4X0 U36471 ( .IN1(\s12/msel/gnt_p1 [1]), .IN2(n33057), .IN3(n33063), 
        .IN4(n33034), .QN(n33037) );
  NAND2X0 U36472 ( .IN1(n33035), .IN2(n33045), .QN(n33036) );
  NAND4X0 U36473 ( .IN1(n34397), .IN2(n33038), .IN3(n33037), .IN4(n33036), 
        .QN(n33041) );
  OA21X1 U36474 ( .IN1(n33039), .IN2(n34397), .IN3(n33041), .Q(n33050) );
  AO221X1 U36475 ( .IN1(n33041), .IN2(\s12/msel/gnt_p1 [0]), .IN3(n33041), 
        .IN4(n33078), .IN5(n33040), .Q(n33049) );
  NOR2X0 U36476 ( .IN1(n33063), .IN2(\s12/msel/gnt_p1 [0]), .QN(n33043) );
  NAND2X0 U36477 ( .IN1(n33057), .IN2(n33050), .QN(n33042) );
  NOR2X0 U36478 ( .IN1(n33043), .IN2(n33042), .QN(n33044) );
  NOR2X0 U36479 ( .IN1(n33044), .IN2(n34397), .QN(n33047) );
  INVX0 U36480 ( .INP(n33066), .ZN(n33059) );
  NAND2X0 U36481 ( .IN1(n33059), .IN2(n33045), .QN(n33046) );
  NAND2X0 U36482 ( .IN1(n33047), .IN2(n33046), .QN(n33048) );
  AO22X1 U36483 ( .IN1(\s12/msel/gnt_p1 [1]), .IN2(n33050), .IN3(n33049), 
        .IN4(n33048), .Q(n17693) );
  INVX0 U36484 ( .INP(n33063), .ZN(n33070) );
  OA21X1 U36485 ( .IN1(n33070), .IN2(n33057), .IN3(n33051), .Q(n33055) );
  OA21X1 U36486 ( .IN1(n33052), .IN2(n33055), .IN3(n33054), .Q(n33071) );
  NOR3X0 U36487 ( .IN1(n33053), .IN2(n33071), .IN3(n33079), .QN(n33062) );
  OA21X1 U36488 ( .IN1(n33054), .IN2(n33053), .IN3(n33080), .Q(n33058) );
  INVX0 U36489 ( .INP(n33058), .ZN(n33064) );
  INVX0 U36490 ( .INP(n33055), .ZN(n33068) );
  OA221X1 U36491 ( .IN1(n33068), .IN2(\s12/msel/gnt_p1 [0]), .IN3(n33068), 
        .IN4(n33063), .IN5(n33065), .Q(n33056) );
  OA221X1 U36492 ( .IN1(n33064), .IN2(n33056), .IN3(n33064), .IN4(n33078), 
        .IN5(n33066), .Q(n33061) );
  OA21X1 U36493 ( .IN1(n33059), .IN2(n33058), .IN3(n33057), .Q(n33069) );
  NOR2X0 U36494 ( .IN1(\s12/msel/gnt_p1 [1]), .IN2(n33069), .QN(n33060) );
  NOR4X0 U36495 ( .IN1(n33062), .IN2(n33061), .IN3(n33060), .IN4(n34397), .QN(
        n33076) );
  OA221X1 U36496 ( .IN1(n33064), .IN2(\s12/msel/gnt_p1 [0]), .IN3(n33064), 
        .IN4(n33078), .IN5(n33063), .Q(n33067) );
  OA221X1 U36497 ( .IN1(n33068), .IN2(n33067), .IN3(n33068), .IN4(n33066), 
        .IN5(n33065), .Q(n33074) );
  NOR3X0 U36498 ( .IN1(n33070), .IN2(n33069), .IN3(n33079), .QN(n33073) );
  NOR2X0 U36499 ( .IN1(\s12/msel/gnt_p1 [1]), .IN2(n33071), .QN(n33072) );
  NOR4X0 U36500 ( .IN1(\s12/msel/gnt_p1 [2]), .IN2(n33074), .IN3(n33073), 
        .IN4(n33072), .QN(n33075) );
  NOR2X0 U36501 ( .IN1(n33076), .IN2(n33075), .QN(n33081) );
  AO221X1 U36502 ( .IN1(n33081), .IN2(\s12/msel/gnt_p1 [1]), .IN3(n33081), 
        .IN4(n33078), .IN5(n33077), .Q(n33085) );
  NOR2X0 U36503 ( .IN1(n33080), .IN2(n33079), .QN(n33084) );
  OA221X1 U36504 ( .IN1(\s12/msel/gnt_p1 [0]), .IN2(\s12/msel/gnt_p1 [2]), 
        .IN3(\s12/msel/gnt_p1 [0]), .IN4(n33082), .IN5(n33081), .Q(n33083) );
  AO221X1 U36505 ( .IN1(n33085), .IN2(n33084), .IN3(n33085), .IN4(n34397), 
        .IN5(n33083), .Q(n17692) );
  NAND3X0 U36506 ( .IN1(n13639), .IN2(n13613), .IN3(m5s12_cyc), .QN(n33138) );
  NAND3X0 U36507 ( .IN1(n13535), .IN2(n13481), .IN3(m7s12_cyc), .QN(n33151) );
  AOI221X1 U36508 ( .IN1(n34278), .IN2(n33138), .IN3(\s12/msel/gnt_p0 [1]), 
        .IN4(n33151), .IN5(n34382), .QN(n33177) );
  NAND3X0 U36509 ( .IN1(n13908), .IN2(n13873), .IN3(m0s12_cyc), .QN(n33175) );
  NAND3X0 U36510 ( .IN1(n13847), .IN2(n13821), .IN3(m1s12_cyc), .QN(n33173) );
  MUX21X1 U36511 ( .IN1(n33175), .IN2(n33173), .S(\s12/msel/gnt_p0 [0]), .Q(
        n33119) );
  NOR2X0 U36512 ( .IN1(n33119), .IN2(\s12/msel/gnt_p0 [1]), .QN(n33092) );
  NAND3X0 U36513 ( .IN1(n13743), .IN2(n13717), .IN3(m3s12_cyc), .QN(n33128) );
  NAND2X0 U36514 ( .IN1(\s12/msel/gnt_p0 [0]), .IN2(\s12/msel/gnt_p0 [1]), 
        .QN(n33089) );
  NOR2X0 U36515 ( .IN1(n33128), .IN2(n33089), .QN(n33182) );
  NOR2X0 U36516 ( .IN1(\s12/msel/gnt_p0 [2]), .IN2(n33182), .QN(n33087) );
  NAND3X0 U36517 ( .IN1(n13795), .IN2(n13769), .IN3(m2s12_cyc), .QN(n33147) );
  INVX0 U36518 ( .INP(n33147), .ZN(n33165) );
  NOR2X0 U36519 ( .IN1(\s12/msel/gnt_p0 [0]), .IN2(n34278), .QN(n33137) );
  NAND2X0 U36520 ( .IN1(n33165), .IN2(n33137), .QN(n33086) );
  NAND2X0 U36521 ( .IN1(n33087), .IN2(n33086), .QN(n33117) );
  NAND3X0 U36522 ( .IN1(n13691), .IN2(n13665), .IN3(m4s12_cyc), .QN(n33130) );
  AND2X1 U36523 ( .IN1(n33138), .IN2(n33130), .Q(n33110) );
  NAND3X0 U36524 ( .IN1(n13587), .IN2(n13561), .IN3(m6s12_cyc), .QN(n33152) );
  INVX0 U36525 ( .INP(n33152), .ZN(n33143) );
  INVX0 U36526 ( .INP(n33151), .ZN(n33132) );
  NOR2X0 U36527 ( .IN1(n33143), .IN2(n33132), .QN(n33098) );
  INVX0 U36528 ( .INP(n33128), .ZN(n33140) );
  INVX0 U36529 ( .INP(n33137), .ZN(n33088) );
  INVX0 U36530 ( .INP(n33173), .ZN(n33145) );
  NAND2X0 U36531 ( .IN1(n34443), .IN2(n34278), .QN(n33162) );
  NAND2X0 U36532 ( .IN1(\s12/msel/gnt_p0 [0]), .IN2(n34278), .QN(n33093) );
  OA21X1 U36533 ( .IN1(n33145), .IN2(n33162), .IN3(n33093), .Q(n33108) );
  NAND2X0 U36534 ( .IN1(n33147), .IN2(n33128), .QN(n33112) );
  OA22X1 U36535 ( .IN1(n33140), .IN2(n33088), .IN3(n33108), .IN4(n33112), .Q(
        n33090) );
  AO22X1 U36536 ( .IN1(n33110), .IN2(n33098), .IN3(n33090), .IN4(n33089), .Q(
        n33091) );
  NOR3X0 U36537 ( .IN1(n33092), .IN2(n33117), .IN3(n33091), .QN(n33097) );
  INVX0 U36538 ( .INP(n33130), .ZN(n33166) );
  MUX21X1 U36539 ( .IN1(n33166), .IN2(n33143), .S(\s12/msel/gnt_p0 [1]), .Q(
        n33176) );
  AND3X1 U36540 ( .IN1(\s12/msel/gnt_p0 [2]), .IN2(n33176), .IN3(n34443), .Q(
        n33096) );
  NAND2X0 U36541 ( .IN1(n33175), .IN2(n33173), .QN(n33101) );
  NOR2X0 U36542 ( .IN1(n33112), .IN2(n33101), .QN(n33094) );
  NOR2X0 U36543 ( .IN1(n33143), .IN2(n33093), .QN(n33136) );
  OAI21X1 U36544 ( .IN1(\s12/msel/gnt_p0 [1]), .IN2(n33136), .IN3(n33151), 
        .QN(n33105) );
  INVX0 U36545 ( .INP(n33098), .ZN(n33111) );
  OA221X1 U36546 ( .IN1(n33094), .IN2(n33105), .IN3(n33094), .IN4(n33111), 
        .IN5(\s12/msel/gnt_p0 [2]), .Q(n33095) );
  OR4X1 U36547 ( .IN1(n33177), .IN2(n33097), .IN3(n33096), .IN4(n33095), .Q(
        n17691) );
  NOR2X0 U36548 ( .IN1(n33112), .IN2(n33111), .QN(n33100) );
  NAND2X0 U36549 ( .IN1(n33098), .IN2(n33101), .QN(n33107) );
  NAND2X0 U36550 ( .IN1(n33107), .IN2(n33138), .QN(n33099) );
  NOR2X0 U36551 ( .IN1(n33100), .IN2(n33099), .QN(n33106) );
  INVX0 U36552 ( .INP(n33136), .ZN(n33103) );
  INVX0 U36553 ( .INP(n33101), .ZN(n33102) );
  OA221X1 U36554 ( .IN1(n33112), .IN2(n33110), .IN3(n33112), .IN4(n33103), 
        .IN5(n33102), .Q(n33104) );
  OA22X1 U36555 ( .IN1(n33106), .IN2(n33162), .IN3(n33105), .IN4(n33104), .Q(
        n33116) );
  NAND4X0 U36556 ( .IN1(\s12/msel/gnt_p0 [1]), .IN2(n33130), .IN3(n33138), 
        .IN4(n33107), .QN(n33115) );
  NAND2X0 U36557 ( .IN1(n33140), .IN2(n33137), .QN(n33114) );
  INVX0 U36558 ( .INP(n33108), .ZN(n33109) );
  OAI221X1 U36559 ( .IN1(n33112), .IN2(n33111), .IN3(n33112), .IN4(n33110), 
        .IN5(n33109), .QN(n33113) );
  NAND4X0 U36560 ( .IN1(n34382), .IN2(n33115), .IN3(n33114), .IN4(n33113), 
        .QN(n33118) );
  OA21X1 U36561 ( .IN1(n33116), .IN2(n34382), .IN3(n33118), .Q(n33127) );
  AO21X1 U36562 ( .IN1(n33119), .IN2(n33118), .IN3(n33117), .Q(n33126) );
  NOR2X0 U36563 ( .IN1(\s12/msel/gnt_p0 [0]), .IN2(n33130), .QN(n33121) );
  NAND2X0 U36564 ( .IN1(n33127), .IN2(n33138), .QN(n33120) );
  NOR2X0 U36565 ( .IN1(n33121), .IN2(n33120), .QN(n33122) );
  NOR2X0 U36566 ( .IN1(n33122), .IN2(n34382), .QN(n33124) );
  NAND2X0 U36567 ( .IN1(n33143), .IN2(n33137), .QN(n33123) );
  NAND2X0 U36568 ( .IN1(n33124), .IN2(n33123), .QN(n33125) );
  AO22X1 U36569 ( .IN1(\s12/msel/gnt_p0 [1]), .IN2(n33127), .IN3(n33126), 
        .IN4(n33125), .Q(n17690) );
  OA21X1 U36570 ( .IN1(n33166), .IN2(n33138), .IN3(n33128), .Q(n33144) );
  NAND2X0 U36571 ( .IN1(n33175), .IN2(n33147), .QN(n33129) );
  NOR2X0 U36572 ( .IN1(n33144), .IN2(n33129), .QN(n33135) );
  INVX0 U36573 ( .INP(n33129), .ZN(n33141) );
  NAND3X0 U36574 ( .IN1(\s12/msel/gnt_p0 [0]), .IN2(n33141), .IN3(n33130), 
        .QN(n33133) );
  INVX0 U36575 ( .INP(n33175), .ZN(n33131) );
  NOR2X0 U36576 ( .IN1(n33131), .IN2(n33173), .QN(n33153) );
  NOR2X0 U36577 ( .IN1(n33153), .IN2(n33132), .QN(n33139) );
  NAND2X0 U36578 ( .IN1(n33133), .IN2(n33139), .QN(n33134) );
  OA22X1 U36579 ( .IN1(n33137), .IN2(n33136), .IN3(n33135), .IN4(n33134), .Q(
        n33172) );
  OA21X1 U36580 ( .IN1(n33143), .IN2(n33139), .IN3(n33138), .Q(n33167) );
  NAND3X0 U36581 ( .IN1(n33141), .IN2(n33140), .IN3(n33152), .QN(n33142) );
  AO21X1 U36582 ( .IN1(n33167), .IN2(n33142), .IN3(n33162), .Q(n33149) );
  NOR2X0 U36583 ( .IN1(n33143), .IN2(n33166), .QN(n33154) );
  INVX0 U36584 ( .INP(n33144), .ZN(n33155) );
  AO21X1 U36585 ( .IN1(\s12/msel/gnt_p0 [0]), .IN2(n33154), .IN3(n33155), .Q(
        n33146) );
  AO21X1 U36586 ( .IN1(n33147), .IN2(n33146), .IN3(n33145), .Q(n33161) );
  NAND3X0 U36587 ( .IN1(\s12/msel/gnt_p0 [1]), .IN2(n33161), .IN3(n33175), 
        .QN(n33148) );
  NAND3X0 U36588 ( .IN1(\s12/msel/gnt_p0 [2]), .IN2(n33149), .IN3(n33148), 
        .QN(n33171) );
  INVX0 U36589 ( .INP(n33154), .ZN(n33150) );
  NOR2X0 U36590 ( .IN1(n33151), .IN2(n33150), .QN(n33160) );
  NAND3X0 U36591 ( .IN1(n33153), .IN2(n33152), .IN3(n33130), .QN(n33158) );
  AND3X1 U36592 ( .IN1(n33175), .IN2(n33154), .IN3(\s12/msel/gnt_p0 [0]), .Q(
        n33156) );
  NOR2X0 U36593 ( .IN1(n33156), .IN2(n33155), .QN(n33157) );
  NAND2X0 U36594 ( .IN1(n33158), .IN2(n33157), .QN(n33159) );
  NOR2X0 U36595 ( .IN1(n33160), .IN2(n33159), .QN(n33164) );
  INVX0 U36596 ( .INP(n33161), .ZN(n33163) );
  OA22X1 U36597 ( .IN1(n33165), .IN2(n33164), .IN3(n33163), .IN4(n33162), .Q(
        n33169) );
  OR4X1 U36598 ( .IN1(n34278), .IN2(n34443), .IN3(n33167), .IN4(n33166), .Q(
        n33168) );
  NAND2X0 U36599 ( .IN1(n33169), .IN2(n33168), .QN(n33170) );
  OA22X1 U36600 ( .IN1(n33172), .IN2(n33171), .IN3(\s12/msel/gnt_p0 [2]), 
        .IN4(n33170), .Q(n33178) );
  NOR2X0 U36601 ( .IN1(n34443), .IN2(n33173), .QN(n33174) );
  AO222X1 U36602 ( .IN1(n33178), .IN2(\s12/msel/gnt_p0 [1]), .IN3(n33178), 
        .IN4(n33175), .IN5(n34278), .IN6(n33174), .Q(n33181) );
  NOR2X0 U36603 ( .IN1(n33176), .IN2(n34382), .QN(n33179) );
  OA22X1 U36604 ( .IN1(\s12/msel/gnt_p0 [0]), .IN2(n33179), .IN3(n33178), 
        .IN4(n33177), .Q(n33180) );
  AO221X1 U36605 ( .IN1(n34382), .IN2(n33182), .IN3(n34382), .IN4(n33181), 
        .IN5(n33180), .Q(n17689) );
  NAND2X0 U36606 ( .IN1(n33219), .IN2(n33220), .QN(n33204) );
  NAND2X0 U36607 ( .IN1(n33183), .IN2(n33209), .QN(n33214) );
  NAND2X0 U36608 ( .IN1(n33191), .IN2(n33184), .QN(n33217) );
  NOR2X0 U36609 ( .IN1(n33214), .IN2(n33217), .QN(n34185) );
  AO221X1 U36610 ( .IN1(n34244), .IN2(n33186), .IN3(n34244), .IN4(n33185), 
        .IN5(n34185), .Q(n33187) );
  AO221X1 U36611 ( .IN1(n33189), .IN2(n33204), .IN3(n33189), .IN4(n33188), 
        .IN5(n33187), .Q(n33202) );
  INVX0 U36612 ( .INP(n33190), .ZN(n33194) );
  AND2X1 U36613 ( .IN1(n34422), .IN2(n33191), .Q(n33216) );
  INVX0 U36614 ( .INP(n33214), .ZN(n33218) );
  AO22X1 U36615 ( .IN1(n33216), .IN2(n33218), .IN3(n33196), .IN4(n33209), .Q(
        n33193) );
  NAND2X0 U36616 ( .IN1(n33192), .IN2(n34244), .QN(n33233) );
  OA22X1 U36617 ( .IN1(n33194), .IN2(n33193), .IN3(\s12/msel/gnt_p2 [1]), 
        .IN4(n33233), .Q(n33201) );
  NAND2X0 U36618 ( .IN1(n33227), .IN2(n33230), .QN(n33203) );
  NOR2X0 U36619 ( .IN1(n33203), .IN2(n33204), .QN(n34186) );
  NOR2X0 U36620 ( .IN1(\s12/msel/gnt_p2 [2]), .IN2(n33195), .QN(n33199) );
  NAND2X0 U36621 ( .IN1(n33197), .IN2(n33196), .QN(n33198) );
  NAND2X0 U36622 ( .IN1(n33199), .IN2(n33198), .QN(n33234) );
  NOR2X0 U36623 ( .IN1(n34186), .IN2(n33234), .QN(n33200) );
  AO22X1 U36624 ( .IN1(\s12/msel/gnt_p2 [2]), .IN2(n33202), .IN3(n33201), 
        .IN4(n33200), .Q(n17688) );
  INVX0 U36625 ( .INP(n33203), .ZN(n33206) );
  NAND2X0 U36626 ( .IN1(n33204), .IN2(n33206), .QN(n33208) );
  INVX0 U36627 ( .INP(n33208), .ZN(n33215) );
  INVX0 U36628 ( .INP(n33217), .ZN(n33207) );
  OA21X1 U36629 ( .IN1(n33207), .IN2(n33204), .IN3(n33206), .Q(n33205) );
  NOR2X0 U36630 ( .IN1(n33205), .IN2(n34244), .QN(n33212) );
  NAND2X0 U36631 ( .IN1(n33207), .IN2(n33206), .QN(n33221) );
  NAND3X0 U36632 ( .IN1(n33209), .IN2(n33221), .IN3(n33208), .QN(n33210) );
  NAND2X0 U36633 ( .IN1(\s12/msel/gnt_p2 [1]), .IN2(n33210), .QN(n33211) );
  NOR2X0 U36634 ( .IN1(n33212), .IN2(n33211), .QN(n33213) );
  AO221X1 U36635 ( .IN1(n33216), .IN2(n33215), .IN3(n33216), .IN4(n33214), 
        .IN5(n33213), .Q(n33226) );
  NOR2X0 U36636 ( .IN1(n33218), .IN2(n33217), .QN(n33224) );
  OAI221X1 U36637 ( .IN1(n34422), .IN2(n33221), .IN3(\s12/msel/gnt_p2 [1]), 
        .IN4(n33220), .IN5(n33219), .QN(n33223) );
  OA22X1 U36638 ( .IN1(n33224), .IN2(n33223), .IN3(n33227), .IN4(n33222), .Q(
        n33225) );
  MUX21X1 U36639 ( .IN1(n33226), .IN2(n33225), .S(\s12/msel/gnt_p2 [2]), .Q(
        n33237) );
  INVX0 U36640 ( .INP(n33227), .ZN(n33228) );
  NAND2X0 U36641 ( .IN1(\s12/msel/gnt_p2 [0]), .IN2(\s12/msel/gnt_p2 [2]), 
        .QN(n33229) );
  NOR2X0 U36642 ( .IN1(n33228), .IN2(n33229), .QN(n33236) );
  OA221X1 U36643 ( .IN1(n33231), .IN2(n33230), .IN3(n33231), .IN4(n33237), 
        .IN5(n33229), .Q(n33232) );
  OA221X1 U36644 ( .IN1(n33234), .IN2(n33237), .IN3(n33234), .IN4(n33233), 
        .IN5(n33232), .Q(n33235) );
  AO221X1 U36645 ( .IN1(n33237), .IN2(\s12/msel/gnt_p2 [1]), .IN3(n33237), 
        .IN4(n33236), .IN5(n33235), .Q(n17687) );
  NOR2X0 U36646 ( .IN1(n33238), .IN2(n34379), .QN(n33239) );
  MUX21X1 U36647 ( .IN1(n34356), .IN2(s15_data_o[0]), .S(n33239), .Q(n17685)
         );
  MUX21X1 U36648 ( .IN1(n34542), .IN2(s15_data_o[1]), .S(n33239), .Q(n17684)
         );
  MUX21X1 U36649 ( .IN1(n34332), .IN2(s15_data_o[2]), .S(n33239), .Q(n17683)
         );
  MUX21X1 U36650 ( .IN1(n34510), .IN2(s15_data_o[3]), .S(n33239), .Q(n17682)
         );
  MUX21X1 U36651 ( .IN1(n34480), .IN2(s15_data_o[4]), .S(n33239), .Q(n17681)
         );
  MUX21X1 U36652 ( .IN1(n34645), .IN2(s15_data_o[5]), .S(n33239), .Q(n17680)
         );
  MUX21X1 U36653 ( .IN1(n34546), .IN2(s15_data_o[6]), .S(n33239), .Q(n17679)
         );
  MUX21X1 U36654 ( .IN1(n34651), .IN2(s15_data_o[7]), .S(n33239), .Q(n17678)
         );
  MUX21X1 U36655 ( .IN1(n34333), .IN2(s15_data_o[8]), .S(n33239), .Q(n17677)
         );
  MUX21X1 U36656 ( .IN1(n34543), .IN2(s15_data_o[9]), .S(n33239), .Q(n17676)
         );
  MUX21X1 U36657 ( .IN1(n34476), .IN2(s15_data_o[10]), .S(n33239), .Q(n17675)
         );
  MUX21X1 U36658 ( .IN1(n34644), .IN2(s15_data_o[11]), .S(n33239), .Q(n17674)
         );
  MUX21X1 U36659 ( .IN1(n34331), .IN2(s15_data_o[12]), .S(n33239), .Q(n17673)
         );
  MUX21X1 U36660 ( .IN1(n34511), .IN2(s15_data_o[13]), .S(n33239), .Q(n17672)
         );
  MUX21X1 U36661 ( .IN1(n34634), .IN2(s15_data_o[14]), .S(n33239), .Q(n17671)
         );
  MUX21X1 U36662 ( .IN1(n34586), .IN2(s15_data_o[15]), .S(n33239), .Q(n17670)
         );
  NAND2X0 U36663 ( .IN1(m5s13_cyc), .IN2(n34644), .QN(n33451) );
  NOR2X0 U36664 ( .IN1(n13640), .IN2(n33451), .QN(n33289) );
  NAND2X0 U36665 ( .IN1(m7s13_cyc), .IN2(n34586), .QN(n33240) );
  NOR2X0 U36666 ( .IN1(n13536), .IN2(n33240), .QN(n33277) );
  MUX21X1 U36667 ( .IN1(n33289), .IN2(n33277), .S(\s13/msel/gnt_p3 [1]), .Q(
        n33312) );
  NAND3X0 U36668 ( .IN1(m4s13_cyc), .IN2(n34333), .IN3(n34543), .QN(n33292) );
  NAND3X0 U36669 ( .IN1(m6s13_cyc), .IN2(n34331), .IN3(n34511), .QN(n33299) );
  MUX21X1 U36670 ( .IN1(n33292), .IN2(n33299), .S(\s13/msel/gnt_p3 [1]), .Q(
        n33271) );
  INVX0 U36671 ( .INP(n33277), .ZN(n33282) );
  NAND2X0 U36672 ( .IN1(n33299), .IN2(n33282), .QN(n33255) );
  INVX0 U36673 ( .INP(n33255), .ZN(n33247) );
  OA22X1 U36674 ( .IN1(\s13/msel/gnt_p3 [0]), .IN2(n33271), .IN3(
        \s13/msel/gnt_p3 [1]), .IN4(n33247), .Q(n33242) );
  NAND3X0 U36675 ( .IN1(m0s13_cyc), .IN2(n34356), .IN3(n34542), .QN(n33280) );
  INVX0 U36676 ( .INP(n33280), .ZN(n33302) );
  NAND3X0 U36677 ( .IN1(m1s13_cyc), .IN2(n34332), .IN3(n34510), .QN(n33273) );
  INVX0 U36678 ( .INP(n33273), .ZN(n33304) );
  NOR2X0 U36679 ( .IN1(n33302), .IN2(n33304), .QN(n34198) );
  NAND2X0 U36680 ( .IN1(m2s13_cyc), .IN2(n34645), .QN(n33448) );
  NOR2X0 U36681 ( .IN1(n13796), .IN2(n33448), .QN(n33303) );
  NAND2X0 U36682 ( .IN1(m3s13_cyc), .IN2(n34651), .QN(n33449) );
  NOR2X0 U36683 ( .IN1(n13744), .IN2(n33449), .QN(n33281) );
  NOR2X0 U36684 ( .IN1(n33303), .IN2(n33281), .QN(n34197) );
  NAND2X0 U36685 ( .IN1(n34198), .IN2(n34197), .QN(n33241) );
  NAND2X0 U36686 ( .IN1(n33242), .IN2(n33241), .QN(n33246) );
  INVX0 U36687 ( .INP(n33289), .ZN(n33274) );
  NAND2X0 U36688 ( .IN1(n33292), .IN2(n33274), .QN(n33250) );
  NOR2X0 U36689 ( .IN1(n33250), .IN2(n33255), .QN(n34196) );
  AO21X1 U36690 ( .IN1(n33302), .IN2(n34267), .IN3(n33304), .Q(n33265) );
  OA22X1 U36691 ( .IN1(n33281), .IN2(n34384), .IN3(n33265), .IN4(
        \s13/msel/gnt_p3 [1]), .Q(n33244) );
  NOR2X0 U36692 ( .IN1(n34267), .IN2(n34384), .QN(n33264) );
  NOR2X0 U36693 ( .IN1(n33264), .IN2(n34197), .QN(n33243) );
  NOR4X0 U36694 ( .IN1(\s13/msel/gnt_p3 [2]), .IN2(n34196), .IN3(n33244), 
        .IN4(n33243), .QN(n33245) );
  AO221X1 U36695 ( .IN1(\s13/msel/gnt_p3 [2]), .IN2(n33312), .IN3(
        \s13/msel/gnt_p3 [2]), .IN4(n33246), .IN5(n33245), .Q(n17669) );
  NOR2X0 U36696 ( .IN1(n34267), .IN2(n34431), .QN(n33311) );
  NOR2X0 U36697 ( .IN1(\s13/msel/gnt_p3 [0]), .IN2(n34384), .QN(n33293) );
  NAND4X0 U36698 ( .IN1(n33293), .IN2(n34198), .IN3(n33292), .IN4(n33274), 
        .QN(n33254) );
  OA221X1 U36699 ( .IN1(n34197), .IN2(\s13/msel/gnt_p3 [1]), .IN3(n34197), 
        .IN4(\s13/msel/gnt_p3 [0]), .IN5(n34431), .Q(n33249) );
  NAND2X0 U36700 ( .IN1(n33264), .IN2(n33280), .QN(n33275) );
  AO221X1 U36701 ( .IN1(n33247), .IN2(n33304), .IN3(n33247), .IN4(n33275), 
        .IN5(n33250), .Q(n33248) );
  NAND3X0 U36702 ( .IN1(n33254), .IN2(n33249), .IN3(n33248), .QN(n33262) );
  NAND2X0 U36703 ( .IN1(n34267), .IN2(n34384), .QN(n33287) );
  NOR2X0 U36704 ( .IN1(n33289), .IN2(n33287), .QN(n33252) );
  OA221X1 U36705 ( .IN1(n33255), .IN2(n34198), .IN3(n33255), .IN4(n33303), 
        .IN5(n33252), .Q(n33260) );
  OA21X1 U36706 ( .IN1(n33250), .IN2(n34384), .IN3(n34197), .Q(n33251) );
  OAI22X1 U36707 ( .IN1(n34267), .IN2(n33251), .IN3(n34197), .IN4(n34384), 
        .QN(n33253) );
  OA221X1 U36708 ( .IN1(n33253), .IN2(n33281), .IN3(n33253), .IN4(n33252), 
        .IN5(n34198), .Q(n33259) );
  NOR2X0 U36709 ( .IN1(\s13/msel/gnt_p3 [1]), .IN2(n34267), .QN(n33257) );
  INVX0 U36710 ( .INP(n33254), .ZN(n33256) );
  OA22X1 U36711 ( .IN1(n33293), .IN2(n33257), .IN3(n33256), .IN4(n33255), .Q(
        n33258) );
  OR4X1 U36712 ( .IN1(n33260), .IN2(n33259), .IN3(n33258), .IN4(n34431), .Q(
        n33261) );
  NAND2X0 U36713 ( .IN1(n33262), .IN2(n33261), .QN(n33266) );
  OAI22X1 U36714 ( .IN1(n34384), .IN2(n33282), .IN3(n33266), .IN4(n33289), 
        .QN(n33263) );
  NAND2X0 U36715 ( .IN1(n33311), .IN2(n33263), .QN(n33270) );
  NAND2X0 U36716 ( .IN1(n33281), .IN2(n33264), .QN(n33305) );
  AO221X1 U36717 ( .IN1(n33305), .IN2(n33266), .IN3(n33305), .IN4(n33265), 
        .IN5(\s13/msel/gnt_p3 [2]), .Q(n33269) );
  NAND3X0 U36718 ( .IN1(\s13/msel/gnt_p3 [2]), .IN2(n34267), .IN3(n33292), 
        .QN(n33267) );
  AO21X1 U36719 ( .IN1(n34384), .IN2(n33267), .IN3(n33266), .Q(n33268) );
  NAND3X0 U36720 ( .IN1(n33270), .IN2(n33269), .IN3(n33268), .QN(n17668) );
  AO21X1 U36721 ( .IN1(\s13/msel/gnt_p3 [2]), .IN2(n33271), .IN3(
        \s13/msel/gnt_p3 [0]), .Q(n33310) );
  OA221X1 U36722 ( .IN1(n33289), .IN2(\s13/msel/gnt_p3 [0]), .IN3(n33289), 
        .IN4(n33299), .IN5(n33292), .Q(n33272) );
  NOR2X0 U36723 ( .IN1(n33281), .IN2(n33272), .QN(n33285) );
  OA21X1 U36724 ( .IN1(n33303), .IN2(n33285), .IN3(n33273), .Q(n33288) );
  OA22X1 U36725 ( .IN1(n33288), .IN2(n33275), .IN3(n33274), .IN4(n33287), .Q(
        n33276) );
  NAND2X0 U36726 ( .IN1(\s13/msel/gnt_p3 [2]), .IN2(n33276), .QN(n33300) );
  NOR2X0 U36727 ( .IN1(n33303), .IN2(n33302), .QN(n33279) );
  OA21X1 U36728 ( .IN1(\s13/msel/gnt_p3 [0]), .IN2(n33289), .IN3(n33292), .Q(
        n33278) );
  AO21X1 U36729 ( .IN1(n33304), .IN2(n33280), .IN3(n33277), .Q(n33291) );
  AO221X1 U36730 ( .IN1(n33279), .IN2(n33281), .IN3(n33279), .IN4(n33278), 
        .IN5(n33291), .Q(n33298) );
  NOR3X0 U36731 ( .IN1(n33281), .IN2(n33289), .IN3(n33280), .QN(n33284) );
  NAND2X0 U36732 ( .IN1(n33292), .IN2(n33299), .QN(n33283) );
  OA22X1 U36733 ( .IN1(n33285), .IN2(n33284), .IN3(n33283), .IN4(n33282), .Q(
        n33286) );
  OA22X1 U36734 ( .IN1(n33288), .IN2(n33287), .IN3(n33303), .IN4(n33286), .Q(
        n33296) );
  AO21X1 U36735 ( .IN1(n33299), .IN2(n33291), .IN3(n33289), .Q(n33290) );
  NAND3X0 U36736 ( .IN1(\s13/msel/gnt_p3 [1]), .IN2(n33290), .IN3(n33292), 
        .QN(n33295) );
  NAND4X0 U36737 ( .IN1(n33293), .IN2(n33292), .IN3(n33299), .IN4(n33291), 
        .QN(n33294) );
  NAND4X0 U36738 ( .IN1(n33296), .IN2(n34431), .IN3(n33295), .IN4(n33294), 
        .QN(n33297) );
  OA221X1 U36739 ( .IN1(n33300), .IN2(n33299), .IN3(n33300), .IN4(n33298), 
        .IN5(n33297), .Q(n33309) );
  INVX0 U36740 ( .INP(n33309), .ZN(n33301) );
  AO221X1 U36741 ( .IN1(\s13/msel/gnt_p3 [1]), .IN2(n33303), .IN3(n34384), 
        .IN4(n33302), .IN5(n33301), .Q(n33307) );
  NAND3X0 U36742 ( .IN1(\s13/msel/gnt_p3 [0]), .IN2(n33304), .IN3(n34384), 
        .QN(n33306) );
  NAND3X0 U36743 ( .IN1(n33307), .IN2(n33306), .IN3(n33305), .QN(n33308) );
  AO222X1 U36744 ( .IN1(n33312), .IN2(n33311), .IN3(n33310), .IN4(n33309), 
        .IN5(n33308), .IN6(n34431), .Q(n17667) );
  NAND3X0 U36745 ( .IN1(n13482), .IN2(m7s13_cyc), .IN3(n34634), .QN(n33345) );
  NAND2X0 U36746 ( .IN1(\s13/msel/gnt_p1 [1]), .IN2(n33345), .QN(n33372) );
  NAND3X0 U36747 ( .IN1(n13614), .IN2(m5s13_cyc), .IN3(n34476), .QN(n33347) );
  NAND2X0 U36748 ( .IN1(n34411), .IN2(n33347), .QN(n33373) );
  NAND3X0 U36749 ( .IN1(n13562), .IN2(m6s13_cyc), .IN3(n34331), .QN(n33313) );
  NAND2X0 U36750 ( .IN1(n33313), .IN2(n33345), .QN(n33326) );
  NAND3X0 U36751 ( .IN1(n13822), .IN2(m1s13_cyc), .IN3(n34332), .QN(n33346) );
  INVX0 U36752 ( .INP(n33346), .ZN(n33344) );
  NAND3X0 U36753 ( .IN1(n13874), .IN2(m0s13_cyc), .IN3(n34356), .QN(n33374) );
  INVX0 U36754 ( .INP(n33374), .ZN(n33357) );
  NOR2X0 U36755 ( .IN1(n33344), .IN2(n33357), .QN(n34202) );
  NAND3X0 U36756 ( .IN1(n13718), .IN2(m3s13_cyc), .IN3(n34546), .QN(n33351) );
  INVX0 U36757 ( .INP(n33351), .ZN(n33316) );
  NAND3X0 U36758 ( .IN1(n13770), .IN2(m2s13_cyc), .IN3(n34480), .QN(n33348) );
  INVX0 U36759 ( .INP(n33348), .ZN(n33359) );
  NOR2X0 U36760 ( .IN1(n33316), .IN2(n33359), .QN(n34203) );
  NAND3X0 U36761 ( .IN1(n13666), .IN2(m4s13_cyc), .IN3(n34333), .QN(n33349) );
  INVX0 U36762 ( .INP(n33349), .ZN(n33365) );
  INVX0 U36763 ( .INP(n33313), .ZN(n33361) );
  MUX21X1 U36764 ( .IN1(n33365), .IN2(n33361), .S(\s13/msel/gnt_p1 [1]), .Q(
        n33371) );
  AO22X1 U36765 ( .IN1(n34202), .IN2(n34203), .IN3(n34248), .IN4(n33371), .Q(
        n33314) );
  AO221X1 U36766 ( .IN1(n33372), .IN2(n33373), .IN3(n33372), .IN4(n33326), 
        .IN5(n33314), .Q(n33320) );
  OA21X1 U36767 ( .IN1(\s13/msel/gnt_p1 [0]), .IN2(n33374), .IN3(n33346), .Q(
        n33335) );
  NOR2X0 U36768 ( .IN1(n34248), .IN2(n34411), .QN(n33315) );
  OA22X1 U36769 ( .IN1(\s13/msel/gnt_p1 [1]), .IN2(n33335), .IN3(n33315), 
        .IN4(n34203), .Q(n33319) );
  NAND2X0 U36770 ( .IN1(n33349), .IN2(n33347), .QN(n33322) );
  NOR2X0 U36771 ( .IN1(n33326), .IN2(n33322), .QN(n34201) );
  NAND2X0 U36772 ( .IN1(n33316), .IN2(n33315), .QN(n33377) );
  NAND3X0 U36773 ( .IN1(\s13/msel/gnt_p1 [1]), .IN2(n33359), .IN3(n34248), 
        .QN(n33317) );
  NAND3X0 U36774 ( .IN1(n34471), .IN2(n33377), .IN3(n33317), .QN(n33334) );
  NOR2X0 U36775 ( .IN1(n34201), .IN2(n33334), .QN(n33318) );
  AO22X1 U36776 ( .IN1(\s13/msel/gnt_p1 [2]), .IN2(n33320), .IN3(n33319), 
        .IN4(n33318), .Q(n17666) );
  OR2X1 U36777 ( .IN1(n33326), .IN2(n34202), .Q(n33321) );
  NAND4X0 U36778 ( .IN1(\s13/msel/gnt_p1 [1]), .IN2(n33347), .IN3(n33349), 
        .IN4(n33321), .QN(n33325) );
  INVX0 U36779 ( .INP(n34203), .ZN(n33327) );
  OR2X1 U36780 ( .IN1(n33327), .IN2(n33326), .Q(n33323) );
  NAND2X0 U36781 ( .IN1(n34203), .IN2(n33322), .QN(n33331) );
  NAND3X0 U36782 ( .IN1(n34411), .IN2(n33323), .IN3(n33331), .QN(n33324) );
  NAND3X0 U36783 ( .IN1(n33351), .IN2(n33325), .IN3(n33324), .QN(n33333) );
  NOR2X0 U36784 ( .IN1(\s13/msel/gnt_p1 [1]), .IN2(n33326), .QN(n33329) );
  NAND2X0 U36785 ( .IN1(n34202), .IN2(n33327), .QN(n33328) );
  NAND2X0 U36786 ( .IN1(n33329), .IN2(n33328), .QN(n33330) );
  OA221X1 U36787 ( .IN1(n33372), .IN2(n34202), .IN3(n33372), .IN4(n33331), 
        .IN5(n33330), .Q(n33332) );
  MUX21X1 U36788 ( .IN1(n33333), .IN2(n33332), .S(\s13/msel/gnt_p1 [2]), .Q(
        n33341) );
  AO21X1 U36789 ( .IN1(n33335), .IN2(n33341), .IN3(n33334), .Q(n33340) );
  NAND2X0 U36790 ( .IN1(n33365), .IN2(n34248), .QN(n33336) );
  NAND3X0 U36791 ( .IN1(n33336), .IN2(n33341), .IN3(n33347), .QN(n33338) );
  NAND3X0 U36792 ( .IN1(\s13/msel/gnt_p1 [1]), .IN2(n33361), .IN3(n34248), 
        .QN(n33337) );
  NAND3X0 U36793 ( .IN1(\s13/msel/gnt_p1 [2]), .IN2(n33338), .IN3(n33337), 
        .QN(n33339) );
  AO22X1 U36794 ( .IN1(\s13/msel/gnt_p1 [1]), .IN2(n33341), .IN3(n33340), 
        .IN4(n33339), .Q(n17665) );
  INVX0 U36795 ( .INP(n33347), .ZN(n33342) );
  NAND2X0 U36796 ( .IN1(n33342), .IN2(n33349), .QN(n33343) );
  NAND2X0 U36797 ( .IN1(n33351), .IN2(n33343), .QN(n33356) );
  AO21X1 U36798 ( .IN1(n33348), .IN2(n33356), .IN3(n33344), .Q(n33363) );
  NAND3X0 U36799 ( .IN1(\s13/msel/gnt_p1 [1]), .IN2(n33363), .IN3(n33374), 
        .QN(n33355) );
  OA21X1 U36800 ( .IN1(n33357), .IN2(n33346), .IN3(n33345), .Q(n33358) );
  OA21X1 U36801 ( .IN1(n33361), .IN2(n33358), .IN3(n33347), .Q(n33364) );
  NAND2X0 U36802 ( .IN1(n33374), .IN2(n33348), .QN(n33352) );
  NAND2X0 U36803 ( .IN1(\s13/msel/gnt_p1 [0]), .IN2(n33349), .QN(n33350) );
  OA221X1 U36804 ( .IN1(n33352), .IN2(n33351), .IN3(n33352), .IN4(n33350), 
        .IN5(n33358), .Q(n33353) );
  OA22X1 U36805 ( .IN1(\s13/msel/gnt_p1 [1]), .IN2(n33364), .IN3(n33361), 
        .IN4(n33353), .Q(n33354) );
  NAND3X0 U36806 ( .IN1(\s13/msel/gnt_p1 [2]), .IN2(n33355), .IN3(n33354), 
        .QN(n33370) );
  INVX0 U36807 ( .INP(n33356), .ZN(n33362) );
  AO221X1 U36808 ( .IN1(n33358), .IN2(n33357), .IN3(n33358), .IN4(n34248), 
        .IN5(n33365), .Q(n33360) );
  AO221X1 U36809 ( .IN1(n33362), .IN2(n33361), .IN3(n33362), .IN4(n33360), 
        .IN5(n33359), .Q(n33368) );
  NAND2X0 U36810 ( .IN1(n34411), .IN2(n33363), .QN(n33367) );
  OR4X1 U36811 ( .IN1(n34411), .IN2(n34248), .IN3(n33365), .IN4(n33364), .Q(
        n33366) );
  NAND4X0 U36812 ( .IN1(n34471), .IN2(n33368), .IN3(n33367), .IN4(n33366), 
        .QN(n33369) );
  NAND2X0 U36813 ( .IN1(n33370), .IN2(n33369), .QN(n33376) );
  AO221X1 U36814 ( .IN1(n34248), .IN2(n34471), .IN3(n34248), .IN4(n33371), 
        .IN5(n33376), .Q(n33382) );
  NAND4X0 U36815 ( .IN1(\s13/msel/gnt_p1 [2]), .IN2(\s13/msel/gnt_p1 [0]), 
        .IN3(n33373), .IN4(n33372), .QN(n33381) );
  NOR2X0 U36816 ( .IN1(\s13/msel/gnt_p1 [1]), .IN2(n33374), .QN(n33375) );
  NOR2X0 U36817 ( .IN1(n33375), .IN2(\s13/msel/gnt_p1 [2]), .QN(n33379) );
  NAND2X0 U36818 ( .IN1(n33377), .IN2(n33376), .QN(n33378) );
  NAND2X0 U36819 ( .IN1(n33379), .IN2(n33378), .QN(n33380) );
  NAND3X0 U36820 ( .IN1(n33382), .IN2(n33381), .IN3(n33380), .QN(n17664) );
  NAND2X0 U36821 ( .IN1(n33383), .IN2(n33385), .QN(n33425) );
  OR2X1 U36822 ( .IN1(n33384), .IN2(n33425), .Q(n33390) );
  NAND2X0 U36823 ( .IN1(n33386), .IN2(n33385), .QN(n33420) );
  AND2X1 U36824 ( .IN1(n33387), .IN2(n33420), .Q(n33422) );
  NOR2X0 U36825 ( .IN1(n33388), .IN2(n33395), .QN(n33427) );
  NOR2X0 U36826 ( .IN1(n33392), .IN2(n33409), .QN(n33416) );
  AO222X1 U36827 ( .IN1(n33390), .IN2(n33422), .IN3(n34653), .IN4(n33389), 
        .IN5(n33427), .IN6(n33416), .Q(n33391) );
  NAND2X0 U36828 ( .IN1(\s13/msel/gnt_p0 [2]), .IN2(n33391), .QN(n33407) );
  NAND2X0 U36829 ( .IN1(n33408), .IN2(n33392), .QN(n33394) );
  NAND3X0 U36830 ( .IN1(n33394), .IN2(n33393), .IN3(n34292), .QN(n33434) );
  INVX0 U36831 ( .INP(n33416), .ZN(n33426) );
  OR2X1 U36832 ( .IN1(n33424), .IN2(n33395), .Q(n33413) );
  OAI22X1 U36833 ( .IN1(n33409), .IN2(n33396), .IN3(n33426), .IN4(n33413), 
        .QN(n33399) );
  OA21X1 U36834 ( .IN1(\s13/msel/gnt_p0 [0]), .IN2(n33398), .IN3(n33397), .Q(
        n33435) );
  OAI22X1 U36835 ( .IN1(n33400), .IN2(n33399), .IN3(\s13/msel/gnt_p0 [1]), 
        .IN4(n33435), .QN(n33401) );
  NOR2X0 U36836 ( .IN1(n33434), .IN2(n33401), .QN(n33404) );
  INVX0 U36837 ( .INP(n33425), .ZN(n33402) );
  NOR2X0 U36838 ( .IN1(n33438), .IN2(n33439), .QN(n33421) );
  NAND2X0 U36839 ( .IN1(n33402), .IN2(n33421), .QN(n33403) );
  NAND2X0 U36840 ( .IN1(n33404), .IN2(n33403), .QN(n33405) );
  NAND3X0 U36841 ( .IN1(n33407), .IN2(n33406), .IN3(n33405), .QN(n17663) );
  NAND2X0 U36842 ( .IN1(n33409), .IN2(n33408), .QN(n33419) );
  OR2X1 U36843 ( .IN1(n33425), .IN2(n33427), .Q(n33410) );
  NAND4X0 U36844 ( .IN1(\s13/msel/gnt_p0 [1]), .IN2(n33412), .IN3(n33411), 
        .IN4(n33410), .QN(n33418) );
  NAND2X0 U36845 ( .IN1(n33421), .IN2(n33425), .QN(n33415) );
  AO22X1 U36846 ( .IN1(n33416), .IN2(n33415), .IN3(n33414), .IN4(n33413), .Q(
        n33417) );
  NAND3X0 U36847 ( .IN1(n33419), .IN2(n33418), .IN3(n33417), .QN(n33433) );
  OA221X1 U36848 ( .IN1(n33426), .IN2(n33421), .IN3(n33426), .IN4(n33420), 
        .IN5(n33427), .Q(n33423) );
  NOR2X0 U36849 ( .IN1(n33423), .IN2(n33422), .QN(n33432) );
  NOR2X0 U36850 ( .IN1(n33425), .IN2(n33424), .QN(n33429) );
  NAND2X0 U36851 ( .IN1(n33427), .IN2(n33426), .QN(n33428) );
  NAND2X0 U36852 ( .IN1(n33429), .IN2(n33428), .QN(n33430) );
  NAND2X0 U36853 ( .IN1(n33430), .IN2(\s13/msel/gnt_p0 [2]), .QN(n33431) );
  NOR2X0 U36854 ( .IN1(n33432), .IN2(n33431), .QN(n33436) );
  AO21X1 U36855 ( .IN1(n34292), .IN2(n33433), .IN3(n33436), .Q(n33447) );
  AO21X1 U36856 ( .IN1(n33435), .IN2(n33447), .IN3(n33434), .Q(n33446) );
  INVX0 U36857 ( .INP(n33436), .ZN(n33437) );
  NOR2X0 U36858 ( .IN1(n33438), .IN2(n33437), .QN(n33441) );
  NAND2X0 U36859 ( .IN1(n34653), .IN2(n33439), .QN(n33440) );
  NAND2X0 U36860 ( .IN1(n33441), .IN2(n33440), .QN(n33444) );
  NAND3X0 U36861 ( .IN1(\s13/msel/gnt_p0 [1]), .IN2(n33442), .IN3(n34653), 
        .QN(n33443) );
  NAND3X0 U36862 ( .IN1(\s13/msel/gnt_p0 [2]), .IN2(n33444), .IN3(n33443), 
        .QN(n33445) );
  AO22X1 U36863 ( .IN1(\s13/msel/gnt_p0 [1]), .IN2(n33447), .IN3(n33446), 
        .IN4(n33445), .Q(n17662) );
  NOR2X0 U36864 ( .IN1(\s13/msel/gnt_p2 [0]), .IN2(n34234), .QN(n33508) );
  INVX0 U36865 ( .INP(n33508), .ZN(n33450) );
  NOR2X0 U36866 ( .IN1(n34480), .IN2(n33448), .QN(n33501) );
  INVX0 U36867 ( .INP(n33501), .ZN(n33514) );
  NOR2X0 U36868 ( .IN1(n34546), .IN2(n33449), .QN(n33515) );
  NAND2X0 U36869 ( .IN1(\s13/msel/gnt_p2 [0]), .IN2(\s13/msel/gnt_p2 [1]), 
        .QN(n33499) );
  INVX0 U36870 ( .INP(n33499), .ZN(n33459) );
  NAND2X0 U36871 ( .IN1(n33515), .IN2(n33459), .QN(n33526) );
  OA21X1 U36872 ( .IN1(n33450), .IN2(n33514), .IN3(n33526), .Q(n33479) );
  NAND3X0 U36873 ( .IN1(n13910), .IN2(m0s13_cyc), .IN3(n34542), .QN(n33513) );
  INVX0 U36874 ( .INP(n33513), .ZN(n33525) );
  NAND3X0 U36875 ( .IN1(n13848), .IN2(m1s13_cyc), .IN3(n34510), .QN(n33491) );
  INVX0 U36876 ( .INP(n33491), .ZN(n33523) );
  MUX21X1 U36877 ( .IN1(n33525), .IN2(n33523), .S(\s13/msel/gnt_p2 [0]), .Q(
        n33480) );
  NAND2X0 U36878 ( .IN1(n34234), .IN2(n33480), .QN(n33453) );
  NAND3X0 U36879 ( .IN1(n13692), .IN2(m4s13_cyc), .IN3(n34543), .QN(n33503) );
  INVX0 U36880 ( .INP(n33503), .ZN(n33487) );
  NOR2X0 U36881 ( .IN1(n34476), .IN2(n33451), .QN(n33478) );
  NOR2X0 U36882 ( .IN1(n33487), .IN2(n33478), .QN(n33462) );
  NAND3X0 U36883 ( .IN1(n13536), .IN2(m7s13_cyc), .IN3(n34586), .QN(n33530) );
  NAND3X0 U36884 ( .IN1(n13588), .IN2(m6s13_cyc), .IN3(n34511), .QN(n33512) );
  NAND2X0 U36885 ( .IN1(n33530), .IN2(n33512), .QN(n33461) );
  INVX0 U36886 ( .INP(n33461), .ZN(n33452) );
  NAND2X0 U36887 ( .IN1(n33462), .IN2(n33452), .QN(n34199) );
  AND4X1 U36888 ( .IN1(n33479), .IN2(n34608), .IN3(n33453), .IN4(n34199), .Q(
        n33460) );
  NOR2X0 U36889 ( .IN1(n33501), .IN2(n33515), .QN(n33468) );
  AND2X1 U36890 ( .IN1(n34234), .IN2(n33491), .Q(n33466) );
  INVX0 U36891 ( .INP(n33515), .ZN(n33486) );
  AO22X1 U36892 ( .IN1(n33468), .IN2(n33466), .IN3(n33508), .IN4(n33486), .Q(
        n33458) );
  NAND2X0 U36893 ( .IN1(\s13/msel/gnt_p2 [1]), .IN2(n33530), .QN(n33455) );
  NOR2X0 U36894 ( .IN1(n33523), .IN2(n33525), .QN(n33470) );
  NAND2X0 U36895 ( .IN1(n33468), .IN2(n33470), .QN(n34200) );
  INVX0 U36896 ( .INP(n34200), .ZN(n33454) );
  AO221X1 U36897 ( .IN1(n33455), .IN2(n33478), .IN3(n33455), .IN4(n33461), 
        .IN5(n33454), .Q(n33456) );
  INVX0 U36898 ( .INP(n33512), .ZN(n33494) );
  MUX21X1 U36899 ( .IN1(n33487), .IN2(n33494), .S(\s13/msel/gnt_p2 [1]), .Q(
        n33532) );
  OA221X1 U36900 ( .IN1(n33456), .IN2(n34288), .IN3(n33456), .IN4(n33532), 
        .IN5(\s13/msel/gnt_p2 [2]), .Q(n33457) );
  AO221X1 U36901 ( .IN1(n33460), .IN2(n33459), .IN3(n33460), .IN4(n33458), 
        .IN5(n33457), .Q(n17660) );
  NAND2X0 U36902 ( .IN1(\s13/msel/gnt_p2 [2]), .IN2(n34288), .QN(n33485) );
  NAND2X0 U36903 ( .IN1(n33462), .IN2(n33461), .QN(n33463) );
  NAND2X0 U36904 ( .IN1(n33468), .IN2(n33463), .QN(n33465) );
  INVX0 U36905 ( .INP(n33478), .ZN(n33529) );
  OA21X1 U36906 ( .IN1(n33470), .IN2(n33461), .IN3(n33529), .Q(n33471) );
  NOR2X0 U36907 ( .IN1(n33487), .IN2(n33499), .QN(n33496) );
  NAND2X0 U36908 ( .IN1(n33470), .IN2(n33462), .QN(n33467) );
  NAND3X0 U36909 ( .IN1(n33486), .IN2(n33467), .IN3(n33463), .QN(n33464) );
  AOI222X1 U36910 ( .IN1(n33466), .IN2(n33465), .IN3(n33471), .IN4(n33496), 
        .IN5(n33464), .IN6(n33508), .QN(n33476) );
  NOR2X0 U36911 ( .IN1(n33494), .IN2(\s13/msel/gnt_p2 [1]), .QN(n33509) );
  OA221X1 U36912 ( .IN1(n33509), .IN2(\s13/msel/gnt_p2 [1]), .IN3(n33509), 
        .IN4(n33467), .IN5(n33530), .Q(n33474) );
  INVX0 U36913 ( .INP(n33468), .ZN(n33469) );
  NAND2X0 U36914 ( .IN1(n33470), .IN2(n33469), .QN(n33473) );
  NAND2X0 U36915 ( .IN1(n34288), .IN2(n34234), .QN(n33497) );
  NOR2X0 U36916 ( .IN1(n33471), .IN2(n33497), .QN(n33472) );
  AO22X1 U36917 ( .IN1(n33474), .IN2(n33473), .IN3(n33478), .IN4(n33472), .Q(
        n33475) );
  MUX21X1 U36918 ( .IN1(n33476), .IN2(n33475), .S(\s13/msel/gnt_p2 [2]), .Q(
        n33483) );
  NAND2X0 U36919 ( .IN1(\s13/msel/gnt_p2 [1]), .IN2(n33494), .QN(n33477) );
  OA21X1 U36920 ( .IN1(n33487), .IN2(n33483), .IN3(n33477), .Q(n33484) );
  NAND2X0 U36921 ( .IN1(\s13/msel/gnt_p2 [0]), .IN2(\s13/msel/gnt_p2 [2]), 
        .QN(n33528) );
  OA21X1 U36922 ( .IN1(n33478), .IN2(n33528), .IN3(n34234), .Q(n33482) );
  OA21X1 U36923 ( .IN1(n33483), .IN2(n33480), .IN3(n33479), .Q(n33481) );
  OAI222X1 U36924 ( .IN1(n33485), .IN2(n33484), .IN3(n33483), .IN4(n33482), 
        .IN5(n33481), .IN6(\s13/msel/gnt_p2 [2]), .QN(n17659) );
  NAND2X0 U36925 ( .IN1(n33503), .IN2(n33512), .QN(n33489) );
  OA21X1 U36926 ( .IN1(n33487), .IN2(n33529), .IN3(n33486), .Q(n33488) );
  OA21X1 U36927 ( .IN1(n34288), .IN2(n33489), .IN3(n33488), .Q(n33492) );
  INVX0 U36928 ( .INP(n33488), .ZN(n33504) );
  NOR2X0 U36929 ( .IN1(n33513), .IN2(n33504), .QN(n33490) );
  OA21X1 U36930 ( .IN1(n33525), .IN2(n33491), .IN3(n33530), .Q(n33505) );
  OA22X1 U36931 ( .IN1(n33492), .IN2(n33490), .IN3(n33505), .IN4(n33489), .Q(
        n33493) );
  OA21X1 U36932 ( .IN1(n33501), .IN2(n33492), .IN3(n33491), .Q(n33500) );
  OA22X1 U36933 ( .IN1(n33501), .IN2(n33493), .IN3(n33500), .IN4(n33497), .Q(
        n33522) );
  OA21X1 U36934 ( .IN1(n33494), .IN2(n33505), .IN3(n33529), .Q(n33498) );
  INVX0 U36935 ( .INP(n33498), .ZN(n33495) );
  NAND2X0 U36936 ( .IN1(n33496), .IN2(n33495), .QN(n33521) );
  NOR2X0 U36937 ( .IN1(n33498), .IN2(n33497), .QN(n33519) );
  NOR3X0 U36938 ( .IN1(n33500), .IN2(n33499), .IN3(n33525), .QN(n33511) );
  NOR2X0 U36939 ( .IN1(n33501), .IN2(n33525), .QN(n33502) );
  OA221X1 U36940 ( .IN1(n33504), .IN2(\s13/msel/gnt_p2 [0]), .IN3(n33504), 
        .IN4(n33503), .IN5(n33502), .Q(n33507) );
  INVX0 U36941 ( .INP(n33505), .ZN(n33506) );
  OA22X1 U36942 ( .IN1(n33509), .IN2(n33508), .IN3(n33507), .IN4(n33506), .Q(
        n33510) );
  NOR2X0 U36943 ( .IN1(n33511), .IN2(n33510), .QN(n33517) );
  NAND4X0 U36944 ( .IN1(n33515), .IN2(n33514), .IN3(n33513), .IN4(n33512), 
        .QN(n33516) );
  NAND2X0 U36945 ( .IN1(n33517), .IN2(n33516), .QN(n33518) );
  NOR2X0 U36946 ( .IN1(n33519), .IN2(n33518), .QN(n33520) );
  OA222X1 U36947 ( .IN1(\s13/msel/gnt_p2 [2]), .IN2(n33522), .IN3(
        \s13/msel/gnt_p2 [2]), .IN4(n33521), .IN5(n33520), .IN6(n34608), .Q(
        n33531) );
  NAND2X0 U36948 ( .IN1(\s13/msel/gnt_p2 [0]), .IN2(n33523), .QN(n33524) );
  OA222X1 U36949 ( .IN1(n33531), .IN2(n33525), .IN3(n33531), .IN4(n34234), 
        .IN5(\s13/msel/gnt_p2 [1]), .IN6(n33524), .Q(n33527) );
  AO21X1 U36950 ( .IN1(n33527), .IN2(n33526), .IN3(\s13/msel/gnt_p2 [2]), .Q(
        n33535) );
  AO221X1 U36951 ( .IN1(\s13/msel/gnt_p2 [1]), .IN2(n33530), .IN3(n34234), 
        .IN4(n33529), .IN5(n33528), .Q(n33534) );
  AO221X1 U36952 ( .IN1(n34288), .IN2(n34608), .IN3(n34288), .IN4(n33532), 
        .IN5(n33531), .Q(n33533) );
  NAND3X0 U36953 ( .IN1(n33535), .IN2(n33534), .IN3(n33533), .QN(n17658) );
  NOR2X0 U36954 ( .IN1(n33536), .IN2(n34379), .QN(n33537) );
  MUX21X1 U36955 ( .IN1(n34367), .IN2(s15_data_o[0]), .S(n33537), .Q(n17657)
         );
  MUX21X1 U36956 ( .IN1(n34604), .IN2(s15_data_o[1]), .S(n33537), .Q(n17656)
         );
  MUX21X1 U36957 ( .IN1(n34334), .IN2(s15_data_o[2]), .S(n33537), .Q(n17655)
         );
  MUX21X1 U36958 ( .IN1(n34512), .IN2(s15_data_o[3]), .S(n33537), .Q(n17654)
         );
  MUX21X1 U36959 ( .IN1(n34477), .IN2(s15_data_o[4]), .S(n33537), .Q(n17653)
         );
  MUX21X1 U36960 ( .IN1(n34646), .IN2(s15_data_o[5]), .S(n33537), .Q(n17652)
         );
  MUX21X1 U36961 ( .IN1(n34481), .IN2(s15_data_o[6]), .S(n33537), .Q(n17651)
         );
  MUX21X1 U36962 ( .IN1(n34648), .IN2(s15_data_o[7]), .S(n33537), .Q(n17650)
         );
  MUX21X1 U36963 ( .IN1(n34635), .IN2(s15_data_o[8]), .S(n33537), .Q(n17649)
         );
  MUX21X1 U36964 ( .IN1(n34571), .IN2(s15_data_o[9]), .S(n33537), .Q(n17648)
         );
  MUX21X1 U36965 ( .IN1(n34547), .IN2(s15_data_o[10]), .S(n33537), .Q(n17647)
         );
  MUX21X1 U36966 ( .IN1(n34652), .IN2(s15_data_o[11]), .S(n33537), .Q(n17646)
         );
  MUX21X1 U36967 ( .IN1(n34357), .IN2(s15_data_o[12]), .S(n33537), .Q(n17645)
         );
  MUX21X1 U36968 ( .IN1(n34544), .IN2(s15_data_o[13]), .S(n33537), .Q(n17644)
         );
  MUX21X1 U36969 ( .IN1(n34358), .IN2(s15_data_o[14]), .S(n33537), .Q(n17643)
         );
  MUX21X1 U36970 ( .IN1(n34513), .IN2(s15_data_o[15]), .S(n33537), .Q(n17642)
         );
  INVX0 U36971 ( .INP(n33564), .ZN(n33574) );
  OA21X1 U36972 ( .IN1(\s14/msel/gnt_p3 [1]), .IN2(n33574), .IN3(n33538), .Q(
        n33606) );
  NOR2X0 U36973 ( .IN1(n34468), .IN2(n34281), .QN(n33542) );
  INVX0 U36974 ( .INP(n33589), .ZN(n33583) );
  NOR2X0 U36975 ( .IN1(n33583), .IN2(\s14/msel/gnt_p3 [1]), .QN(n33541) );
  NAND2X0 U36976 ( .IN1(n33539), .IN2(\s14/msel/gnt_p3 [2]), .QN(n33540) );
  NOR2X0 U36977 ( .IN1(n33541), .IN2(n33540), .QN(n33609) );
  OA22X1 U36978 ( .IN1(\s14/msel/gnt_p3 [1]), .IN2(n33543), .IN3(n33542), 
        .IN4(n33609), .Q(n33544) );
  NAND2X0 U36979 ( .IN1(n33606), .IN2(n33544), .QN(n33553) );
  AND2X1 U36980 ( .IN1(n33595), .IN2(n33554), .Q(n33585) );
  OA21X1 U36981 ( .IN1(n33579), .IN2(n33585), .IN3(n33573), .Q(n33547) );
  NOR2X0 U36982 ( .IN1(n33560), .IN2(n33545), .QN(n33546) );
  NOR3X0 U36983 ( .IN1(n33572), .IN2(n33547), .IN3(n33546), .QN(n33551) );
  INVX0 U36984 ( .INP(n33579), .ZN(n33549) );
  OA222X1 U36985 ( .IN1(n33549), .IN2(n33601), .IN3(n33548), .IN4(
        \s14/msel/gnt_p3 [1]), .IN5(n33587), .IN6(n33566), .Q(n33550) );
  NOR3X0 U36986 ( .IN1(n34211), .IN2(n33551), .IN3(n33550), .QN(n33552) );
  OA22X1 U36987 ( .IN1(n34210), .IN2(n33553), .IN3(\s14/msel/gnt_p3 [2]), 
        .IN4(n33552), .Q(n17641) );
  NAND2X0 U36988 ( .IN1(n33560), .IN2(n33554), .QN(n33604) );
  NAND2X0 U36989 ( .IN1(n33577), .IN2(n33595), .QN(n33562) );
  AO221X1 U36990 ( .IN1(n33573), .IN2(n33555), .IN3(n33573), .IN4(n33589), 
        .IN5(n33562), .Q(n33558) );
  OA21X1 U36991 ( .IN1(n33600), .IN2(n33557), .IN3(n33556), .Q(n33561) );
  NAND2X0 U36992 ( .IN1(\s14/msel/gnt_p3 [0]), .IN2(n33584), .QN(n33559) );
  AO22X1 U36993 ( .IN1(n33558), .IN2(n33561), .IN3(n34447), .IN4(n33559), .Q(
        n33571) );
  OAI221X1 U36994 ( .IN1(n33589), .IN2(n33574), .IN3(n33589), .IN4(n33559), 
        .IN5(n33573), .QN(n33575) );
  AO21X1 U36995 ( .IN1(n33575), .IN2(n33595), .IN3(n33560), .Q(n33596) );
  NAND2X0 U36996 ( .IN1(n33577), .IN2(n33596), .QN(n33570) );
  INVX0 U36997 ( .INP(n33561), .ZN(n33580) );
  INVX0 U36998 ( .INP(n33562), .ZN(n33565) );
  OA221X1 U36999 ( .IN1(n33580), .IN2(\s14/msel/gnt_p3 [0]), .IN3(n33580), 
        .IN4(n33565), .IN5(n33584), .Q(n33563) );
  NOR2X0 U37000 ( .IN1(n33564), .IN2(n33563), .QN(n33588) );
  NAND2X0 U37001 ( .IN1(n33566), .IN2(n33565), .QN(n33568) );
  AO221X1 U37002 ( .IN1(n33588), .IN2(n33578), .IN3(n33588), .IN4(n33568), 
        .IN5(n33567), .Q(n33569) );
  OA221X1 U37003 ( .IN1(n33572), .IN2(n33571), .IN3(n33587), .IN4(n33570), 
        .IN5(n33569), .Q(n33599) );
  NAND2X0 U37004 ( .IN1(n33574), .IN2(n33573), .QN(n33576) );
  OA21X1 U37005 ( .IN1(n33577), .IN2(n33576), .IN3(n33575), .Q(n33586) );
  NOR2X0 U37006 ( .IN1(n33578), .IN2(n33589), .QN(n33581) );
  OA221X1 U37007 ( .IN1(n33586), .IN2(n33581), .IN3(n33586), .IN4(n33580), 
        .IN5(n33579), .Q(n33592) );
  AND3X1 U37008 ( .IN1(n33584), .IN2(n33583), .IN3(n33582), .Q(n33594) );
  OA21X1 U37009 ( .IN1(n33594), .IN2(n33586), .IN3(n33585), .Q(n33591) );
  NOR3X0 U37010 ( .IN1(n33589), .IN2(n33588), .IN3(n33587), .QN(n33590) );
  NOR4X0 U37011 ( .IN1(\s14/msel/gnt_p3 [2]), .IN2(n33592), .IN3(n33591), 
        .IN4(n33590), .QN(n33598) );
  OAI221X1 U37012 ( .IN1(n33596), .IN2(n33595), .IN3(n33596), .IN4(n33594), 
        .IN5(n33593), .QN(n33597) );
  AO22X1 U37013 ( .IN1(\s14/msel/gnt_p3 [2]), .IN2(n33599), .IN3(n33598), 
        .IN4(n33597), .Q(n33605) );
  AO221X1 U37014 ( .IN1(\s14/msel/gnt_p3 [1]), .IN2(n33601), .IN3(n34447), 
        .IN4(n33600), .IN5(n33605), .Q(n33603) );
  NAND3X0 U37015 ( .IN1(n33604), .IN2(n33603), .IN3(n33602), .QN(n33611) );
  INVX0 U37016 ( .INP(n33605), .ZN(n33608) );
  NOR2X0 U37017 ( .IN1(n33606), .IN2(n34281), .QN(n33607) );
  OA22X1 U37018 ( .IN1(\s14/msel/gnt_p3 [0]), .IN2(n33609), .IN3(n33608), 
        .IN4(n33607), .Q(n33610) );
  AO21X1 U37019 ( .IN1(n34281), .IN2(n33611), .IN3(n33610), .Q(n17639) );
  NOR2X0 U37020 ( .IN1(\s14/msel/gnt_p1 [0]), .IN2(n34242), .QN(n33634) );
  NOR2X0 U37021 ( .IN1(n34214), .IN2(n33612), .QN(n33621) );
  NOR2X0 U37022 ( .IN1(n33621), .IN2(n33613), .QN(n33618) );
  INVX0 U37023 ( .INP(n33613), .ZN(n33615) );
  OA21X1 U37024 ( .IN1(n33615), .IN2(n33614), .IN3(n33632), .Q(n33620) );
  OA22X1 U37025 ( .IN1(n33618), .IN2(n33617), .IN3(n33620), .IN4(n33616), .Q(
        n33619) );
  NOR2X0 U37026 ( .IN1(n33619), .IN2(n34386), .QN(n33630) );
  NAND3X0 U37027 ( .IN1(\s14/msel/gnt_p1 [1]), .IN2(n33620), .IN3(n33631), 
        .QN(n33624) );
  INVX0 U37028 ( .INP(n33621), .ZN(n33622) );
  NAND2X0 U37029 ( .IN1(n33622), .IN2(n34242), .QN(n33623) );
  NAND4X0 U37030 ( .IN1(n34386), .IN2(n33625), .IN3(n33624), .IN4(n33623), 
        .QN(n33628) );
  NAND3X0 U37031 ( .IN1(n33626), .IN2(n34215), .IN3(n34242), .QN(n33627) );
  NAND2X0 U37032 ( .IN1(n33628), .IN2(n33627), .QN(n33629) );
  NOR2X0 U37033 ( .IN1(n33630), .IN2(n33629), .QN(n33639) );
  OA21X1 U37034 ( .IN1(\s14/msel/gnt_p1 [0]), .IN2(n33631), .IN3(n33639), .Q(
        n33633) );
  AO22X1 U37035 ( .IN1(n33635), .IN2(n33634), .IN3(n33633), .IN4(n33632), .Q(
        n33642) );
  INVX0 U37036 ( .INP(n33636), .ZN(n33637) );
  AO21X1 U37037 ( .IN1(n33639), .IN2(n33638), .IN3(n33637), .Q(n33641) );
  AND2X1 U37038 ( .IN1(\s14/msel/gnt_p1 [1]), .IN2(n33639), .Q(n33640) );
  AO221X1 U37039 ( .IN1(\s14/msel/gnt_p1 [2]), .IN2(n33642), .IN3(n34386), 
        .IN4(n33641), .IN5(n33640), .Q(n17637) );
  NAND2X0 U37040 ( .IN1(n33659), .IN2(n33668), .QN(n33648) );
  INVX0 U37041 ( .INP(n33643), .ZN(n33645) );
  NOR2X0 U37042 ( .IN1(n33649), .IN2(n33644), .QN(n33651) );
  OR3X1 U37043 ( .IN1(n34247), .IN2(n33645), .IN3(n33651), .Q(n33647) );
  NAND2X0 U37044 ( .IN1(n33645), .IN2(n33654), .QN(n33650) );
  NAND3X0 U37045 ( .IN1(n34247), .IN2(n33650), .IN3(n33672), .QN(n33646) );
  NAND3X0 U37046 ( .IN1(n33648), .IN2(n33647), .IN3(n33646), .QN(n33657) );
  AND2X1 U37047 ( .IN1(n33650), .IN2(n33649), .Q(n33653) );
  NOR2X0 U37048 ( .IN1(n33684), .IN2(n33651), .QN(n33652) );
  AO222X1 U37049 ( .IN1(\s14/msel/gnt_p0 [1]), .IN2(n33667), .IN3(
        \s14/msel/gnt_p0 [1]), .IN4(n33653), .IN5(n33652), .IN6(n34247), .Q(
        n33656) );
  NAND4X0 U37050 ( .IN1(n33654), .IN2(n34247), .IN3(n33686), .IN4(n33676), 
        .QN(n33655) );
  OA221X1 U37051 ( .IN1(\s14/msel/gnt_p0 [2]), .IN2(n33657), .IN3(n34387), 
        .IN4(n33656), .IN5(n33655), .Q(n33666) );
  OA21X1 U37052 ( .IN1(\s14/msel/gnt_p0 [0]), .IN2(n33688), .IN3(n33666), .Q(
        n33658) );
  NOR2X0 U37053 ( .IN1(n33658), .IN2(n34387), .QN(n33662) );
  NAND2X0 U37054 ( .IN1(n33660), .IN2(n33659), .QN(n33661) );
  NAND2X0 U37055 ( .IN1(n33662), .IN2(n33661), .QN(n33665) );
  AO221X1 U37056 ( .IN1(n33666), .IN2(\s14/msel/gnt_p0 [0]), .IN3(n33666), 
        .IN4(n33694), .IN5(n33663), .Q(n33664) );
  AO22X1 U37057 ( .IN1(\s14/msel/gnt_p0 [1]), .IN2(n33666), .IN3(n33665), 
        .IN4(n33664), .Q(n17634) );
  INVX0 U37058 ( .INP(n33694), .ZN(n33675) );
  NOR2X0 U37059 ( .IN1(n33672), .IN2(n33675), .QN(n33677) );
  OR2X1 U37060 ( .IN1(n33667), .IN2(n33677), .Q(n33685) );
  AO21X1 U37061 ( .IN1(n33684), .IN2(n33688), .IN3(n33668), .Q(n33671) );
  OA221X1 U37062 ( .IN1(n33671), .IN2(\s14/msel/gnt_p0 [0]), .IN3(n33671), 
        .IN4(n33688), .IN5(n33669), .Q(n33670) );
  OA221X1 U37063 ( .IN1(n33685), .IN2(n33670), .IN3(n33685), .IN4(n33694), 
        .IN5(n33686), .Q(n33693) );
  INVX0 U37064 ( .INP(n33671), .ZN(n33680) );
  OA21X1 U37065 ( .IN1(n33680), .IN2(n33682), .IN3(n33672), .Q(n33683) );
  NOR3X0 U37066 ( .IN1(n33675), .IN2(n33683), .IN3(n33673), .QN(n33692) );
  NAND2X0 U37067 ( .IN1(n33686), .IN2(n33688), .QN(n33674) );
  AO221X1 U37068 ( .IN1(n33676), .IN2(n33675), .IN3(n33676), .IN4(n34639), 
        .IN5(n33674), .Q(n33679) );
  NAND3X0 U37069 ( .IN1(n33677), .IN2(n33688), .IN3(n33686), .QN(n33678) );
  AND3X1 U37070 ( .IN1(n33680), .IN2(n33679), .IN3(n33678), .Q(n33681) );
  OA22X1 U37071 ( .IN1(\s14/msel/gnt_p0 [1]), .IN2(n33683), .IN3(n33682), 
        .IN4(n33681), .Q(n33690) );
  AO21X1 U37072 ( .IN1(n33686), .IN2(n33685), .IN3(n33684), .Q(n33687) );
  NAND4X0 U37073 ( .IN1(\s14/msel/gnt_p0 [1]), .IN2(\s14/msel/gnt_p0 [0]), 
        .IN3(n33688), .IN4(n33687), .QN(n33689) );
  NAND2X0 U37074 ( .IN1(n33690), .IN2(n33689), .QN(n33691) );
  AO222X1 U37075 ( .IN1(\s14/msel/gnt_p0 [2]), .IN2(n33693), .IN3(
        \s14/msel/gnt_p0 [2]), .IN4(n33692), .IN5(n33691), .IN6(n34387), .Q(
        n33697) );
  OA21X1 U37076 ( .IN1(\s14/msel/gnt_p0 [1]), .IN2(n33694), .IN3(n33697), .Q(
        n33701) );
  NOR2X0 U37077 ( .IN1(n33695), .IN2(n34387), .QN(n33698) );
  OA22X1 U37078 ( .IN1(\s14/msel/gnt_p0 [0]), .IN2(n33698), .IN3(n33697), 
        .IN4(n33696), .Q(n33699) );
  AO221X1 U37079 ( .IN1(n34387), .IN2(n33701), .IN3(n34387), .IN4(n33700), 
        .IN5(n33699), .Q(n17633) );
  MUX21X1 U37080 ( .IN1(n33702), .IN2(n33717), .S(\s14/msel/gnt_p2 [1]), .Q(
        n33758) );
  NAND2X0 U37081 ( .IN1(\s14/msel/gnt_p2 [1]), .IN2(n33756), .QN(n33704) );
  NAND2X0 U37082 ( .IN1(n33707), .IN2(n33755), .QN(n33703) );
  AO22X1 U37083 ( .IN1(n34271), .IN2(n33758), .IN3(n33704), .IN4(n33703), .Q(
        n33715) );
  OAI22X1 U37084 ( .IN1(n33731), .IN2(n34381), .IN3(n33706), .IN4(n33705), 
        .QN(n33712) );
  NAND2X0 U37085 ( .IN1(n33708), .IN2(n33707), .QN(n33711) );
  NAND2X0 U37086 ( .IN1(n34381), .IN2(n33709), .QN(n33710) );
  AND4X1 U37087 ( .IN1(n33713), .IN2(n33712), .IN3(n33711), .IN4(n33710), .Q(
        n33714) );
  AO221X1 U37088 ( .IN1(\s14/msel/gnt_p2 [2]), .IN2(n33716), .IN3(
        \s14/msel/gnt_p2 [2]), .IN4(n33715), .IN5(n33714), .Q(n17632) );
  OA21X1 U37089 ( .IN1(n33751), .IN2(n33719), .IN3(n33756), .Q(n33736) );
  OA21X1 U37090 ( .IN1(n33717), .IN2(n33736), .IN3(n33755), .Q(n33734) );
  NAND2X0 U37091 ( .IN1(n33730), .IN2(n33735), .QN(n33724) );
  AO21X1 U37092 ( .IN1(n33718), .IN2(n33735), .IN3(n33731), .Q(n33722) );
  INVX0 U37093 ( .INP(n33722), .ZN(n33742) );
  OA21X1 U37094 ( .IN1(n34271), .IN2(n33724), .IN3(n33742), .Q(n33720) );
  OA21X1 U37095 ( .IN1(n33729), .IN2(n33720), .IN3(n33719), .Q(n33728) );
  OA22X1 U37096 ( .IN1(n33734), .IN2(n33721), .IN3(n33728), .IN4(n33732), .Q(
        n33727) );
  NOR3X0 U37097 ( .IN1(n33751), .IN2(n33724), .IN3(n34271), .QN(n33723) );
  NOR2X0 U37098 ( .IN1(n33723), .IN2(n33722), .QN(n33725) );
  AO221X1 U37099 ( .IN1(n33725), .IN2(n33736), .IN3(n33725), .IN4(n33724), 
        .IN5(n33729), .Q(n33726) );
  NAND3X0 U37100 ( .IN1(n34460), .IN2(n33727), .IN3(n33726), .QN(n33748) );
  OR3X1 U37101 ( .IN1(n34381), .IN2(n33751), .IN3(n33728), .Q(n33746) );
  NOR2X0 U37102 ( .IN1(n33751), .IN2(n33729), .QN(n33739) );
  NAND3X0 U37103 ( .IN1(n33739), .IN2(n33731), .IN3(n33730), .QN(n33733) );
  AO21X1 U37104 ( .IN1(n33734), .IN2(n33733), .IN3(n33732), .Q(n33745) );
  AND3X1 U37105 ( .IN1(n33735), .IN2(n33739), .IN3(\s14/msel/gnt_p2 [0]), .Q(
        n33738) );
  INVX0 U37106 ( .INP(n33736), .ZN(n33737) );
  NOR2X0 U37107 ( .IN1(n33738), .IN2(n33737), .QN(n33743) );
  INVX0 U37108 ( .INP(n33739), .ZN(n33741) );
  AO221X1 U37109 ( .IN1(n33743), .IN2(n33742), .IN3(n33743), .IN4(n33741), 
        .IN5(n33740), .Q(n33744) );
  NAND4X0 U37110 ( .IN1(\s14/msel/gnt_p2 [2]), .IN2(n33746), .IN3(n33745), 
        .IN4(n33744), .QN(n33747) );
  NAND2X0 U37111 ( .IN1(n33748), .IN2(n33747), .QN(n33757) );
  NAND2X0 U37112 ( .IN1(\s14/msel/gnt_p2 [0]), .IN2(n33749), .QN(n33750) );
  OA222X1 U37113 ( .IN1(n33757), .IN2(n33751), .IN3(n33757), .IN4(n34381), 
        .IN5(\s14/msel/gnt_p2 [1]), .IN6(n33750), .Q(n33753) );
  AO21X1 U37114 ( .IN1(n33753), .IN2(n33752), .IN3(\s14/msel/gnt_p2 [2]), .Q(
        n33761) );
  AO221X1 U37115 ( .IN1(\s14/msel/gnt_p2 [1]), .IN2(n33756), .IN3(n34381), 
        .IN4(n33755), .IN5(n33754), .Q(n33760) );
  AO221X1 U37116 ( .IN1(n34271), .IN2(n34460), .IN3(n34271), .IN4(n33758), 
        .IN5(n33757), .Q(n33759) );
  NAND3X0 U37117 ( .IN1(n33761), .IN2(n33760), .IN3(n33759), .QN(n17630) );
  NOR2X0 U37118 ( .IN1(n33762), .IN2(n34379), .QN(n33763) );
  MUX21X1 U37119 ( .IN1(n34298), .IN2(s15_data_o[0]), .S(n33763), .Q(n17629)
         );
  MUX21X1 U37120 ( .IN1(n34482), .IN2(s15_data_o[1]), .S(n33763), .Q(n17628)
         );
  MUX21X1 U37121 ( .IN1(n34302), .IN2(s15_data_o[2]), .S(n33763), .Q(n17627)
         );
  MUX21X1 U37122 ( .IN1(n34514), .IN2(s15_data_o[3]), .S(n33763), .Q(n17626)
         );
  MUX21X1 U37123 ( .IN1(n34359), .IN2(s15_data_o[4]), .S(n33763), .Q(n17625)
         );
  MUX21X1 U37124 ( .IN1(n34602), .IN2(s15_data_o[5]), .S(n33763), .Q(n17624)
         );
  MUX21X1 U37125 ( .IN1(n34303), .IN2(s15_data_o[6]), .S(n33763), .Q(n17623)
         );
  MUX21X1 U37126 ( .IN1(n34515), .IN2(s15_data_o[7]), .S(n33763), .Q(n17622)
         );
  MUX21X1 U37127 ( .IN1(n34299), .IN2(s15_data_o[8]), .S(n33763), .Q(n17621)
         );
  MUX21X1 U37128 ( .IN1(n34516), .IN2(s15_data_o[9]), .S(n33763), .Q(n17620)
         );
  MUX21X1 U37129 ( .IN1(n34300), .IN2(s15_data_o[10]), .S(n33763), .Q(n17619)
         );
  MUX21X1 U37130 ( .IN1(n34517), .IN2(s15_data_o[11]), .S(n33763), .Q(n17618)
         );
  MUX21X1 U37131 ( .IN1(n34360), .IN2(s15_data_o[12]), .S(n33763), .Q(n17617)
         );
  MUX21X1 U37132 ( .IN1(n34598), .IN2(s15_data_o[13]), .S(n33763), .Q(n17616)
         );
  MUX21X1 U37133 ( .IN1(n34301), .IN2(s15_data_o[14]), .S(n33763), .Q(n17615)
         );
  MUX21X1 U37134 ( .IN1(n34518), .IN2(s15_data_o[15]), .S(n33763), .Q(n17614)
         );
  NAND2X0 U37135 ( .IN1(\s15/msel/gnt_p3 [0]), .IN2(\s15/msel/gnt_p3 [1]), 
        .QN(n33816) );
  INVX0 U37136 ( .INP(n33852), .ZN(n33813) );
  INVX0 U37137 ( .INP(n33833), .ZN(n33854) );
  MUX21X1 U37138 ( .IN1(n33813), .IN2(n33854), .S(\s15/msel/gnt_p3 [0]), .Q(
        n33801) );
  NAND2X0 U37139 ( .IN1(\s15/msel/gnt_p3 [1]), .IN2(n33853), .QN(n33764) );
  OA21X1 U37140 ( .IN1(n33801), .IN2(\s15/msel/gnt_p3 [1]), .IN3(n33764), .Q(
        n33765) );
  NAND2X0 U37141 ( .IN1(n33816), .IN2(n33765), .QN(n33768) );
  NOR2X0 U37142 ( .IN1(\s15/msel/gnt_p3 [1]), .IN2(n34283), .QN(n33777) );
  NOR2X0 U37143 ( .IN1(\s15/msel/gnt_p3 [0]), .IN2(\s15/msel/gnt_p3 [1]), .QN(
        n33791) );
  NAND2X0 U37144 ( .IN1(n33791), .IN2(n33833), .QN(n33788) );
  INVX0 U37145 ( .INP(n33788), .ZN(n33766) );
  AND2X1 U37146 ( .IN1(\s15/msel/gnt_p3 [1]), .IN2(n33803), .Q(n33787) );
  AO221X1 U37147 ( .IN1(n33773), .IN2(n33777), .IN3(n33773), .IN4(n33766), 
        .IN5(n33787), .Q(n33767) );
  AND3X1 U37148 ( .IN1(n33769), .IN2(n33768), .IN3(n33767), .Q(n33772) );
  MUX21X1 U37149 ( .IN1(n33822), .IN2(n33827), .S(\s15/msel/gnt_p3 [1]), .Q(
        n33811) );
  OA22X1 U37150 ( .IN1(\s15/msel/gnt_p3 [0]), .IN2(n33811), .IN3(n33774), 
        .IN4(n33779), .Q(n33770) );
  NAND2X0 U37151 ( .IN1(n33815), .IN2(n34421), .QN(n33842) );
  NAND2X0 U37152 ( .IN1(n33817), .IN2(n34421), .QN(n33850) );
  NAND4X0 U37153 ( .IN1(n33770), .IN2(n33812), .IN3(n33842), .IN4(n33850), 
        .QN(n33771) );
  MUX21X1 U37154 ( .IN1(n33772), .IN2(n33771), .S(\s15/msel/gnt_p3 [2]), .Q(
        n17613) );
  NAND2X0 U37155 ( .IN1(\s15/msel/gnt_p3 [1]), .IN2(n33793), .QN(n33778) );
  NAND2X0 U37156 ( .IN1(n33773), .IN2(n33778), .QN(n33785) );
  NAND2X0 U37157 ( .IN1(n33791), .IN2(n33814), .QN(n33782) );
  INVX0 U37158 ( .INP(n33791), .ZN(n33829) );
  NAND2X0 U37159 ( .IN1(n33829), .IN2(n33774), .QN(n33786) );
  NAND3X0 U37160 ( .IN1(n33782), .IN2(n33816), .IN3(n33786), .QN(n33775) );
  NAND3X0 U37161 ( .IN1(n33776), .IN2(n33785), .IN3(n33775), .QN(n33784) );
  NAND2X0 U37162 ( .IN1(\s15/msel/gnt_p3 [1]), .IN2(n34283), .QN(n33802) );
  INVX0 U37163 ( .INP(n33802), .ZN(n33821) );
  NOR2X0 U37164 ( .IN1(n33821), .IN2(n33777), .QN(n33836) );
  NOR2X0 U37165 ( .IN1(n33779), .IN2(n33778), .QN(n33790) );
  NAND2X0 U37166 ( .IN1(n33812), .IN2(n33842), .QN(n33780) );
  NOR2X0 U37167 ( .IN1(n33790), .IN2(n33780), .QN(n33781) );
  OA22X1 U37168 ( .IN1(n33792), .IN2(n33782), .IN3(n33836), .IN4(n33781), .Q(
        n33783) );
  NAND3X0 U37169 ( .IN1(n33784), .IN2(n33783), .IN3(\s15/msel/gnt_p3 [2]), 
        .QN(n33800) );
  INVX0 U37170 ( .INP(n33785), .ZN(n33789) );
  OA22X1 U37171 ( .IN1(n33789), .IN2(n33788), .IN3(n33787), .IN4(n33786), .Q(
        n33798) );
  INVX0 U37172 ( .INP(n33790), .ZN(n33797) );
  NAND2X0 U37173 ( .IN1(n33791), .IN2(n33854), .QN(n33795) );
  INVX0 U37174 ( .INP(n33792), .ZN(n33794) );
  NAND3X0 U37175 ( .IN1(n33795), .IN2(n33794), .IN3(n33793), .QN(n33796) );
  NAND4X0 U37176 ( .IN1(n33798), .IN2(n34433), .IN3(n33797), .IN4(n33796), 
        .QN(n33799) );
  NAND2X0 U37177 ( .IN1(n33800), .IN2(n33799), .QN(n33805) );
  OR2X1 U37178 ( .IN1(n34421), .IN2(n33805), .Q(n33810) );
  OA22X1 U37179 ( .IN1(n33802), .IN2(n33853), .IN3(n33805), .IN4(n33801), .Q(
        n33804) );
  INVX0 U37180 ( .INP(n33803), .ZN(n33828) );
  INVX0 U37181 ( .INP(n33816), .ZN(n33835) );
  NAND2X0 U37182 ( .IN1(n33828), .IN2(n33835), .QN(n33857) );
  AO21X1 U37183 ( .IN1(n33804), .IN2(n33857), .IN3(\s15/msel/gnt_p3 [2]), .Q(
        n33809) );
  NAND2X0 U37184 ( .IN1(\s15/msel/gnt_p3 [1]), .IN2(n33823), .QN(n33851) );
  OA21X1 U37185 ( .IN1(n33817), .IN2(n33805), .IN3(n33851), .Q(n33807) );
  OA22X1 U37186 ( .IN1(n33818), .IN2(n33805), .IN3(n34421), .IN4(n33827), .Q(
        n33806) );
  AO221X1 U37187 ( .IN1(\s15/msel/gnt_p3 [0]), .IN2(n33807), .IN3(n34283), 
        .IN4(n33806), .IN5(n34433), .Q(n33808) );
  NAND3X0 U37188 ( .IN1(n33810), .IN2(n33809), .IN3(n33808), .QN(n17612) );
  AO21X1 U37189 ( .IN1(\s15/msel/gnt_p3 [2]), .IN2(n33811), .IN3(
        \s15/msel/gnt_p3 [0]), .Q(n33862) );
  OA21X1 U37190 ( .IN1(n33813), .IN2(n33833), .IN3(n33812), .Q(n33820) );
  OA21X1 U37191 ( .IN1(n33815), .IN2(n33820), .IN3(n33814), .Q(n33831) );
  NOR3X0 U37192 ( .IN1(n33818), .IN2(n33831), .IN3(n33816), .QN(n33849) );
  AO21X1 U37193 ( .IN1(n33822), .IN2(n33817), .IN3(n33828), .Q(n33838) );
  NOR2X0 U37194 ( .IN1(n34283), .IN2(n33818), .QN(n33839) );
  OAI221X1 U37195 ( .IN1(n33838), .IN2(n33827), .IN3(n33838), .IN4(n33839), 
        .IN5(n33853), .QN(n33832) );
  NOR2X0 U37196 ( .IN1(n33852), .IN2(n33838), .QN(n33819) );
  AO221X1 U37197 ( .IN1(n33832), .IN2(n33833), .IN3(n33832), .IN4(n33829), 
        .IN5(n33819), .Q(n33826) );
  INVX0 U37198 ( .INP(n33820), .ZN(n33837) );
  NAND4X0 U37199 ( .IN1(n33821), .IN2(n33827), .IN3(n33822), .IN4(n33837), 
        .QN(n33825) );
  NAND4X0 U37200 ( .IN1(n33823), .IN2(n33827), .IN3(n33822), .IN4(n33853), 
        .QN(n33824) );
  NAND4X0 U37201 ( .IN1(n33826), .IN2(n34433), .IN3(n33825), .IN4(n33824), 
        .QN(n33848) );
  NAND4X0 U37202 ( .IN1(n33828), .IN2(n33827), .IN3(n33852), .IN4(n33853), 
        .QN(n33830) );
  AO21X1 U37203 ( .IN1(n33831), .IN2(n33830), .IN3(n33829), .Q(n33846) );
  NAND2X0 U37204 ( .IN1(n33833), .IN2(n33832), .QN(n33834) );
  NAND3X0 U37205 ( .IN1(n33835), .IN2(n33852), .IN3(n33834), .QN(n33845) );
  INVX0 U37206 ( .INP(n33836), .ZN(n33843) );
  AND2X1 U37207 ( .IN1(n33852), .IN2(n33853), .Q(n33840) );
  AO221X1 U37208 ( .IN1(n33840), .IN2(n33839), .IN3(n33840), .IN4(n33838), 
        .IN5(n33837), .Q(n33841) );
  NAND3X0 U37209 ( .IN1(n33843), .IN2(n33842), .IN3(n33841), .QN(n33844) );
  NAND4X0 U37210 ( .IN1(\s15/msel/gnt_p3 [2]), .IN2(n33846), .IN3(n33845), 
        .IN4(n33844), .QN(n33847) );
  OA21X1 U37211 ( .IN1(n33849), .IN2(n33848), .IN3(n33847), .Q(n33861) );
  NAND2X0 U37212 ( .IN1(n33851), .IN2(n33850), .QN(n33860) );
  NOR2X0 U37213 ( .IN1(n34283), .IN2(n34433), .QN(n33859) );
  OAI221X1 U37214 ( .IN1(n34421), .IN2(n33853), .IN3(\s15/msel/gnt_p3 [1]), 
        .IN4(n33852), .IN5(n33861), .QN(n33856) );
  NAND3X0 U37215 ( .IN1(\s15/msel/gnt_p3 [0]), .IN2(n33854), .IN3(n34421), 
        .QN(n33855) );
  NAND3X0 U37216 ( .IN1(n33857), .IN2(n33856), .IN3(n33855), .QN(n33858) );
  AO222X1 U37217 ( .IN1(n33862), .IN2(n33861), .IN3(n33860), .IN4(n33859), 
        .IN5(n33858), .IN6(n34433), .Q(n17611) );
  NOR2X0 U37218 ( .IN1(n33864), .IN2(n33863), .QN(n33865) );
  INVX0 U37219 ( .INP(n33887), .ZN(n33890) );
  OA22X1 U37220 ( .IN1(\s15/msel/gnt_p1 [0]), .IN2(n33865), .IN3(
        \s15/msel/gnt_p1 [1]), .IN4(n33890), .Q(n33867) );
  AO21X1 U37221 ( .IN1(n33867), .IN2(n33866), .IN3(n34448), .Q(n33876) );
  NAND3X0 U37222 ( .IN1(n34272), .IN2(n33868), .IN3(\s15/msel/gnt_p1 [1]), 
        .QN(n33869) );
  NAND2X0 U37223 ( .IN1(n33869), .IN2(n34448), .QN(n33900) );
  INVX0 U37224 ( .INP(n33900), .ZN(n33874) );
  OA21X1 U37225 ( .IN1(\s15/msel/gnt_p1 [0]), .IN2(n33871), .IN3(n33870), .Q(
        n33901) );
  AO21X1 U37226 ( .IN1(n33901), .IN2(n33889), .IN3(\s15/msel/gnt_p1 [1]), .Q(
        n33872) );
  NAND4X0 U37227 ( .IN1(n33874), .IN2(n33888), .IN3(n33873), .IN4(n33872), 
        .QN(n33875) );
  NAND3X0 U37228 ( .IN1(n33877), .IN2(n33876), .IN3(n33875), .QN(n17610) );
  NAND2X0 U37229 ( .IN1(n33890), .IN2(n33878), .QN(n33879) );
  NAND4X0 U37230 ( .IN1(\s15/msel/gnt_p1 [1]), .IN2(n33895), .IN3(n33880), 
        .IN4(n33879), .QN(n33883) );
  NAND3X0 U37231 ( .IN1(n33889), .IN2(n33888), .IN3(n33881), .QN(n33885) );
  NAND2X0 U37232 ( .IN1(n33885), .IN2(n34412), .QN(n33882) );
  NAND3X0 U37233 ( .IN1(n33888), .IN2(n33883), .IN3(n33882), .QN(n33893) );
  AO22X1 U37234 ( .IN1(n33887), .IN2(n33886), .IN3(n33885), .IN4(n33884), .Q(
        n33892) );
  NAND4X0 U37235 ( .IN1(n33890), .IN2(n34412), .IN3(n33889), .IN4(n33888), 
        .QN(n33891) );
  OA221X1 U37236 ( .IN1(\s15/msel/gnt_p1 [2]), .IN2(n33893), .IN3(n34448), 
        .IN4(n33892), .IN5(n33891), .Q(n33904) );
  NAND2X0 U37237 ( .IN1(n33894), .IN2(n34272), .QN(n33896) );
  NAND3X0 U37238 ( .IN1(n33896), .IN2(n33904), .IN3(n33895), .QN(n33899) );
  NAND3X0 U37239 ( .IN1(\s15/msel/gnt_p1 [1]), .IN2(n33897), .IN3(n34272), 
        .QN(n33898) );
  NAND3X0 U37240 ( .IN1(\s15/msel/gnt_p1 [2]), .IN2(n33899), .IN3(n33898), 
        .QN(n33903) );
  AO21X1 U37241 ( .IN1(n33901), .IN2(n33904), .IN3(n33900), .Q(n33902) );
  AO22X1 U37242 ( .IN1(\s15/msel/gnt_p1 [1]), .IN2(n33904), .IN3(n33903), 
        .IN4(n33902), .Q(n17609) );
  NAND3X0 U37243 ( .IN1(m6s15_cyc), .IN2(n13590), .IN3(n13564), .QN(n33964) );
  INVX0 U37244 ( .INP(n33964), .ZN(n33958) );
  NAND3X0 U37245 ( .IN1(m7s15_cyc), .IN2(n13538), .IN3(n13485), .QN(n33949) );
  INVX0 U37246 ( .INP(n33949), .ZN(n33960) );
  NOR2X0 U37247 ( .IN1(n33958), .IN2(n33960), .QN(n33919) );
  NOR2X0 U37248 ( .IN1(\s15/msel/gnt_p0 [1]), .IN2(n33919), .QN(n33918) );
  NAND3X0 U37249 ( .IN1(m5s15_cyc), .IN2(n13642), .IN3(n13616), .QN(n33952) );
  MUX21X1 U37250 ( .IN1(n33952), .IN2(n33949), .S(\s15/msel/gnt_p0 [1]), .Q(
        n33905) );
  INVX0 U37251 ( .INP(n33905), .ZN(n33910) );
  NAND3X0 U37252 ( .IN1(m4s15_cyc), .IN2(n13694), .IN3(n13668), .QN(n33965) );
  INVX0 U37253 ( .INP(n33965), .ZN(n33953) );
  MUX21X1 U37254 ( .IN1(n33953), .IN2(n33958), .S(\s15/msel/gnt_p0 [1]), .Q(
        n33983) );
  OA21X1 U37255 ( .IN1(n33910), .IN2(n33983), .IN3(n34261), .Q(n33906) );
  NOR2X0 U37256 ( .IN1(n33918), .IN2(n33906), .QN(n33908) );
  NAND3X0 U37257 ( .IN1(m2s15_cyc), .IN2(n13798), .IN3(n13772), .QN(n33948) );
  INVX0 U37258 ( .INP(n33948), .ZN(n33974) );
  NAND3X0 U37259 ( .IN1(m3s15_cyc), .IN2(n13746), .IN3(n13720), .QN(n33951) );
  INVX0 U37260 ( .INP(n33951), .ZN(n33933) );
  NOR2X0 U37261 ( .IN1(n33974), .IN2(n33933), .QN(n33921) );
  NAND3X0 U37262 ( .IN1(m0s15_cyc), .IN2(n13914), .IN3(n13876), .QN(n33962) );
  INVX0 U37263 ( .INP(n33962), .ZN(n33979) );
  NAND3X0 U37264 ( .IN1(m1s15_cyc), .IN2(n13850), .IN3(n13824), .QN(n33959) );
  INVX0 U37265 ( .INP(n33959), .ZN(n33961) );
  NOR2X0 U37266 ( .IN1(n33979), .IN2(n33961), .QN(n33925) );
  NAND2X0 U37267 ( .IN1(n33921), .IN2(n33925), .QN(n33907) );
  NAND2X0 U37268 ( .IN1(n33908), .IN2(n33907), .QN(n33909) );
  NAND2X0 U37269 ( .IN1(\s15/msel/gnt_p0 [2]), .IN2(n33909), .QN(n33917) );
  NAND3X0 U37270 ( .IN1(\s15/msel/gnt_p0 [0]), .IN2(\s15/msel/gnt_p0 [2]), 
        .IN3(n33910), .QN(n33984) );
  INVX0 U37271 ( .INP(n33919), .ZN(n33924) );
  NAND2X0 U37272 ( .IN1(n33952), .IN2(n33965), .QN(n33920) );
  NOR2X0 U37273 ( .IN1(n33924), .IN2(n33920), .QN(n33915) );
  NOR2X0 U37274 ( .IN1(n34261), .IN2(n34226), .QN(n33966) );
  AND2X1 U37275 ( .IN1(n34226), .IN2(n33959), .Q(n33929) );
  NOR2X0 U37276 ( .IN1(\s15/msel/gnt_p0 [0]), .IN2(n34226), .QN(n33932) );
  AO22X1 U37277 ( .IN1(n33921), .IN2(n33929), .IN3(n33932), .IN4(n33951), .Q(
        n33911) );
  NOR2X0 U37278 ( .IN1(n33966), .IN2(n33911), .QN(n33914) );
  NAND2X0 U37279 ( .IN1(\s15/msel/gnt_p0 [0]), .IN2(n33961), .QN(n33978) );
  OA21X1 U37280 ( .IN1(\s15/msel/gnt_p0 [0]), .IN2(n33962), .IN3(n33978), .Q(
        n33941) );
  NOR2X0 U37281 ( .IN1(\s15/msel/gnt_p0 [1]), .IN2(n33941), .QN(n33913) );
  NAND2X0 U37282 ( .IN1(n33932), .IN2(n33974), .QN(n33912) );
  NAND2X0 U37283 ( .IN1(n33933), .IN2(n33966), .QN(n33980) );
  NAND3X0 U37284 ( .IN1(n33912), .IN2(n33980), .IN3(n34441), .QN(n33940) );
  OR4X1 U37285 ( .IN1(n33915), .IN2(n33914), .IN3(n33913), .IN4(n33940), .Q(
        n33916) );
  NAND3X0 U37286 ( .IN1(n33917), .IN2(n33984), .IN3(n33916), .QN(n17607) );
  OA22X1 U37287 ( .IN1(n33960), .IN2(n34226), .IN3(n33918), .IN4(n34261), .Q(
        n33928) );
  NAND2X0 U37288 ( .IN1(n33919), .IN2(n33921), .QN(n33931) );
  NOR2X0 U37289 ( .IN1(n33931), .IN2(\s15/msel/gnt_p0 [1]), .QN(n33923) );
  NAND2X0 U37290 ( .IN1(n33921), .IN2(n33920), .QN(n33930) );
  NAND2X0 U37291 ( .IN1(n33930), .IN2(n33925), .QN(n33922) );
  NOR2X0 U37292 ( .IN1(n33923), .IN2(n33922), .QN(n33927) );
  OR2X1 U37293 ( .IN1(n33925), .IN2(n33924), .Q(n33934) );
  AND2X1 U37294 ( .IN1(n33931), .IN2(n33934), .Q(n33926) );
  NAND2X0 U37295 ( .IN1(n34261), .IN2(n34226), .QN(n33967) );
  OA22X1 U37296 ( .IN1(n33928), .IN2(n33927), .IN3(n33926), .IN4(n33967), .Q(
        n33939) );
  NAND3X0 U37297 ( .IN1(n33931), .IN2(n33930), .IN3(n33929), .QN(n33937) );
  NAND2X0 U37298 ( .IN1(n33933), .IN2(n33932), .QN(n33936) );
  NAND4X0 U37299 ( .IN1(\s15/msel/gnt_p0 [1]), .IN2(n33965), .IN3(n33952), 
        .IN4(n33934), .QN(n33935) );
  NAND4X0 U37300 ( .IN1(n34441), .IN2(n33937), .IN3(n33936), .IN4(n33935), 
        .QN(n33938) );
  OA21X1 U37301 ( .IN1(n33939), .IN2(n34441), .IN3(n33938), .Q(n33945) );
  AO21X1 U37302 ( .IN1(n33945), .IN2(n33941), .IN3(n33940), .Q(n33947) );
  AO221X1 U37303 ( .IN1(\s15/msel/gnt_p0 [0]), .IN2(n33949), .IN3(n34261), 
        .IN4(n33964), .IN5(n34226), .Q(n33944) );
  NAND2X0 U37304 ( .IN1(n33953), .IN2(n34261), .QN(n33942) );
  NAND3X0 U37305 ( .IN1(n33942), .IN2(n33952), .IN3(n33945), .QN(n33943) );
  NAND3X0 U37306 ( .IN1(\s15/msel/gnt_p0 [2]), .IN2(n33944), .IN3(n33943), 
        .QN(n33946) );
  AO22X1 U37307 ( .IN1(n33947), .IN2(n33946), .IN3(\s15/msel/gnt_p0 [1]), 
        .IN4(n33945), .Q(n17606) );
  NAND2X0 U37308 ( .IN1(n33962), .IN2(n33948), .QN(n33954) );
  OA21X1 U37309 ( .IN1(n33979), .IN2(n33959), .IN3(n33949), .Q(n33950) );
  OA21X1 U37310 ( .IN1(n34261), .IN2(n33954), .IN3(n33950), .Q(n33956) );
  OA21X1 U37311 ( .IN1(n33958), .IN2(n33956), .IN3(n33952), .Q(n33970) );
  AND2X1 U37312 ( .IN1(n33950), .IN2(n33953), .Q(n33955) );
  OA21X1 U37313 ( .IN1(n33953), .IN2(n33952), .IN3(n33951), .Q(n33973) );
  OA22X1 U37314 ( .IN1(n33956), .IN2(n33955), .IN3(n33973), .IN4(n33954), .Q(
        n33957) );
  OA22X1 U37315 ( .IN1(n33970), .IN2(n33967), .IN3(n33958), .IN4(n33957), .Q(
        n33977) );
  OA21X1 U37316 ( .IN1(n33974), .IN2(n33973), .IN3(n33959), .Q(n33968) );
  OR3X1 U37317 ( .IN1(n34226), .IN2(n33979), .IN3(n33968), .Q(n33976) );
  AO221X1 U37318 ( .IN1(n33962), .IN2(\s15/msel/gnt_p0 [0]), .IN3(n33962), 
        .IN4(n33961), .IN5(n33960), .Q(n33963) );
  NAND3X0 U37319 ( .IN1(n33964), .IN2(n33965), .IN3(n33963), .QN(n33972) );
  NAND2X0 U37320 ( .IN1(n33966), .IN2(n33965), .QN(n33969) );
  OA22X1 U37321 ( .IN1(n33970), .IN2(n33969), .IN3(n33968), .IN4(n33967), .Q(
        n33971) );
  OA221X1 U37322 ( .IN1(n33974), .IN2(n33973), .IN3(n33974), .IN4(n33972), 
        .IN5(n33971), .Q(n33975) );
  OA222X1 U37323 ( .IN1(n34441), .IN2(n33977), .IN3(n34441), .IN4(n33976), 
        .IN5(n33975), .IN6(\s15/msel/gnt_p0 [2]), .Q(n33982) );
  OA222X1 U37324 ( .IN1(n33982), .IN2(n33979), .IN3(n33982), .IN4(n34226), 
        .IN5(\s15/msel/gnt_p0 [1]), .IN6(n33978), .Q(n33981) );
  AO21X1 U37325 ( .IN1(n33981), .IN2(n33980), .IN3(\s15/msel/gnt_p0 [2]), .Q(
        n33986) );
  AO221X1 U37326 ( .IN1(n34261), .IN2(n34441), .IN3(n34261), .IN4(n33983), 
        .IN5(n33982), .Q(n33985) );
  NAND3X0 U37327 ( .IN1(n33986), .IN2(n33985), .IN3(n33984), .QN(n17605) );
  NOR2X0 U37328 ( .IN1(n33987), .IN2(n34265), .QN(n34060) );
  INVX0 U37329 ( .INP(n33988), .ZN(n33989) );
  INVX0 U37330 ( .INP(n34022), .ZN(n34036) );
  OA221X1 U37331 ( .IN1(\s15/msel/gnt_p2 [1]), .IN2(n34036), .IN3(n34265), 
        .IN4(n34043), .IN5(n34231), .Q(n34055) );
  NOR2X0 U37332 ( .IN1(n33989), .IN2(n34055), .QN(n33990) );
  OA221X1 U37333 ( .IN1(n34060), .IN2(n34005), .IN3(n34060), .IN4(n34061), 
        .IN5(n33990), .Q(n34000) );
  NAND2X0 U37334 ( .IN1(\s15/msel/gnt_p2 [0]), .IN2(\s15/msel/gnt_p2 [1]), 
        .QN(n34033) );
  NOR2X0 U37335 ( .IN1(n34029), .IN2(n34033), .QN(n34053) );
  NOR2X0 U37336 ( .IN1(\s15/msel/gnt_p2 [2]), .IN2(n34053), .QN(n33993) );
  NOR2X0 U37337 ( .IN1(\s15/msel/gnt_p2 [0]), .IN2(n34265), .QN(n33991) );
  NAND2X0 U37338 ( .IN1(n34040), .IN2(n33991), .QN(n33992) );
  NAND2X0 U37339 ( .IN1(n33993), .IN2(n33992), .QN(n34021) );
  NOR2X0 U37340 ( .IN1(\s15/msel/gnt_p2 [1]), .IN2(n34231), .QN(n34015) );
  NOR2X0 U37341 ( .IN1(n33994), .IN2(\s15/msel/gnt_p2 [1]), .QN(n34014) );
  OA21X1 U37342 ( .IN1(n34015), .IN2(n34014), .IN3(n34008), .Q(n33996) );
  AND2X1 U37343 ( .IN1(\s15/msel/gnt_p2 [1]), .IN2(n34029), .Q(n33995) );
  MUX21X1 U37344 ( .IN1(n34051), .IN2(n34049), .S(\s15/msel/gnt_p2 [0]), .Q(
        n34020) );
  OA22X1 U37345 ( .IN1(n33996), .IN2(n33995), .IN3(\s15/msel/gnt_p2 [1]), 
        .IN4(n34020), .Q(n33998) );
  NAND2X0 U37346 ( .IN1(n33998), .IN2(n33997), .QN(n33999) );
  OAI22X1 U37347 ( .IN1(n34000), .IN2(n34406), .IN3(n34021), .IN4(n33999), 
        .QN(n17604) );
  INVX0 U37348 ( .INP(n34008), .ZN(n34001) );
  NAND2X0 U37349 ( .IN1(n34003), .IN2(n34001), .QN(n34004) );
  NAND2X0 U37350 ( .IN1(n34005), .IN2(n34004), .QN(n34002) );
  AO21X1 U37351 ( .IN1(n34002), .IN2(n34061), .IN3(\s15/msel/gnt_p2 [1]), .Q(
        n34019) );
  NAND2X0 U37352 ( .IN1(n34003), .IN2(n34007), .QN(n34010) );
  NAND3X0 U37353 ( .IN1(n34060), .IN2(n34004), .IN3(n34010), .QN(n34018) );
  INVX0 U37354 ( .INP(n34005), .ZN(n34006) );
  NAND2X0 U37355 ( .IN1(n34007), .IN2(n34006), .QN(n34009) );
  NAND2X0 U37356 ( .IN1(n34008), .IN2(n34009), .QN(n34016) );
  NAND2X0 U37357 ( .IN1(n34010), .IN2(n34009), .QN(n34011) );
  OA21X1 U37358 ( .IN1(n34012), .IN2(n34011), .IN3(\s15/msel/gnt_p2 [1]), .Q(
        n34013) );
  AO221X1 U37359 ( .IN1(n34016), .IN2(n34015), .IN3(n34016), .IN4(n34014), 
        .IN5(n34013), .Q(n34017) );
  OA222X1 U37360 ( .IN1(n34406), .IN2(n34019), .IN3(n34406), .IN4(n34018), 
        .IN5(\s15/msel/gnt_p2 [2]), .IN6(n34017), .Q(n34023) );
  NAND2X0 U37361 ( .IN1(\s15/msel/gnt_p2 [0]), .IN2(\s15/msel/gnt_p2 [2]), 
        .QN(n34059) );
  OA221X1 U37362 ( .IN1(n34021), .IN2(n34020), .IN3(n34021), .IN4(n34023), 
        .IN5(n34059), .Q(n34027) );
  AO22X1 U37363 ( .IN1(\s15/msel/gnt_p2 [1]), .IN2(n34043), .IN3(n34022), 
        .IN4(n34023), .Q(n34026) );
  INVX0 U37364 ( .INP(n34059), .ZN(n34024) );
  OA221X1 U37365 ( .IN1(\s15/msel/gnt_p2 [1]), .IN2(n34024), .IN3(
        \s15/msel/gnt_p2 [1]), .IN4(n34061), .IN5(n34023), .Q(n34025) );
  AO221X1 U37366 ( .IN1(n34027), .IN2(n34406), .IN3(n34027), .IN4(n34026), 
        .IN5(n34025), .Q(n17603) );
  OA21X1 U37367 ( .IN1(n34035), .IN2(n34049), .IN3(n34028), .Q(n34038) );
  OA21X1 U37368 ( .IN1(n34043), .IN2(n34038), .IN3(n34061), .Q(n34041) );
  NOR3X0 U37369 ( .IN1(n34036), .IN2(n34041), .IN3(n34033), .QN(n34048) );
  AO221X1 U37370 ( .IN1(n34038), .IN2(n34035), .IN3(n34038), .IN4(n34231), 
        .IN5(n34036), .Q(n34030) );
  OA21X1 U37371 ( .IN1(n34036), .IN2(n34061), .IN3(n34029), .Q(n34037) );
  OA21X1 U37372 ( .IN1(n34043), .IN2(n34030), .IN3(n34037), .Q(n34031) );
  OA21X1 U37373 ( .IN1(n34040), .IN2(n34037), .IN3(n34049), .Q(n34034) );
  OA22X1 U37374 ( .IN1(n34040), .IN2(n34031), .IN3(n34034), .IN4(
        \s15/msel/gnt_p2 [1]), .Q(n34032) );
  NAND2X0 U37375 ( .IN1(n34032), .IN2(n34406), .QN(n34047) );
  NOR3X0 U37376 ( .IN1(n34035), .IN2(n34034), .IN3(n34033), .QN(n34046) );
  AO221X1 U37377 ( .IN1(n34037), .IN2(n34036), .IN3(n34037), .IN4(n34231), 
        .IN5(n34035), .Q(n34039) );
  OA21X1 U37378 ( .IN1(n34040), .IN2(n34039), .IN3(n34038), .Q(n34042) );
  OA22X1 U37379 ( .IN1(n34043), .IN2(n34042), .IN3(n34041), .IN4(
        \s15/msel/gnt_p2 [1]), .Q(n34044) );
  NAND2X0 U37380 ( .IN1(\s15/msel/gnt_p2 [2]), .IN2(n34044), .QN(n34045) );
  OA22X1 U37381 ( .IN1(n34048), .IN2(n34047), .IN3(n34046), .IN4(n34045), .Q(
        n34054) );
  NOR2X0 U37382 ( .IN1(n34231), .IN2(n34049), .QN(n34050) );
  AO222X1 U37383 ( .IN1(n34054), .IN2(\s15/msel/gnt_p2 [1]), .IN3(n34054), 
        .IN4(n34051), .IN5(n34265), .IN6(n34050), .Q(n34052) );
  OAI21X1 U37384 ( .IN1(n34053), .IN2(n34052), .IN3(n34406), .QN(n34066) );
  INVX0 U37385 ( .INP(n34054), .ZN(n34056) );
  NOR2X0 U37386 ( .IN1(n34056), .IN2(n34055), .QN(n34058) );
  NAND2X0 U37387 ( .IN1(n34231), .IN2(n34406), .QN(n34057) );
  NAND2X0 U37388 ( .IN1(n34058), .IN2(n34057), .QN(n34065) );
  NOR2X0 U37389 ( .IN1(n34060), .IN2(n34059), .QN(n34063) );
  NAND2X0 U37390 ( .IN1(n34265), .IN2(n34061), .QN(n34062) );
  NAND2X0 U37391 ( .IN1(n34063), .IN2(n34062), .QN(n34064) );
  NAND3X0 U37392 ( .IN1(n34066), .IN2(n34065), .IN3(n34064), .QN(n17601) );
  INVX0 U37393 ( .INP(n34067), .ZN(n34069) );
  OAI22X1 U37394 ( .IN1(\s0/msel/pri_out [1]), .IN2(\s0/next ), .IN3(n34069), 
        .IN4(n34068), .QN(n34070) );
  NOR2X0 U37395 ( .IN1(rst_i), .IN2(n34070), .QN(n17598) );
  NAND3X0 U37396 ( .IN1(n34072), .IN2(n34071), .IN3(\s1/next ), .QN(n34082) );
  OA21X1 U37397 ( .IN1(\s1/msel/pri_out [0]), .IN2(\s1/next ), .IN3(n34082), 
        .Q(n34079) );
  NAND4X0 U37398 ( .IN1(n34076), .IN2(n34075), .IN3(n34074), .IN4(n34073), 
        .QN(n34077) );
  AND4X1 U37399 ( .IN1(n34080), .IN2(n34081), .IN3(\s1/next ), .IN4(n34077), 
        .Q(n34078) );
  OA21X1 U37400 ( .IN1(n34079), .IN2(n34078), .IN3(n34690), .Q(n17597) );
  NAND2X0 U37401 ( .IN1(n34081), .IN2(n34080), .QN(n34083) );
  OAI22X1 U37402 ( .IN1(\s1/msel/pri_out [1]), .IN2(\s1/next ), .IN3(n34083), 
        .IN4(n34082), .QN(n34084) );
  NOR2X0 U37403 ( .IN1(rst_i), .IN2(n34084), .QN(n17596) );
  NOR2X0 U37404 ( .IN1(\s2/msel/pri_out [0]), .IN2(\s2/next ), .QN(n34091) );
  NAND2X0 U37405 ( .IN1(n34086), .IN2(n34085), .QN(n34087) );
  NAND4X0 U37406 ( .IN1(n34089), .IN2(n34088), .IN3(\s2/next ), .IN4(n34087), 
        .QN(n34090) );
  OA21X1 U37407 ( .IN1(n34092), .IN2(n34091), .IN3(n34090), .Q(n34093) );
  NOR2X0 U37408 ( .IN1(rst_i), .IN2(n34093), .QN(n17595) );
  OAI22X1 U37409 ( .IN1(\s3/msel/pri_out [1]), .IN2(\s3/next ), .IN3(n34095), 
        .IN4(n34094), .QN(n34096) );
  NOR2X0 U37410 ( .IN1(rst_i), .IN2(n34096), .QN(n17592) );
  OA21X1 U37411 ( .IN1(n34099), .IN2(n34098), .IN3(n34097), .Q(n34104) );
  NAND2X0 U37412 ( .IN1(n34101), .IN2(n34100), .QN(n34102) );
  MUX21X1 U37413 ( .IN1(\s4/msel/pri_out [0]), .IN2(n34102), .S(\s4/next ), 
        .Q(n34103) );
  OA21X1 U37414 ( .IN1(n34104), .IN2(n34103), .IN3(n34678), .Q(n17591) );
  NAND2X0 U37415 ( .IN1(n34106), .IN2(n34105), .QN(n34110) );
  OA221X1 U37416 ( .IN1(n34110), .IN2(n34109), .IN3(n34110), .IN4(n34108), 
        .IN5(n34107), .Q(n34112) );
  NOR2X0 U37417 ( .IN1(\s5/msel/pri_out [0]), .IN2(\s5/next ), .QN(n34111) );
  NOR3X0 U37418 ( .IN1(rst_i), .IN2(n34112), .IN3(n34111), .QN(n17589) );
  NAND3X0 U37419 ( .IN1(n34115), .IN2(n34114), .IN3(n34113), .QN(n34125) );
  MUX21X1 U37420 ( .IN1(\s6/msel/pri_out [0]), .IN2(n34125), .S(\s6/next ), 
        .Q(n34124) );
  NAND4X0 U37421 ( .IN1(n34118), .IN2(n34117), .IN3(n34116), .IN4(\s6/next ), 
        .QN(n34126) );
  INVX0 U37422 ( .INP(n34126), .ZN(n34123) );
  NAND3X0 U37423 ( .IN1(n34121), .IN2(n34120), .IN3(n34119), .QN(n34122) );
  OA221X1 U37424 ( .IN1(n34124), .IN2(n34123), .IN3(n34124), .IN4(n34122), 
        .IN5(n34677), .Q(n17587) );
  OAI22X1 U37425 ( .IN1(\s6/msel/pri_out [1]), .IN2(\s6/next ), .IN3(n34126), 
        .IN4(n34125), .QN(n34127) );
  NOR2X0 U37426 ( .IN1(rst_i), .IN2(n34127), .QN(n17586) );
  NAND3X0 U37427 ( .IN1(n34130), .IN2(n34129), .IN3(n34128), .QN(n34131) );
  NAND4X0 U37428 ( .IN1(n34134), .IN2(n34133), .IN3(n34132), .IN4(n34131), 
        .QN(n34136) );
  AO22X1 U37429 ( .IN1(n34676), .IN2(n34377), .IN3(n34136), .IN4(n34135), .Q(
        n34137) );
  NOR2X0 U37430 ( .IN1(rst_i), .IN2(n34137), .QN(n17585) );
  NOR2X0 U37431 ( .IN1(\s8/msel/pri_out [0]), .IN2(\s8/next ), .QN(n34147) );
  NAND3X0 U37432 ( .IN1(n34140), .IN2(n34139), .IN3(n34138), .QN(n34150) );
  INVX0 U37433 ( .INP(n34141), .ZN(n34144) );
  NOR3X0 U37434 ( .IN1(n34143), .IN2(n34142), .IN3(n34674), .QN(n34148) );
  OA221X1 U37435 ( .IN1(n34150), .IN2(n34145), .IN3(n34150), .IN4(n34144), 
        .IN5(n34148), .Q(n34146) );
  NOR3X0 U37436 ( .IN1(n34147), .IN2(n34146), .IN3(rst_i), .QN(n17583) );
  INVX0 U37437 ( .INP(n34148), .ZN(n34149) );
  OAI22X1 U37438 ( .IN1(n34150), .IN2(n34149), .IN3(\s8/msel/pri_out [1]), 
        .IN4(\s8/next ), .QN(n34151) );
  NOR2X0 U37439 ( .IN1(rst_i), .IN2(n34151), .QN(n17582) );
  NAND4X0 U37440 ( .IN1(n34154), .IN2(n34153), .IN3(n34152), .IN4(\s9/next ), 
        .QN(n34163) );
  INVX0 U37441 ( .INP(n34163), .ZN(n34155) );
  OA21X1 U37442 ( .IN1(n34157), .IN2(n34156), .IN3(n34155), .Q(n34161) );
  OR2X1 U37443 ( .IN1(n34159), .IN2(n34158), .Q(n34162) );
  MUX21X1 U37444 ( .IN1(\s9/msel/pri_out [0]), .IN2(n34162), .S(\s9/next ), 
        .Q(n34160) );
  OA21X1 U37445 ( .IN1(n34161), .IN2(n34160), .IN3(n34681), .Q(n17581) );
  OAI22X1 U37446 ( .IN1(\s9/msel/pri_out [1]), .IN2(\s9/next ), .IN3(n34163), 
        .IN4(n34162), .QN(n34164) );
  NOR2X0 U37447 ( .IN1(rst_i), .IN2(n34164), .QN(n17580) );
  AO22X1 U37448 ( .IN1(n34166), .IN2(n34165), .IN3(n34672), .IN4(n34376), .Q(
        n34167) );
  NOR2X0 U37449 ( .IN1(rst_i), .IN2(n34167), .QN(n17578) );
  NAND3X0 U37450 ( .IN1(n34169), .IN2(n34168), .IN3(\s11/next ), .QN(n34179)
         );
  NOR3X0 U37451 ( .IN1(n34172), .IN2(n34171), .IN3(n34170), .QN(n34178) );
  NAND3X0 U37452 ( .IN1(n34175), .IN2(n34174), .IN3(n34173), .QN(n34176) );
  OA221X1 U37453 ( .IN1(n34179), .IN2(n34178), .IN3(n34179), .IN4(n34176), 
        .IN5(n34690), .Q(n34177) );
  OA21X1 U37454 ( .IN1(\s11/msel/pri_out [0]), .IN2(\s11/next ), .IN3(n34177), 
        .Q(n17577) );
  INVX0 U37455 ( .INP(n34178), .ZN(n34180) );
  OAI22X1 U37456 ( .IN1(\s11/msel/pri_out [1]), .IN2(\s11/next ), .IN3(n34180), 
        .IN4(n34179), .QN(n34181) );
  NOR2X0 U37457 ( .IN1(rst_i), .IN2(n34181), .QN(n17576) );
  NAND3X0 U37458 ( .IN1(n34184), .IN2(n34183), .IN3(n34182), .QN(n34193) );
  MUX21X1 U37459 ( .IN1(\s12/msel/pri_out [0]), .IN2(n34193), .S(\s12/next ), 
        .Q(n34192) );
  NAND3X0 U37460 ( .IN1(n34186), .IN2(n34185), .IN3(\s12/next ), .QN(n34194)
         );
  INVX0 U37461 ( .INP(n34194), .ZN(n34191) );
  NAND3X0 U37462 ( .IN1(n34189), .IN2(n34188), .IN3(n34187), .QN(n34190) );
  OA221X1 U37463 ( .IN1(n34192), .IN2(n34191), .IN3(n34192), .IN4(n34190), 
        .IN5(n34686), .Q(n17575) );
  OAI22X1 U37464 ( .IN1(\s12/msel/pri_out [1]), .IN2(\s12/next ), .IN3(n34194), 
        .IN4(n34193), .QN(n34195) );
  NOR2X0 U37465 ( .IN1(rst_i), .IN2(n34195), .QN(n17574) );
  NAND4X0 U37466 ( .IN1(n34198), .IN2(n34197), .IN3(n34196), .IN4(\s13/next ), 
        .QN(n34207) );
  NOR2X0 U37467 ( .IN1(n34200), .IN2(n34199), .QN(n34206) );
  NAND3X0 U37468 ( .IN1(n34203), .IN2(n34202), .IN3(n34201), .QN(n34204) );
  OA221X1 U37469 ( .IN1(n34207), .IN2(n34206), .IN3(n34207), .IN4(n34204), 
        .IN5(n34683), .Q(n34205) );
  OA21X1 U37470 ( .IN1(\s13/msel/pri_out [0]), .IN2(\s13/next ), .IN3(n34205), 
        .Q(n17573) );
  INVX0 U37471 ( .INP(n34206), .ZN(n34208) );
  OAI22X1 U37472 ( .IN1(\s13/msel/pri_out [1]), .IN2(\s13/next ), .IN3(n34208), 
        .IN4(n34207), .QN(n34209) );
  NOR2X0 U37473 ( .IN1(rst_i), .IN2(n34209), .QN(n17572) );
  NAND2X0 U37474 ( .IN1(n34211), .IN2(n34210), .QN(n34212) );
  MUX21X1 U37475 ( .IN1(\s14/msel/pri_out [0]), .IN2(n34212), .S(\s14/next ), 
        .Q(n34218) );
  NAND3X0 U37476 ( .IN1(n34215), .IN2(n34214), .IN3(n34213), .QN(n34216) );
  OA221X1 U37477 ( .IN1(n34218), .IN2(n34217), .IN3(n34218), .IN4(n34216), 
        .IN5(n34692), .Q(n17571) );
  INVX0 U37478 ( .INP(n34219), .ZN(n34221) );
  OAI22X1 U37479 ( .IN1(\s15/msel/pri_out [1]), .IN2(\s15/next ), .IN3(n34221), 
        .IN4(n34220), .QN(n34222) );
  NOR2X0 U37480 ( .IN1(rst_i), .IN2(n34222), .QN(n17568) );
endmodule

