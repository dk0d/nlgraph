module b14 ( clock, reset, \addr[19] , \addr[18] , \addr[17] , 
        \addr[16] , \addr[15] , \addr[14] , \addr[13] , \addr[12] , \addr[11] , 
        \addr[10] , \addr[9] , \addr[8] , \addr[7] , \addr[6] , \addr[5] , 
        \addr[4] , \addr[3] , \addr[2] , \addr[1] , \addr[0] ,
        \datai[31] , \datai[30] , \datai[29] , \datai[28] , \datai[27] , 
        \datai[26] , \datai[25] , \datai[24] , \datai[23] , \datai[22] , 
        \datai[21] , \datai[20] , \datai[19] , \datai[18] , \datai[17] , 
        \datai[16] , \datai[15] , \datai[14] , \datai[13] , \datai[12] , 
        \datai[11] , \datai[10] , \datai[9] , \datai[8] , \datai[7] , 
        \datai[6] , \datai[5] , \datai[4] , \datai[3] , \datai[2] , \datai[1] , 
        \datai[0] , \datao[31] , \datao[30] , \datao[29] , 
        \datao[28] , \datao[27] , \datao[26] , \datao[25] , \datao[24] , 
        \datao[23] , \datao[22] , \datao[21] , \datao[20] , \datao[19] , 
        \datao[18] , \datao[17] , \datao[16] , \datao[15] , \datao[14] , 
        \datao[13] , \datao[12] , \datao[11] , \datao[10] , \datao[9] , 
        \datao[8] , \datao[7] , \datao[6] , \datao[5] , \datao[4] , \datao[3] , 
        \datao[2] , \datao[1] , \datao[0] , rd, wr );
  input clock, reset, \datai[31] , \datai[30] , \datai[29] , \datai[28] ,
         \datai[27] , \datai[26] , \datai[25] , \datai[24] , \datai[23] ,
         \datai[22] , \datai[21] , \datai[20] , \datai[19] , \datai[18] ,
         \datai[17] , \datai[16] , \datai[15] , \datai[14] , \datai[13] ,
         \datai[12] , \datai[11] , \datai[10] , \datai[9] , \datai[8] ,
         \datai[7] , \datai[6] , \datai[5] , \datai[4] , \datai[3] ,
         \datai[2] , \datai[1] , \datai[0] ;
  output \addr[19] , \addr[18] , \addr[17] , \addr[16] , \addr[15] ,
         \addr[14] , \addr[13] , \addr[12] , \addr[11] , \addr[10] , \addr[9] ,
         \addr[8] , \addr[7] , \addr[6] , \addr[5] , \addr[4] , \addr[3] ,
         \addr[2] , \addr[1] , \addr[0] , \datao[31] , \datao[30] ,
         \datao[29] , \datao[28] , \datao[27] , \datao[26] , \datao[25] ,
         \datao[24] , \datao[23] , \datao[22] , \datao[21] , \datao[20] ,
         \datao[19] , \datao[18] , \datao[17] , \datao[16] , \datao[15] ,
         \datao[14] , \datao[13] , \datao[12] , \datao[11] , \datao[10] ,
         \datao[9] , \datao[8] , \datao[7] , \datao[6] , \datao[5] ,
         \datao[4] , \datao[3] , \datao[2] , \datao[1] , \datao[0] , rd, wr;
  wire   B, state, N5560, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736;
  wire   [19:0] addr;
  wire   [31:0] datai;
  wire   [31:0] datao;
  wire   [31:0] IR;
  wire   [31:0] d;
  wire   [31:0] reg0;
  wire   [31:0] reg1;
  wire   [31:0] reg2;
  wire   [28:0] reg3;

  DFFARX1 state_reg ( .D(n2703), .CLK(clock), .RSTB(n2735), .Q(state), .QN(
        n2703) );
  DFFARX1 \IR_reg[0]  ( .D(n893), .CLK(clock), .RSTB(n2729), .Q(IR[0]), .QN(
        n2702) );
  DFFARX1 \IR_reg[1]  ( .D(n892), .CLK(clock), .RSTB(n2732), .Q(IR[1]) );
  DFFARX1 \IR_reg[2]  ( .D(n891), .CLK(clock), .RSTB(n2734), .Q(IR[2]), .QN(
        n2701) );
  DFFARX1 \IR_reg[3]  ( .D(n890), .CLK(clock), .RSTB(n2728), .Q(IR[3]) );
  DFFARX1 \IR_reg[4]  ( .D(n889), .CLK(clock), .RSTB(n2734), .Q(IR[4]) );
  DFFARX1 \IR_reg[5]  ( .D(n888), .CLK(clock), .RSTB(n2730), .Q(IR[5]) );
  DFFARX1 \IR_reg[6]  ( .D(n887), .CLK(clock), .RSTB(n2732), .Q(IR[6]) );
  DFFARX1 \IR_reg[7]  ( .D(n886), .CLK(clock), .RSTB(n2732), .Q(IR[7]) );
  DFFARX1 \IR_reg[8]  ( .D(n885), .CLK(clock), .RSTB(n2732), .Q(IR[8]) );
  DFFARX1 \IR_reg[9]  ( .D(n884), .CLK(clock), .RSTB(n2734), .Q(IR[9]) );
  DFFARX1 \IR_reg[10]  ( .D(n883), .CLK(clock), .RSTB(n2732), .Q(IR[10]) );
  DFFARX1 \IR_reg[11]  ( .D(n882), .CLK(clock), .RSTB(n2734), .Q(IR[11]) );
  DFFARX1 \IR_reg[12]  ( .D(n881), .CLK(clock), .RSTB(n2735), .Q(IR[12]) );
  DFFARX1 \IR_reg[13]  ( .D(n880), .CLK(clock), .RSTB(n2734), .Q(IR[13]) );
  DFFARX1 \IR_reg[14]  ( .D(n879), .CLK(clock), .RSTB(n2731), .Q(IR[14]) );
  DFFARX1 \IR_reg[15]  ( .D(n878), .CLK(clock), .RSTB(n2730), .Q(IR[15]) );
  DFFARX1 \IR_reg[16]  ( .D(n877), .CLK(clock), .RSTB(n2733), .Q(IR[16]) );
  DFFARX1 \IR_reg[17]  ( .D(n876), .CLK(clock), .RSTB(n2729), .Q(IR[17]) );
  DFFARX1 \IR_reg[18]  ( .D(n875), .CLK(clock), .RSTB(n2728), .Q(IR[18]) );
  DFFARX1 \IR_reg[19]  ( .D(n874), .CLK(clock), .RSTB(n2729), .Q(IR[19]) );
  DFFARX1 \IR_reg[20]  ( .D(n873), .CLK(clock), .RSTB(n2731), .Q(IR[20]), .QN(
        n2706) );
  DFFARX1 \IR_reg[21]  ( .D(n872), .CLK(clock), .RSTB(n2731), .Q(IR[21]), .QN(
        n2712) );
  DFFARX1 \IR_reg[22]  ( .D(n871), .CLK(clock), .RSTB(n2728), .Q(IR[22]), .QN(
        n2708) );
  DFFARX1 \IR_reg[23]  ( .D(n870), .CLK(clock), .RSTB(n2732), .Q(IR[23]), .QN(
        n2710) );
  DFFARX1 \IR_reg[24]  ( .D(n869), .CLK(clock), .RSTB(n2728), .Q(IR[24]), .QN(
        n2705) );
  DFFARX1 \IR_reg[25]  ( .D(n868), .CLK(clock), .RSTB(n2728), .Q(IR[25]), .QN(
        n2711) );
  DFFARX1 \IR_reg[26]  ( .D(n867), .CLK(clock), .RSTB(n2729), .Q(IR[26]), .QN(
        n2707) );
  DFFARX1 \IR_reg[27]  ( .D(n866), .CLK(clock), .RSTB(n2733), .Q(IR[27]), .QN(
        n2724) );
  DFFARX1 \IR_reg[28]  ( .D(n865), .CLK(clock), .RSTB(n2730), .Q(IR[28]), .QN(
        n2725) );
  DFFARX1 \IR_reg[29]  ( .D(n864), .CLK(clock), .RSTB(n2731), .Q(IR[29]) );
  DFFARX1 \IR_reg[30]  ( .D(n863), .CLK(clock), .RSTB(n2735), .Q(IR[30]), .QN(
        n2726) );
  DFFARX1 \IR_reg[31]  ( .D(n862), .CLK(clock), .RSTB(n2728), .Q(n2699), .QN(
        n2727) );
  DFFARX1 \reg2_reg[0]  ( .D(n989), .CLK(clock), .RSTB(n2728), .Q(reg2[0]) );
  DFFARX1 \reg2_reg[1]  ( .D(n988), .CLK(clock), .RSTB(n2735), .Q(reg2[1]) );
  DFFARX1 \reg2_reg[2]  ( .D(n987), .CLK(clock), .RSTB(n2730), .Q(reg2[2]) );
  DFFARX1 \reg2_reg[3]  ( .D(n986), .CLK(clock), .RSTB(n2734), .Q(reg2[3]) );
  DFFARX1 \reg2_reg[4]  ( .D(n985), .CLK(clock), .RSTB(n2730), .Q(reg2[4]) );
  DFFARX1 \reg2_reg[5]  ( .D(n984), .CLK(clock), .RSTB(n2730), .Q(reg2[5]) );
  DFFARX1 \reg2_reg[6]  ( .D(n983), .CLK(clock), .RSTB(n2729), .Q(reg2[6]) );
  DFFARX1 \reg2_reg[7]  ( .D(n982), .CLK(clock), .RSTB(n2730), .Q(reg2[7]) );
  DFFARX1 \reg2_reg[8]  ( .D(n981), .CLK(clock), .RSTB(n2735), .Q(reg2[8]) );
  DFFARX1 \reg2_reg[9]  ( .D(n980), .CLK(clock), .RSTB(n2730), .Q(reg2[9]) );
  DFFARX1 \reg2_reg[10]  ( .D(n979), .CLK(clock), .RSTB(n2735), .Q(reg2[10])
         );
  DFFARX1 \reg2_reg[11]  ( .D(n978), .CLK(clock), .RSTB(n2732), .Q(reg2[11])
         );
  DFFARX1 \reg2_reg[12]  ( .D(n977), .CLK(clock), .RSTB(n2731), .Q(reg2[12])
         );
  DFFARX1 \reg2_reg[13]  ( .D(n976), .CLK(clock), .RSTB(n2731), .Q(reg2[13])
         );
  DFFARX1 \reg2_reg[14]  ( .D(n975), .CLK(clock), .RSTB(n2729), .Q(reg2[14])
         );
  DFFARX1 \reg2_reg[15]  ( .D(n974), .CLK(clock), .RSTB(n2732), .Q(reg2[15])
         );
  DFFARX1 \reg2_reg[16]  ( .D(n973), .CLK(clock), .RSTB(n2730), .Q(reg2[16])
         );
  DFFARX1 \reg2_reg[17]  ( .D(n972), .CLK(clock), .RSTB(n2728), .Q(reg2[17])
         );
  DFFARX1 \reg2_reg[18]  ( .D(n971), .CLK(clock), .RSTB(n2733), .Q(reg2[18])
         );
  DFFARX1 \reg2_reg[19]  ( .D(n970), .CLK(clock), .RSTB(n2731), .Q(reg2[19])
         );
  DFFARX1 \reg2_reg[20]  ( .D(n969), .CLK(clock), .RSTB(n2732), .Q(reg2[20])
         );
  DFFARX1 \reg2_reg[21]  ( .D(n968), .CLK(clock), .RSTB(n2735), .Q(reg2[21])
         );
  DFFARX1 \reg2_reg[22]  ( .D(n967), .CLK(clock), .RSTB(n2732), .Q(reg2[22])
         );
  DFFARX1 \reg2_reg[23]  ( .D(n966), .CLK(clock), .RSTB(n2728), .Q(reg2[23])
         );
  DFFARX1 \reg2_reg[24]  ( .D(n965), .CLK(clock), .RSTB(n2729), .Q(reg2[24])
         );
  DFFARX1 \reg2_reg[25]  ( .D(n964), .CLK(clock), .RSTB(n2733), .Q(reg2[25])
         );
  DFFARX1 \reg2_reg[26]  ( .D(n963), .CLK(clock), .RSTB(n2730), .Q(reg2[26])
         );
  DFFARX1 \reg2_reg[27]  ( .D(n962), .CLK(clock), .RSTB(n2731), .Q(reg2[27])
         );
  DFFARX1 \reg2_reg[28]  ( .D(n961), .CLK(clock), .RSTB(n2735), .Q(reg2[28])
         );
  DFFARX1 \reg2_reg[29]  ( .D(n960), .CLK(clock), .RSTB(n2734), .Q(reg2[29])
         );
  DFFARX1 \reg2_reg[30]  ( .D(n959), .CLK(clock), .RSTB(n2732), .Q(reg2[30])
         );
  DFFARX1 \reg2_reg[31]  ( .D(n958), .CLK(clock), .RSTB(n2734), .Q(reg2[31])
         );
  DFFARX1 \reg1_reg[0]  ( .D(n957), .CLK(clock), .RSTB(n2733), .Q(reg1[0]) );
  DFFARX1 \reg1_reg[1]  ( .D(n956), .CLK(clock), .RSTB(n2732), .Q(reg1[1]) );
  DFFARX1 \reg1_reg[2]  ( .D(n955), .CLK(clock), .RSTB(n2729), .Q(reg1[2]) );
  DFFARX1 \reg1_reg[3]  ( .D(n954), .CLK(clock), .RSTB(n2728), .Q(reg1[3]) );
  DFFARX1 \reg1_reg[4]  ( .D(n953), .CLK(clock), .RSTB(n2729), .Q(reg1[4]) );
  DFFARX1 \reg1_reg[5]  ( .D(n952), .CLK(clock), .RSTB(n2728), .Q(reg1[5]) );
  DFFARX1 \reg1_reg[6]  ( .D(n951), .CLK(clock), .RSTB(n2733), .Q(reg1[6]) );
  DFFARX1 \reg1_reg[7]  ( .D(n950), .CLK(clock), .RSTB(n2731), .Q(reg1[7]) );
  DFFARX1 \reg1_reg[8]  ( .D(n949), .CLK(clock), .RSTB(n2734), .Q(reg1[8]) );
  DFFARX1 \reg1_reg[9]  ( .D(n948), .CLK(clock), .RSTB(n2731), .Q(reg1[9]) );
  DFFARX1 \reg1_reg[10]  ( .D(n947), .CLK(clock), .RSTB(n2734), .Q(reg1[10])
         );
  DFFARX1 \reg1_reg[11]  ( .D(n946), .CLK(clock), .RSTB(n2733), .Q(reg1[11])
         );
  DFFARX1 \reg1_reg[12]  ( .D(n945), .CLK(clock), .RSTB(n2733), .Q(reg1[12])
         );
  DFFARX1 \reg1_reg[13]  ( .D(n944), .CLK(clock), .RSTB(n2728), .Q(reg1[13])
         );
  DFFARX1 \reg1_reg[14]  ( .D(n943), .CLK(clock), .RSTB(n2733), .Q(reg1[14])
         );
  DFFARX1 \reg1_reg[15]  ( .D(n942), .CLK(clock), .RSTB(n2735), .Q(reg1[15])
         );
  DFFARX1 \reg1_reg[16]  ( .D(n941), .CLK(clock), .RSTB(n2735), .Q(reg1[16])
         );
  DFFARX1 \reg1_reg[17]  ( .D(n940), .CLK(clock), .RSTB(n2729), .Q(reg1[17])
         );
  DFFARX1 \reg1_reg[18]  ( .D(n939), .CLK(clock), .RSTB(n2730), .Q(reg1[18])
         );
  DFFARX1 \reg1_reg[19]  ( .D(n938), .CLK(clock), .RSTB(n2735), .Q(reg1[19])
         );
  DFFARX1 \reg1_reg[20]  ( .D(n937), .CLK(clock), .RSTB(n2730), .Q(reg1[20])
         );
  DFFARX1 \reg1_reg[21]  ( .D(n936), .CLK(clock), .RSTB(n2734), .Q(reg1[21])
         );
  DFFARX1 \reg1_reg[22]  ( .D(n935), .CLK(clock), .RSTB(n2731), .Q(reg1[22])
         );
  DFFARX1 \reg1_reg[23]  ( .D(n934), .CLK(clock), .RSTB(n2732), .Q(reg1[23])
         );
  DFFARX1 \reg1_reg[24]  ( .D(n933), .CLK(clock), .RSTB(n2735), .Q(reg1[24])
         );
  DFFARX1 \reg1_reg[25]  ( .D(n932), .CLK(clock), .RSTB(n2729), .Q(reg1[25])
         );
  DFFARX1 \reg1_reg[26]  ( .D(n931), .CLK(clock), .RSTB(n2734), .Q(reg1[26])
         );
  DFFARX1 \reg1_reg[27]  ( .D(n930), .CLK(clock), .RSTB(n2733), .Q(reg1[27])
         );
  DFFARX1 \reg1_reg[28]  ( .D(n929), .CLK(clock), .RSTB(n2732), .Q(reg1[28])
         );
  DFFARX1 \reg1_reg[29]  ( .D(n928), .CLK(clock), .RSTB(n2729), .Q(reg1[29])
         );
  DFFARX1 \reg1_reg[30]  ( .D(n927), .CLK(clock), .RSTB(n2728), .Q(reg1[30])
         );
  DFFARX1 \reg1_reg[31]  ( .D(n926), .CLK(clock), .RSTB(n2729), .Q(reg1[31])
         );
  DFFARX1 \reg0_reg[0]  ( .D(n925), .CLK(clock), .RSTB(n2733), .Q(reg0[0]) );
  DFFARX1 \reg0_reg[1]  ( .D(n924), .CLK(clock), .RSTB(n2730), .Q(reg0[1]) );
  DFFARX1 \reg0_reg[2]  ( .D(n923), .CLK(clock), .RSTB(n2731), .Q(reg0[2]) );
  DFFARX1 \reg0_reg[3]  ( .D(n922), .CLK(clock), .RSTB(n2735), .Q(reg0[3]) );
  DFFARX1 \reg0_reg[4]  ( .D(n921), .CLK(clock), .RSTB(n2730), .Q(reg0[4]) );
  DFFARX1 \reg0_reg[5]  ( .D(n920), .CLK(clock), .RSTB(n2731), .Q(reg0[5]) );
  DFFARX1 \reg0_reg[6]  ( .D(n919), .CLK(clock), .RSTB(n2735), .Q(reg0[6]) );
  DFFARX1 \reg0_reg[7]  ( .D(n918), .CLK(clock), .RSTB(n2734), .Q(reg0[7]) );
  DFFARX1 \reg0_reg[8]  ( .D(n917), .CLK(clock), .RSTB(n2732), .Q(reg0[8]) );
  DFFARX1 \reg0_reg[9]  ( .D(n916), .CLK(clock), .RSTB(n2728), .Q(reg0[9]) );
  DFFARX1 \reg0_reg[10]  ( .D(n915), .CLK(clock), .RSTB(n2729), .Q(reg0[10])
         );
  DFFARX1 \reg0_reg[11]  ( .D(n914), .CLK(clock), .RSTB(n2733), .Q(reg0[11])
         );
  DFFARX1 \reg0_reg[12]  ( .D(n913), .CLK(clock), .RSTB(n2730), .Q(reg0[12])
         );
  DFFARX1 \reg0_reg[13]  ( .D(n912), .CLK(clock), .RSTB(n2731), .Q(reg0[13])
         );
  DFFARX1 \reg0_reg[14]  ( .D(n911), .CLK(clock), .RSTB(n2735), .Q(reg0[14])
         );
  DFFARX1 \reg0_reg[15]  ( .D(n910), .CLK(clock), .RSTB(n2734), .Q(reg0[15])
         );
  DFFARX1 \reg0_reg[16]  ( .D(n909), .CLK(clock), .RSTB(n2728), .Q(reg0[16])
         );
  DFFARX1 \reg0_reg[17]  ( .D(n908), .CLK(clock), .RSTB(n2728), .Q(reg0[17])
         );
  DFFARX1 \reg0_reg[18]  ( .D(n907), .CLK(clock), .RSTB(n2728), .Q(reg0[18])
         );
  DFFARX1 \reg0_reg[19]  ( .D(n906), .CLK(clock), .RSTB(n2728), .Q(reg0[19])
         );
  DFFARX1 \reg0_reg[20]  ( .D(n905), .CLK(clock), .RSTB(n2728), .Q(reg0[20])
         );
  DFFARX1 \reg0_reg[21]  ( .D(n904), .CLK(clock), .RSTB(n2728), .Q(reg0[21])
         );
  DFFARX1 \reg0_reg[22]  ( .D(n903), .CLK(clock), .RSTB(n2728), .Q(reg0[22])
         );
  DFFARX1 \reg0_reg[23]  ( .D(n902), .CLK(clock), .RSTB(n2728), .Q(reg0[23])
         );
  DFFARX1 \reg0_reg[24]  ( .D(n901), .CLK(clock), .RSTB(n2728), .Q(reg0[24])
         );
  DFFARX1 \reg0_reg[25]  ( .D(n900), .CLK(clock), .RSTB(n2728), .Q(reg0[25])
         );
  DFFARX1 \reg0_reg[26]  ( .D(n899), .CLK(clock), .RSTB(n2728), .Q(reg0[26])
         );
  DFFARX1 \reg0_reg[27]  ( .D(n898), .CLK(clock), .RSTB(n2728), .Q(reg0[27])
         );
  DFFARX1 \reg0_reg[28]  ( .D(n897), .CLK(clock), .RSTB(n2729), .Q(reg0[28])
         );
  DFFARX1 \reg0_reg[29]  ( .D(n896), .CLK(clock), .RSTB(n2729), .Q(reg0[29])
         );
  DFFARX1 \reg0_reg[30]  ( .D(n895), .CLK(clock), .RSTB(n2729), .Q(reg0[30])
         );
  DFFARX1 \reg0_reg[31]  ( .D(n894), .CLK(clock), .RSTB(n2729), .Q(reg0[31])
         );
  DFFARX1 \datao_reg[0]  ( .D(n861), .CLK(clock), .RSTB(n2729), .Q(datao[0])
         );
  DFFARX1 \datao_reg[1]  ( .D(n860), .CLK(clock), .RSTB(n2729), .Q(datao[1])
         );
  DFFARX1 \datao_reg[2]  ( .D(n859), .CLK(clock), .RSTB(n2729), .Q(datao[2])
         );
  DFFARX1 \datao_reg[3]  ( .D(n858), .CLK(clock), .RSTB(n2729), .Q(datao[3])
         );
  DFFARX1 \datao_reg[4]  ( .D(n857), .CLK(clock), .RSTB(n2729), .Q(datao[4])
         );
  DFFARX1 \datao_reg[5]  ( .D(n856), .CLK(clock), .RSTB(n2729), .Q(datao[5])
         );
  DFFARX1 \datao_reg[6]  ( .D(n855), .CLK(clock), .RSTB(n2729), .Q(datao[6])
         );
  DFFARX1 \datao_reg[7]  ( .D(n854), .CLK(clock), .RSTB(n2729), .Q(datao[7])
         );
  DFFARX1 \datao_reg[8]  ( .D(n853), .CLK(clock), .RSTB(n2730), .Q(datao[8])
         );
  DFFARX1 \datao_reg[9]  ( .D(n852), .CLK(clock), .RSTB(n2730), .Q(datao[9])
         );
  DFFARX1 \datao_reg[10]  ( .D(n851), .CLK(clock), .RSTB(n2730), .Q(datao[10])
         );
  DFFARX1 \datao_reg[11]  ( .D(n850), .CLK(clock), .RSTB(n2730), .Q(datao[11])
         );
  DFFARX1 \datao_reg[12]  ( .D(n849), .CLK(clock), .RSTB(n2730), .Q(datao[12])
         );
  DFFARX1 \datao_reg[13]  ( .D(n848), .CLK(clock), .RSTB(n2730), .Q(datao[13])
         );
  DFFARX1 \datao_reg[14]  ( .D(n847), .CLK(clock), .RSTB(n2730), .Q(datao[14])
         );
  DFFARX1 \datao_reg[15]  ( .D(n846), .CLK(clock), .RSTB(n2730), .Q(datao[15])
         );
  DFFARX1 \datao_reg[16]  ( .D(n845), .CLK(clock), .RSTB(n2730), .Q(datao[16])
         );
  DFFARX1 \datao_reg[17]  ( .D(n844), .CLK(clock), .RSTB(n2730), .Q(datao[17])
         );
  DFFARX1 \datao_reg[18]  ( .D(n843), .CLK(clock), .RSTB(n2730), .Q(datao[18])
         );
  DFFARX1 \datao_reg[19]  ( .D(n842), .CLK(clock), .RSTB(n2730), .Q(datao[19])
         );
  DFFARX1 \datao_reg[20]  ( .D(n841), .CLK(clock), .RSTB(n2731), .Q(datao[20])
         );
  DFFARX1 \datao_reg[21]  ( .D(n840), .CLK(clock), .RSTB(n2731), .Q(datao[21])
         );
  DFFARX1 \datao_reg[22]  ( .D(n839), .CLK(clock), .RSTB(n2731), .Q(datao[22])
         );
  DFFARX1 \datao_reg[23]  ( .D(n838), .CLK(clock), .RSTB(n2731), .Q(datao[23])
         );
  DFFARX1 \datao_reg[24]  ( .D(n837), .CLK(clock), .RSTB(n2731), .Q(datao[24])
         );
  DFFARX1 \datao_reg[25]  ( .D(n836), .CLK(clock), .RSTB(n2731), .Q(datao[25])
         );
  DFFARX1 \datao_reg[26]  ( .D(n835), .CLK(clock), .RSTB(n2731), .Q(datao[26])
         );
  DFFARX1 \datao_reg[27]  ( .D(n834), .CLK(clock), .RSTB(n2731), .Q(datao[27])
         );
  DFFARX1 \datao_reg[28]  ( .D(n833), .CLK(clock), .RSTB(n2731), .Q(datao[28])
         );
  DFFARX1 \datao_reg[29]  ( .D(n832), .CLK(clock), .RSTB(n2731), .Q(datao[29])
         );
  DFFARX1 \datao_reg[30]  ( .D(n831), .CLK(clock), .RSTB(n2731), .Q(datao[30])
         );
  DFFARX1 \datao_reg[31]  ( .D(n830), .CLK(clock), .RSTB(n2731), .Q(datao[31])
         );
  DFFARX1 wr_reg ( .D(n2736), .CLK(clock), .RSTB(n2732), .Q(wr) );
  DFFARX1 B_reg ( .D(n829), .CLK(clock), .RSTB(n2732), .Q(B), .QN(n2704) );
  DFFARX1 \d_reg[0]  ( .D(n828), .CLK(clock), .RSTB(n2732), .Q(d[0]), .QN(
        n2700) );
  DFFARX1 \d_reg[1]  ( .D(n827), .CLK(clock), .RSTB(n2732), .Q(d[1]), .QN(
        n2709) );
  DFFARX1 rd_reg ( .D(N5560), .CLK(clock), .RSTB(n2732), .Q(rd) );
  DFFARX1 \addr_reg[0]  ( .D(n826), .CLK(clock), .RSTB(n2732), .Q(addr[0]) );
  DFFARX1 \addr_reg[1]  ( .D(n825), .CLK(clock), .RSTB(n2732), .Q(addr[1]) );
  DFFARX1 \addr_reg[2]  ( .D(n824), .CLK(clock), .RSTB(n2732), .Q(addr[2]) );
  DFFARX1 \addr_reg[3]  ( .D(n823), .CLK(clock), .RSTB(n2732), .Q(addr[3]) );
  DFFARX1 \addr_reg[4]  ( .D(n822), .CLK(clock), .RSTB(n2735), .Q(addr[4]) );
  DFFARX1 \addr_reg[5]  ( .D(n821), .CLK(clock), .RSTB(n2732), .Q(addr[5]) );
  DFFARX1 \addr_reg[6]  ( .D(n820), .CLK(clock), .RSTB(n2732), .Q(addr[6]) );
  DFFARX1 \addr_reg[7]  ( .D(n819), .CLK(clock), .RSTB(n2732), .Q(addr[7]) );
  DFFARX1 \addr_reg[8]  ( .D(n818), .CLK(clock), .RSTB(n2733), .Q(addr[8]) );
  DFFARX1 \addr_reg[9]  ( .D(n817), .CLK(clock), .RSTB(n2733), .Q(addr[9]) );
  DFFARX1 \addr_reg[10]  ( .D(n816), .CLK(clock), .RSTB(n2733), .Q(addr[10])
         );
  DFFARX1 \addr_reg[11]  ( .D(n815), .CLK(clock), .RSTB(n2733), .Q(addr[11])
         );
  DFFARX1 \addr_reg[12]  ( .D(n814), .CLK(clock), .RSTB(n2733), .Q(addr[12])
         );
  DFFARX1 \addr_reg[13]  ( .D(n813), .CLK(clock), .RSTB(n2733), .Q(addr[13])
         );
  DFFARX1 \addr_reg[14]  ( .D(n812), .CLK(clock), .RSTB(n2733), .Q(addr[14])
         );
  DFFARX1 \addr_reg[15]  ( .D(n811), .CLK(clock), .RSTB(n2733), .Q(addr[15])
         );
  DFFARX1 \addr_reg[16]  ( .D(n810), .CLK(clock), .RSTB(n2733), .Q(addr[16])
         );
  DFFARX1 \addr_reg[17]  ( .D(n809), .CLK(clock), .RSTB(n2733), .Q(addr[17])
         );
  DFFARX1 \addr_reg[18]  ( .D(n808), .CLK(clock), .RSTB(n2733), .Q(addr[18])
         );
  DFFARX1 \addr_reg[19]  ( .D(n806), .CLK(clock), .RSTB(n2733), .Q(addr[19])
         );
  DFFARX1 \reg3_reg[0]  ( .D(n805), .CLK(clock), .RSTB(n2729), .Q(reg3[0]) );
  DFFARX1 \reg3_reg[1]  ( .D(n804), .CLK(clock), .RSTB(n2734), .Q(reg3[1]) );
  DFFARX1 \reg3_reg[2]  ( .D(n803), .CLK(clock), .RSTB(n2731), .Q(reg3[2]) );
  DFFARX1 \reg3_reg[3]  ( .D(n802), .CLK(clock), .RSTB(n2733), .Q(reg3[3]), 
        .QN(n2698) );
  DFFARX1 \reg3_reg[4]  ( .D(n801), .CLK(clock), .RSTB(n2734), .Q(reg3[4]) );
  DFFARX1 \reg3_reg[5]  ( .D(n800), .CLK(clock), .RSTB(n2734), .Q(reg3[5]) );
  DFFARX1 \reg3_reg[6]  ( .D(n799), .CLK(clock), .RSTB(n2734), .Q(reg3[6]) );
  DFFARX1 \reg3_reg[7]  ( .D(n798), .CLK(clock), .RSTB(n2734), .Q(reg3[7]), 
        .QN(n2713) );
  DFFARX1 \reg3_reg[8]  ( .D(n797), .CLK(clock), .RSTB(n2734), .Q(reg3[8]) );
  DFFARX1 \reg3_reg[9]  ( .D(n796), .CLK(clock), .RSTB(n2734), .Q(reg3[9]), 
        .QN(n2714) );
  DFFARX1 \reg3_reg[10]  ( .D(n795), .CLK(clock), .RSTB(n2734), .Q(reg3[10])
         );
  DFFARX1 \reg3_reg[11]  ( .D(n794), .CLK(clock), .RSTB(n2734), .Q(reg3[11]), 
        .QN(n2715) );
  DFFARX1 \reg3_reg[12]  ( .D(n793), .CLK(clock), .RSTB(n2734), .Q(reg3[12])
         );
  DFFARX1 \reg3_reg[13]  ( .D(n792), .CLK(clock), .RSTB(n2734), .Q(reg3[13]), 
        .QN(n2716) );
  DFFARX1 \reg3_reg[14]  ( .D(n791), .CLK(clock), .RSTB(n2734), .Q(reg3[14])
         );
  DFFARX1 \reg3_reg[15]  ( .D(n790), .CLK(clock), .RSTB(n2734), .Q(reg3[15]), 
        .QN(n2717) );
  DFFARX1 \reg3_reg[16]  ( .D(n789), .CLK(clock), .RSTB(n2735), .Q(reg3[16])
         );
  DFFARX1 \reg3_reg[17]  ( .D(n788), .CLK(clock), .RSTB(n2735), .Q(reg3[17]), 
        .QN(n2718) );
  DFFARX1 \reg3_reg[18]  ( .D(n787), .CLK(clock), .RSTB(n2735), .Q(reg3[18])
         );
  DFFARX1 \reg3_reg[19]  ( .D(n786), .CLK(clock), .RSTB(n2735), .Q(reg3[19]), 
        .QN(n2719) );
  DFFARX1 \reg3_reg[20]  ( .D(n785), .CLK(clock), .RSTB(n2728), .Q(reg3[20])
         );
  DFFARX1 \reg3_reg[21]  ( .D(n784), .CLK(clock), .RSTB(n2735), .Q(reg3[21]), 
        .QN(n2720) );
  DFFARX1 \reg3_reg[22]  ( .D(n783), .CLK(clock), .RSTB(n2733), .Q(reg3[22])
         );
  DFFARX1 \reg3_reg[23]  ( .D(n782), .CLK(clock), .RSTB(n2735), .Q(reg3[23]), 
        .QN(n2721) );
  DFFARX1 \reg3_reg[24]  ( .D(n781), .CLK(clock), .RSTB(n2735), .Q(reg3[24])
         );
  DFFARX1 \reg3_reg[25]  ( .D(n780), .CLK(clock), .RSTB(n2735), .Q(reg3[25]), 
        .QN(n2722) );
  DFFARX1 \reg3_reg[26]  ( .D(n779), .CLK(clock), .RSTB(n2735), .Q(reg3[26])
         );
  DFFARX1 \reg3_reg[27]  ( .D(n778), .CLK(clock), .RSTB(n2735), .Q(reg3[27]), 
        .QN(n2723) );
  DFFARX1 \reg3_reg[28]  ( .D(n777), .CLK(clock), .RSTB(n2735), .Q(reg3[28])
         );
  NOR2X0 U1087 ( .IN1(n1019), .IN2(n1020), .QN(n997) );
  NOR2X0 U1088 ( .IN1(n1017), .IN2(n1020), .QN(n998) );
  NOR2X0 U1089 ( .IN1(n1018), .IN2(n1019), .QN(n999) );
  NOR4X0 U1090 ( .IN1(n1846), .IN2(n2391), .IN3(n1842), .IN4(n2703), .QN(n1000) );
  INVX0 U1091 ( .INP(reset), .ZN(n2729) );
  INVX0 U1092 ( .INP(reset), .ZN(n2728) );
  INVX0 U1093 ( .INP(reset), .ZN(n2732) );
  INVX0 U1094 ( .INP(reset), .ZN(n2734) );
  INVX0 U1095 ( .INP(reset), .ZN(n2735) );
  INVX0 U1096 ( .INP(reset), .ZN(n2731) );
  INVX0 U1097 ( .INP(reset), .ZN(n2730) );
  INVX0 U1098 ( .INP(reset), .ZN(n2733) );
  NOR2X0 U1099 ( .IN1(IR[0]), .IN2(IR[1]), .QN(n1153) );
  NAND2X0 U1100 ( .IN1(n1153), .IN2(n2701), .QN(n1186) );
  OR3X1 U1101 ( .IN1(IR[3]), .IN2(IR[4]), .IN3(n1186), .Q(n1185) );
  OR3X1 U1102 ( .IN1(IR[5]), .IN2(IR[6]), .IN3(n1185), .Q(n1170) );
  OR3X1 U1103 ( .IN1(IR[7]), .IN2(IR[8]), .IN3(n1170), .Q(n1066) );
  OR3X1 U1104 ( .IN1(IR[9]), .IN2(IR[10]), .IN3(n1066), .Q(n1052) );
  OR3X1 U1105 ( .IN1(IR[11]), .IN2(IR[12]), .IN3(n1052), .Q(n1038) );
  OR3X1 U1106 ( .IN1(IR[13]), .IN2(IR[14]), .IN3(n1038), .Q(n1115) );
  OR3X1 U1107 ( .IN1(IR[15]), .IN2(IR[16]), .IN3(n1115), .Q(n1114) );
  OR3X1 U1108 ( .IN1(IR[17]), .IN2(IR[18]), .IN3(n1114), .Q(n1100) );
  NOR2X0 U1109 ( .IN1(IR[19]), .IN2(n1100), .QN(n1005) );
  NAND2X0 U1110 ( .IN1(n1005), .IN2(n2706), .QN(n1260) );
  NOR2X0 U1111 ( .IN1(IR[21]), .IN2(n1260), .QN(n1004) );
  NAND2X0 U1112 ( .IN1(n1004), .IN2(n2708), .QN(n1003) );
  NOR2X0 U1113 ( .IN1(IR[23]), .IN2(n1003), .QN(n1001) );
  NAND2X0 U1114 ( .IN1(n1001), .IN2(n2705), .QN(n1002) );
  NOR2X0 U1115 ( .IN1(IR[25]), .IN2(n1002), .QN(n1006) );
  MUX21X1 U1116 ( .IN1(n2707), .IN2(IR[26]), .S(n1006), .Q(n2650) );
  MUX21X1 U1117 ( .IN1(n2650), .IN2(IR[26]), .S(n2727), .Q(n1405) );
  MUX21X1 U1118 ( .IN1(n2705), .IN2(IR[24]), .S(n1001), .Q(n2648) );
  MUX21X1 U1119 ( .IN1(n2648), .IN2(IR[24]), .S(n2727), .Q(n1404) );
  MUX21X1 U1120 ( .IN1(IR[25]), .IN2(n2711), .S(n1002), .Q(n2649) );
  MUX21X1 U1121 ( .IN1(IR[25]), .IN2(n2649), .S(n2699), .Q(n1468) );
  AND3X1 U1122 ( .IN1(n1405), .IN2(n1404), .IN3(n1468), .Q(n1988) );
  MUX21X1 U1123 ( .IN1(IR[23]), .IN2(n2710), .S(n1003), .Q(n2647) );
  MUX21X1 U1124 ( .IN1(n2647), .IN2(IR[23]), .S(n2727), .Q(n1992) );
  INVX0 U1125 ( .INP(n1992), .ZN(n1987) );
  NAND2X0 U1126 ( .IN1(n1988), .IN2(n1987), .QN(n1994) );
  OR2X1 U1127 ( .IN1(n2703), .IN2(n1994), .Q(n2659) );
  INVX0 U1128 ( .INP(n2659), .ZN(n2736) );
  MUX21X1 U1129 ( .IN1(n2708), .IN2(IR[22]), .S(n1004), .Q(n2646) );
  MUX21X1 U1130 ( .IN1(IR[22]), .IN2(n2646), .S(n2699), .Q(n1831) );
  INVX0 U1131 ( .INP(n1831), .ZN(n2519) );
  MUX21X1 U1132 ( .IN1(n2706), .IN2(IR[20]), .S(n1005), .Q(n2644) );
  MUX21X1 U1133 ( .IN1(n2644), .IN2(IR[20]), .S(n2727), .Q(n1361) );
  INVX0 U1134 ( .INP(n1361), .ZN(n1363) );
  XNOR2X1 U1135 ( .IN1(IR[19]), .IN2(n1100), .Q(n1094) );
  NAND2X0 U1136 ( .IN1(n1006), .IN2(n2707), .QN(n1012) );
  NOR2X0 U1137 ( .IN1(IR[27]), .IN2(n1012), .QN(n1010) );
  NAND2X0 U1138 ( .IN1(n1010), .IN2(n2725), .QN(n1014) );
  NOR2X0 U1139 ( .IN1(IR[29]), .IN2(n1014), .QN(n1015) );
  NAND2X0 U1140 ( .IN1(n1015), .IN2(n2726), .QN(n1007) );
  NAND2X0 U1141 ( .IN1(n1007), .IN2(n2699), .QN(n2657) );
  NAND2X0 U1142 ( .IN1(IR[19]), .IN2(n2727), .QN(n1008) );
  OA21X1 U1143 ( .IN1(n1094), .IN2(n2657), .IN3(n1008), .Q(n2555) );
  INVX0 U1144 ( .INP(n2555), .ZN(n1265) );
  NAND2X0 U1145 ( .IN1(n2699), .IN2(n1115), .QN(n1009) );
  XNOR2X1 U1146 ( .IN1(IR[15]), .IN2(n1009), .Q(n2270) );
  MUX21X1 U1147 ( .IN1(n2725), .IN2(IR[28]), .S(n1010), .Q(n2653) );
  INVX0 U1148 ( .INP(n2653), .ZN(n1011) );
  MUX21X1 U1149 ( .IN1(n2725), .IN2(n1011), .S(n2699), .Q(n1996) );
  MUX21X1 U1150 ( .IN1(n2724), .IN2(IR[27]), .S(n1012), .Q(n2651) );
  NOR2X0 U1151 ( .IN1(n2651), .IN2(n2727), .QN(n1013) );
  AOI21X1 U1152 ( .IN1(n2727), .IN2(IR[27]), .IN3(n1013), .QN(n1989) );
  NAND2X0 U1153 ( .IN1(n1996), .IN2(n1989), .QN(n2520) );
  MUX21X1 U1154 ( .IN1(n2270), .IN2(datai[15]), .S(n2520), .Q(n2103) );
  INVX0 U1155 ( .INP(n2103), .ZN(n1543) );
  AOI21X1 U1156 ( .IN1(IR[29]), .IN2(n1014), .IN3(n1015), .QN(n2654) );
  MUX21X1 U1157 ( .IN1(IR[29]), .IN2(n2654), .S(n2699), .Q(n1019) );
  INVX0 U1158 ( .INP(n1019), .ZN(n1017) );
  MUX21X1 U1159 ( .IN1(n2726), .IN2(IR[30]), .S(n1015), .Q(n2655) );
  INVX0 U1160 ( .INP(n2655), .ZN(n1016) );
  MUX21X1 U1161 ( .IN1(n2726), .IN2(n1016), .S(n2699), .Q(n1018) );
  INVX0 U1162 ( .INP(n1018), .ZN(n1020) );
  NAND2X0 U1163 ( .IN1(n998), .IN2(reg1[15]), .QN(n1024) );
  NAND2X0 U1164 ( .IN1(n997), .IN2(reg0[15]), .QN(n1023) );
  NAND2X0 U1165 ( .IN1(n999), .IN2(reg2[15]), .QN(n1022) );
  NAND2X0 U1166 ( .IN1(n1020), .IN2(n1019), .QN(n1206) );
  NAND3X0 U1167 ( .IN1(reg3[3]), .IN2(reg3[4]), .IN3(reg3[5]), .QN(n1164) );
  INVX0 U1168 ( .INP(n1164), .ZN(n1174) );
  NAND2X0 U1169 ( .IN1(n1174), .IN2(reg3[6]), .QN(n1173) );
  NOR2X0 U1170 ( .IN1(n1173), .IN2(n2713), .QN(n1148) );
  NAND2X0 U1171 ( .IN1(n1148), .IN2(reg3[8]), .QN(n1069) );
  NOR2X0 U1172 ( .IN1(n1069), .IN2(n2714), .QN(n1061) );
  NAND2X0 U1173 ( .IN1(n1061), .IN2(reg3[10]), .QN(n1055) );
  NOR2X0 U1174 ( .IN1(n1055), .IN2(n2715), .QN(n1047) );
  NAND2X0 U1175 ( .IN1(n1047), .IN2(reg3[12]), .QN(n1041) );
  NOR2X0 U1176 ( .IN1(n1041), .IN2(n2716), .QN(n1033) );
  NAND2X0 U1177 ( .IN1(n1033), .IN2(reg3[14]), .QN(n1027) );
  NOR2X0 U1178 ( .IN1(n1027), .IN2(n2717), .QN(n1119) );
  AO21X1 U1179 ( .IN1(n1027), .IN2(n2717), .IN3(n1119), .Q(n1555) );
  OR2X1 U1180 ( .IN1(n1206), .IN2(n1555), .Q(n1021) );
  NAND4X0 U1181 ( .IN1(n1024), .IN2(n1023), .IN3(n1022), .IN4(n1021), .QN(
        n2675) );
  NAND2X0 U1182 ( .IN1(n1543), .IN2(n2675), .QN(n1545) );
  INVX0 U1183 ( .INP(n1115), .ZN(n1026) );
  OA21X1 U1184 ( .IN1(IR[13]), .IN2(n1038), .IN3(IR[14]), .Q(n1025) );
  NOR2X0 U1185 ( .IN1(n1026), .IN2(n1025), .QN(n1354) );
  MUX21X1 U1186 ( .IN1(IR[14]), .IN2(n1354), .S(n2699), .Q(n2278) );
  MUX21X1 U1187 ( .IN1(n2278), .IN2(datai[14]), .S(n2520), .Q(n2114) );
  INVX0 U1188 ( .INP(n2114), .ZN(n1574) );
  NAND2X0 U1189 ( .IN1(n998), .IN2(reg1[14]), .QN(n1031) );
  NAND2X0 U1190 ( .IN1(n997), .IN2(reg0[14]), .QN(n1030) );
  NAND2X0 U1191 ( .IN1(n999), .IN2(reg2[14]), .QN(n1029) );
  OA21X1 U1192 ( .IN1(n1033), .IN2(reg3[14]), .IN3(n1027), .Q(n2109) );
  INVX0 U1193 ( .INP(n1206), .ZN(n1201) );
  NAND2X0 U1194 ( .IN1(n2109), .IN2(n1201), .QN(n1028) );
  NAND4X0 U1195 ( .IN1(n1031), .IN2(n1030), .IN3(n1029), .IN4(n1028), .QN(
        n2674) );
  NAND2X0 U1196 ( .IN1(n1574), .IN2(n2674), .QN(n1563) );
  NAND2X0 U1197 ( .IN1(n2699), .IN2(n1038), .QN(n1032) );
  XNOR2X1 U1198 ( .IN1(IR[13]), .IN2(n1032), .Q(n2286) );
  MUX21X1 U1199 ( .IN1(n2286), .IN2(datai[13]), .S(n2520), .Q(n2125) );
  INVX0 U1200 ( .INP(n2125), .ZN(n1584) );
  NAND2X0 U1201 ( .IN1(n998), .IN2(reg1[13]), .QN(n1037) );
  NAND2X0 U1202 ( .IN1(n997), .IN2(reg0[13]), .QN(n1036) );
  NAND2X0 U1203 ( .IN1(n999), .IN2(reg2[13]), .QN(n1035) );
  AO21X1 U1204 ( .IN1(n1041), .IN2(n2716), .IN3(n1033), .Q(n1596) );
  OR2X1 U1205 ( .IN1(n1206), .IN2(n1596), .Q(n1034) );
  NAND4X0 U1206 ( .IN1(n1037), .IN2(n1036), .IN3(n1035), .IN4(n1034), .QN(
        n2673) );
  NAND2X0 U1207 ( .IN1(n1584), .IN2(n2673), .QN(n1586) );
  INVX0 U1208 ( .INP(n1038), .ZN(n1040) );
  OA21X1 U1209 ( .IN1(IR[11]), .IN2(n1052), .IN3(IR[12]), .Q(n1039) );
  NOR2X0 U1210 ( .IN1(n1040), .IN2(n1039), .QN(n1352) );
  MUX21X1 U1211 ( .IN1(IR[12]), .IN2(n1352), .S(n2699), .Q(n2294) );
  MUX21X1 U1212 ( .IN1(n2294), .IN2(datai[12]), .S(n2520), .Q(n2136) );
  INVX0 U1213 ( .INP(n2136), .ZN(n1615) );
  NAND2X0 U1214 ( .IN1(n998), .IN2(reg1[12]), .QN(n1045) );
  NAND2X0 U1215 ( .IN1(n997), .IN2(reg0[12]), .QN(n1044) );
  NAND2X0 U1216 ( .IN1(n999), .IN2(reg2[12]), .QN(n1043) );
  OA21X1 U1217 ( .IN1(n1047), .IN2(reg3[12]), .IN3(n1041), .Q(n2131) );
  NAND2X0 U1218 ( .IN1(n2131), .IN2(n1201), .QN(n1042) );
  NAND4X0 U1219 ( .IN1(n1045), .IN2(n1044), .IN3(n1043), .IN4(n1042), .QN(
        n2672) );
  NAND2X0 U1220 ( .IN1(n1615), .IN2(n2672), .QN(n1604) );
  AND4X1 U1221 ( .IN1(n1545), .IN2(n1563), .IN3(n1586), .IN4(n1604), .Q(n1074)
         );
  NAND2X0 U1222 ( .IN1(n2699), .IN2(n1052), .QN(n1046) );
  XNOR2X1 U1223 ( .IN1(IR[11]), .IN2(n1046), .Q(n2302) );
  MUX21X1 U1224 ( .IN1(n2302), .IN2(datai[11]), .S(n2520), .Q(n2147) );
  INVX0 U1225 ( .INP(n2147), .ZN(n1625) );
  NAND2X0 U1226 ( .IN1(n998), .IN2(reg1[11]), .QN(n1051) );
  NAND2X0 U1227 ( .IN1(n997), .IN2(reg0[11]), .QN(n1050) );
  NAND2X0 U1228 ( .IN1(n999), .IN2(reg2[11]), .QN(n1049) );
  AO21X1 U1229 ( .IN1(n1055), .IN2(n2715), .IN3(n1047), .Q(n1637) );
  OR2X1 U1230 ( .IN1(n1206), .IN2(n1637), .Q(n1048) );
  NAND4X0 U1231 ( .IN1(n1051), .IN2(n1050), .IN3(n1049), .IN4(n1048), .QN(
        n2671) );
  NAND2X0 U1232 ( .IN1(n1625), .IN2(n2671), .QN(n1627) );
  INVX0 U1233 ( .INP(n1052), .ZN(n1054) );
  OA21X1 U1234 ( .IN1(IR[9]), .IN2(n1066), .IN3(IR[10]), .Q(n1053) );
  NOR2X0 U1235 ( .IN1(n1054), .IN2(n1053), .QN(n1350) );
  MUX21X1 U1236 ( .IN1(IR[10]), .IN2(n1350), .S(n2699), .Q(n2310) );
  MUX21X1 U1237 ( .IN1(n2310), .IN2(datai[10]), .S(n2520), .Q(n2158) );
  INVX0 U1238 ( .INP(n2158), .ZN(n1656) );
  NAND2X0 U1239 ( .IN1(n998), .IN2(reg1[10]), .QN(n1059) );
  NAND2X0 U1240 ( .IN1(n997), .IN2(reg0[10]), .QN(n1058) );
  NAND2X0 U1241 ( .IN1(n999), .IN2(reg2[10]), .QN(n1057) );
  OA21X1 U1242 ( .IN1(n1061), .IN2(reg3[10]), .IN3(n1055), .Q(n2153) );
  NAND2X0 U1243 ( .IN1(n2153), .IN2(n1201), .QN(n1056) );
  NAND4X0 U1244 ( .IN1(n1059), .IN2(n1058), .IN3(n1057), .IN4(n1056), .QN(
        n2670) );
  NAND2X0 U1245 ( .IN1(n1656), .IN2(n2670), .QN(n1645) );
  NAND2X0 U1246 ( .IN1(n2699), .IN2(n1066), .QN(n1060) );
  XNOR2X1 U1247 ( .IN1(IR[9]), .IN2(n1060), .Q(n2318) );
  MUX21X1 U1248 ( .IN1(n2318), .IN2(datai[9]), .S(n2520), .Q(n2169) );
  INVX0 U1249 ( .INP(n2169), .ZN(n1666) );
  NAND2X0 U1250 ( .IN1(n998), .IN2(reg1[9]), .QN(n1065) );
  NAND2X0 U1251 ( .IN1(n997), .IN2(reg0[9]), .QN(n1064) );
  NAND2X0 U1252 ( .IN1(n999), .IN2(reg2[9]), .QN(n1063) );
  AO21X1 U1253 ( .IN1(n1069), .IN2(n2714), .IN3(n1061), .Q(n1678) );
  OR2X1 U1254 ( .IN1(n1206), .IN2(n1678), .Q(n1062) );
  NAND4X0 U1255 ( .IN1(n1065), .IN2(n1064), .IN3(n1063), .IN4(n1062), .QN(
        n2669) );
  NAND2X0 U1256 ( .IN1(n1666), .IN2(n2669), .QN(n1668) );
  AND3X1 U1257 ( .IN1(n1627), .IN2(n1645), .IN3(n1668), .Q(n1221) );
  INVX0 U1258 ( .INP(n1066), .ZN(n1068) );
  OA21X1 U1259 ( .IN1(IR[7]), .IN2(n1170), .IN3(IR[8]), .Q(n1067) );
  NOR2X0 U1260 ( .IN1(n1068), .IN2(n1067), .QN(n1348) );
  MUX21X1 U1261 ( .IN1(IR[8]), .IN2(n1348), .S(n2699), .Q(n2326) );
  MUX21X1 U1262 ( .IN1(n2326), .IN2(datai[8]), .S(n2520), .Q(n2180) );
  INVX0 U1263 ( .INP(n2180), .ZN(n1697) );
  NAND2X0 U1264 ( .IN1(n998), .IN2(reg1[8]), .QN(n1073) );
  NAND2X0 U1265 ( .IN1(n997), .IN2(reg0[8]), .QN(n1072) );
  NAND2X0 U1266 ( .IN1(n999), .IN2(reg2[8]), .QN(n1071) );
  OA21X1 U1267 ( .IN1(n1148), .IN2(reg3[8]), .IN3(n1069), .Q(n2175) );
  NAND2X0 U1268 ( .IN1(n2175), .IN2(n1201), .QN(n1070) );
  NAND4X0 U1269 ( .IN1(n1073), .IN2(n1072), .IN3(n1071), .IN4(n1070), .QN(
        n2668) );
  NAND2X0 U1270 ( .IN1(n1697), .IN2(n2668), .QN(n1684) );
  NAND3X0 U1271 ( .IN1(n1074), .IN2(n1221), .IN3(n1684), .QN(n1225) );
  AND2X1 U1272 ( .IN1(datai[23]), .IN2(n2520), .Q(n2036) );
  INVX0 U1273 ( .INP(n2036), .ZN(n1426) );
  NAND2X0 U1274 ( .IN1(n998), .IN2(reg1[23]), .QN(n1078) );
  NAND2X0 U1275 ( .IN1(n997), .IN2(reg0[23]), .QN(n1077) );
  NAND2X0 U1276 ( .IN1(n999), .IN2(reg2[23]), .QN(n1076) );
  NAND2X0 U1277 ( .IN1(n1119), .IN2(reg3[16]), .QN(n1118) );
  NOR2X0 U1278 ( .IN1(n1118), .IN2(n2718), .QN(n1109) );
  NAND2X0 U1279 ( .IN1(n1109), .IN2(reg3[18]), .QN(n1103) );
  NOR2X0 U1280 ( .IN1(n1103), .IN2(n2719), .QN(n1095) );
  NAND2X0 U1281 ( .IN1(n1095), .IN2(reg3[20]), .QN(n1089) );
  NOR2X0 U1282 ( .IN1(n1089), .IN2(n2720), .QN(n1084) );
  NAND2X0 U1283 ( .IN1(n1084), .IN2(reg3[22]), .QN(n1079) );
  NOR2X0 U1284 ( .IN1(n1079), .IN2(n2721), .QN(n1142) );
  AO21X1 U1285 ( .IN1(n1079), .IN2(n2721), .IN3(n1142), .Q(n2025) );
  OR2X1 U1286 ( .IN1(n1206), .IN2(n2025), .Q(n1075) );
  NAND4X0 U1287 ( .IN1(n1078), .IN2(n1077), .IN3(n1076), .IN4(n1075), .QN(
        n2684) );
  NAND2X0 U1288 ( .IN1(n1426), .IN2(n2684), .QN(n1428) );
  AND2X1 U1289 ( .IN1(datai[22]), .IN2(n2520), .Q(n2429) );
  INVX0 U1290 ( .INP(n2429), .ZN(n2430) );
  NAND2X0 U1291 ( .IN1(n998), .IN2(reg1[22]), .QN(n1083) );
  NAND2X0 U1292 ( .IN1(n997), .IN2(reg0[22]), .QN(n1082) );
  NAND2X0 U1293 ( .IN1(n999), .IN2(reg2[22]), .QN(n1081) );
  OA21X1 U1294 ( .IN1(n1084), .IN2(reg3[22]), .IN3(n1079), .Q(n2432) );
  NAND2X0 U1295 ( .IN1(n2432), .IN2(n1201), .QN(n1080) );
  NAND4X0 U1296 ( .IN1(n1083), .IN2(n1082), .IN3(n1081), .IN4(n1080), .QN(
        n2683) );
  NAND2X0 U1297 ( .IN1(n2430), .IN2(n2683), .QN(n2417) );
  AND2X1 U1298 ( .IN1(datai[21]), .IN2(n2520), .Q(n2048) );
  INVX0 U1299 ( .INP(n2048), .ZN(n1440) );
  NAND2X0 U1300 ( .IN1(n998), .IN2(reg1[21]), .QN(n1088) );
  NAND2X0 U1301 ( .IN1(n997), .IN2(reg0[21]), .QN(n1087) );
  NAND2X0 U1302 ( .IN1(n999), .IN2(reg2[21]), .QN(n1086) );
  AO21X1 U1303 ( .IN1(n1089), .IN2(n2720), .IN3(n1084), .Q(n2037) );
  OR2X1 U1304 ( .IN1(n1206), .IN2(n2037), .Q(n1085) );
  NAND4X0 U1305 ( .IN1(n1088), .IN2(n1087), .IN3(n1086), .IN4(n1085), .QN(
        n2681) );
  NAND2X0 U1306 ( .IN1(n1440), .IN2(n2681), .QN(n1442) );
  AND2X1 U1307 ( .IN1(datai[20]), .IN2(n2520), .Q(n2406) );
  INVX0 U1308 ( .INP(n2406), .ZN(n2407) );
  NAND2X0 U1309 ( .IN1(n998), .IN2(reg1[20]), .QN(n1093) );
  NAND2X0 U1310 ( .IN1(n997), .IN2(reg0[20]), .QN(n1092) );
  NAND2X0 U1311 ( .IN1(n999), .IN2(reg2[20]), .QN(n1091) );
  OA21X1 U1312 ( .IN1(n1095), .IN2(reg3[20]), .IN3(n1089), .Q(n2409) );
  NAND2X0 U1313 ( .IN1(n2409), .IN2(n1201), .QN(n1090) );
  NAND4X0 U1314 ( .IN1(n1093), .IN2(n1092), .IN3(n1091), .IN4(n1090), .QN(
        n2680) );
  NAND2X0 U1315 ( .IN1(n2407), .IN2(n2680), .QN(n2394) );
  AND4X1 U1316 ( .IN1(n1428), .IN2(n2417), .IN3(n1442), .IN4(n2394), .Q(n1124)
         );
  INVX0 U1317 ( .INP(n1094), .ZN(n1360) );
  MUX21X1 U1318 ( .IN1(IR[19]), .IN2(n1360), .S(n2699), .Q(n2238) );
  MUX21X1 U1319 ( .IN1(n2238), .IN2(datai[19]), .S(n2520), .Q(n2059) );
  INVX0 U1320 ( .INP(n2059), .ZN(n1454) );
  NAND2X0 U1321 ( .IN1(n998), .IN2(reg1[19]), .QN(n1099) );
  NAND2X0 U1322 ( .IN1(n997), .IN2(reg0[19]), .QN(n1098) );
  NAND2X0 U1323 ( .IN1(n999), .IN2(reg2[19]), .QN(n1097) );
  AO21X1 U1324 ( .IN1(n1103), .IN2(n2719), .IN3(n1095), .Q(n1471) );
  OR2X1 U1325 ( .IN1(n1206), .IN2(n1471), .Q(n1096) );
  NAND4X0 U1326 ( .IN1(n1099), .IN2(n1098), .IN3(n1097), .IN4(n1096), .QN(
        n2679) );
  NAND2X0 U1327 ( .IN1(n1454), .IN2(n2679), .QN(n1456) );
  INVX0 U1328 ( .INP(n1100), .ZN(n1102) );
  OA21X1 U1329 ( .IN1(IR[17]), .IN2(n1114), .IN3(IR[18]), .Q(n1101) );
  NOR2X0 U1330 ( .IN1(n1102), .IN2(n1101), .QN(n1358) );
  MUX21X1 U1331 ( .IN1(IR[18]), .IN2(n1358), .S(n2699), .Q(n2246) );
  MUX21X1 U1332 ( .IN1(n2246), .IN2(datai[18]), .S(n2520), .Q(n2070) );
  INVX0 U1333 ( .INP(n2070), .ZN(n1492) );
  NAND2X0 U1334 ( .IN1(n998), .IN2(reg1[18]), .QN(n1107) );
  NAND2X0 U1335 ( .IN1(n997), .IN2(reg0[18]), .QN(n1106) );
  NAND2X0 U1336 ( .IN1(n999), .IN2(reg2[18]), .QN(n1105) );
  OA21X1 U1337 ( .IN1(n1109), .IN2(reg3[18]), .IN3(n1103), .Q(n2065) );
  NAND2X0 U1338 ( .IN1(n2065), .IN2(n1201), .QN(n1104) );
  NAND4X0 U1339 ( .IN1(n1107), .IN2(n1106), .IN3(n1105), .IN4(n1104), .QN(
        n2678) );
  NAND2X0 U1340 ( .IN1(n1492), .IN2(n2678), .QN(n1481) );
  NAND2X0 U1341 ( .IN1(n2699), .IN2(n1114), .QN(n1108) );
  XNOR2X1 U1342 ( .IN1(IR[17]), .IN2(n1108), .Q(n2254) );
  MUX21X1 U1343 ( .IN1(n2254), .IN2(datai[17]), .S(n2520), .Q(n2081) );
  INVX0 U1344 ( .INP(n2081), .ZN(n1502) );
  NAND2X0 U1345 ( .IN1(n998), .IN2(reg1[17]), .QN(n1113) );
  NAND2X0 U1346 ( .IN1(n997), .IN2(reg0[17]), .QN(n1112) );
  NAND2X0 U1347 ( .IN1(n999), .IN2(reg2[17]), .QN(n1111) );
  AO21X1 U1348 ( .IN1(n1118), .IN2(n2718), .IN3(n1109), .Q(n1514) );
  OR2X1 U1349 ( .IN1(n1206), .IN2(n1514), .Q(n1110) );
  NAND4X0 U1350 ( .IN1(n1113), .IN2(n1112), .IN3(n1111), .IN4(n1110), .QN(
        n2677) );
  NAND2X0 U1351 ( .IN1(n1502), .IN2(n2677), .QN(n1504) );
  AND3X1 U1352 ( .IN1(n1456), .IN2(n1481), .IN3(n1504), .Q(n1239) );
  INVX0 U1353 ( .INP(n1114), .ZN(n1117) );
  OA21X1 U1354 ( .IN1(IR[15]), .IN2(n1115), .IN3(IR[16]), .Q(n1116) );
  NOR2X0 U1355 ( .IN1(n1117), .IN2(n1116), .QN(n1356) );
  MUX21X1 U1356 ( .IN1(IR[16]), .IN2(n1356), .S(n2699), .Q(n2262) );
  MUX21X1 U1357 ( .IN1(n2262), .IN2(datai[16]), .S(n2520), .Q(n2092) );
  INVX0 U1358 ( .INP(n2092), .ZN(n1533) );
  NAND2X0 U1359 ( .IN1(n998), .IN2(reg1[16]), .QN(n1123) );
  NAND2X0 U1360 ( .IN1(n997), .IN2(reg0[16]), .QN(n1122) );
  NAND2X0 U1361 ( .IN1(n999), .IN2(reg2[16]), .QN(n1121) );
  OA21X1 U1362 ( .IN1(n1119), .IN2(reg3[16]), .IN3(n1118), .Q(n2087) );
  NAND2X0 U1363 ( .IN1(n2087), .IN2(n1201), .QN(n1120) );
  NAND4X0 U1364 ( .IN1(n1123), .IN2(n1122), .IN3(n1121), .IN4(n1120), .QN(
        n2676) );
  NAND2X0 U1365 ( .IN1(n1533), .IN2(n2676), .QN(n1522) );
  NAND3X0 U1366 ( .IN1(n1124), .IN2(n1239), .IN3(n1522), .QN(n1233) );
  NOR2X0 U1367 ( .IN1(n1225), .IN2(n1233), .QN(n1215) );
  INVX0 U1368 ( .INP(n2668), .ZN(n1918) );
  NAND2X0 U1369 ( .IN1(n2180), .IN2(n1918), .QN(n1683) );
  INVX0 U1370 ( .INP(n1683), .ZN(n1374) );
  NOR2X0 U1371 ( .IN1(n1543), .IN2(n2675), .QN(n1381) );
  INVX0 U1372 ( .INP(n1381), .ZN(n1544) );
  INVX0 U1373 ( .INP(n2674), .ZN(n1912) );
  NAND2X0 U1374 ( .IN1(n2114), .IN2(n1912), .QN(n1562) );
  NOR2X0 U1375 ( .IN1(n1584), .IN2(n2673), .QN(n1379) );
  INVX0 U1376 ( .INP(n1379), .ZN(n1585) );
  INVX0 U1377 ( .INP(n2672), .ZN(n1914) );
  NAND2X0 U1378 ( .IN1(n2136), .IN2(n1914), .QN(n1603) );
  NAND4X0 U1379 ( .IN1(n1544), .IN2(n1562), .IN3(n1585), .IN4(n1603), .QN(
        n1125) );
  NOR2X0 U1380 ( .IN1(n1625), .IN2(n2671), .QN(n1377) );
  INVX0 U1381 ( .INP(n1377), .ZN(n1626) );
  INVX0 U1382 ( .INP(n2670), .ZN(n1916) );
  NAND2X0 U1383 ( .IN1(n2158), .IN2(n1916), .QN(n1644) );
  NOR2X0 U1384 ( .IN1(n1666), .IN2(n2669), .QN(n1375) );
  INVX0 U1385 ( .INP(n1375), .ZN(n1667) );
  NAND3X0 U1386 ( .IN1(n1626), .IN2(n1644), .IN3(n1667), .QN(n1272) );
  NOR3X0 U1387 ( .IN1(n1374), .IN2(n1125), .IN3(n1272), .QN(n1300) );
  INVX0 U1388 ( .INP(n2676), .ZN(n1910) );
  NAND2X0 U1389 ( .IN1(n2092), .IN2(n1910), .QN(n1521) );
  INVX0 U1390 ( .INP(n1521), .ZN(n1382) );
  NOR2X0 U1391 ( .IN1(n1426), .IN2(n2684), .QN(n1389) );
  INVX0 U1392 ( .INP(n1389), .ZN(n1427) );
  INVX0 U1393 ( .INP(n2683), .ZN(n1934) );
  NAND2X0 U1394 ( .IN1(n2429), .IN2(n1934), .QN(n2416) );
  NOR2X0 U1395 ( .IN1(n1440), .IN2(n2681), .QN(n1387) );
  INVX0 U1396 ( .INP(n1387), .ZN(n1441) );
  INVX0 U1397 ( .INP(n2680), .ZN(n1905) );
  NAND2X0 U1398 ( .IN1(n2406), .IN2(n1905), .QN(n2393) );
  NAND4X0 U1399 ( .IN1(n1427), .IN2(n2416), .IN3(n1441), .IN4(n2393), .QN(
        n1126) );
  NOR2X0 U1400 ( .IN1(n1454), .IN2(n2679), .QN(n1385) );
  INVX0 U1401 ( .INP(n1385), .ZN(n1455) );
  INVX0 U1402 ( .INP(n2678), .ZN(n1907) );
  NAND2X0 U1403 ( .IN1(n2070), .IN2(n1907), .QN(n1480) );
  NOR2X0 U1404 ( .IN1(n1502), .IN2(n2677), .QN(n1383) );
  INVX0 U1405 ( .INP(n1383), .ZN(n1503) );
  NAND3X0 U1406 ( .IN1(n1455), .IN2(n1480), .IN3(n1503), .QN(n1301) );
  NOR3X0 U1407 ( .IN1(n1382), .IN2(n1126), .IN3(n1301), .QN(n1311) );
  AND2X1 U1408 ( .IN1(datai[27]), .IN2(n2520), .Q(n2492) );
  INVX0 U1409 ( .INP(n2492), .ZN(n1365) );
  NAND2X0 U1410 ( .IN1(n998), .IN2(reg1[27]), .QN(n1130) );
  NAND2X0 U1411 ( .IN1(n997), .IN2(reg0[27]), .QN(n1129) );
  NAND2X0 U1412 ( .IN1(n999), .IN2(reg2[27]), .QN(n1128) );
  NAND2X0 U1413 ( .IN1(n1142), .IN2(reg3[24]), .QN(n1141) );
  NOR2X0 U1414 ( .IN1(n1141), .IN2(n2722), .QN(n1136) );
  NAND2X0 U1415 ( .IN1(n1136), .IN2(reg3[26]), .QN(n1131) );
  NOR2X0 U1416 ( .IN1(n1131), .IN2(n2723), .QN(n1200) );
  AO21X1 U1417 ( .IN1(n1131), .IN2(n2723), .IN3(n1200), .Q(n2002) );
  OR2X1 U1418 ( .IN1(n1206), .IN2(n2002), .Q(n1127) );
  NAND4X0 U1419 ( .IN1(n1130), .IN2(n1129), .IN3(n1128), .IN4(n1127), .QN(
        n2688) );
  NAND2X0 U1420 ( .IN1(n1365), .IN2(n2688), .QN(n2486) );
  AND2X1 U1421 ( .IN1(datai[26]), .IN2(n2520), .Q(n2475) );
  INVX0 U1422 ( .INP(n2475), .ZN(n2476) );
  NAND2X0 U1423 ( .IN1(n998), .IN2(reg1[26]), .QN(n1135) );
  NAND2X0 U1424 ( .IN1(n997), .IN2(reg0[26]), .QN(n1134) );
  NAND2X0 U1425 ( .IN1(n999), .IN2(reg2[26]), .QN(n1133) );
  OA21X1 U1426 ( .IN1(n1136), .IN2(reg3[26]), .IN3(n1131), .Q(n2478) );
  NAND2X0 U1427 ( .IN1(n2478), .IN2(n1201), .QN(n1132) );
  NAND4X0 U1428 ( .IN1(n1135), .IN2(n1134), .IN3(n1133), .IN4(n1132), .QN(
        n2687) );
  NAND2X0 U1429 ( .IN1(n2476), .IN2(n2687), .QN(n2463) );
  AND2X1 U1430 ( .IN1(datai[25]), .IN2(n2520), .Q(n2024) );
  INVX0 U1431 ( .INP(n2024), .ZN(n1412) );
  NAND2X0 U1432 ( .IN1(n998), .IN2(reg1[25]), .QN(n1140) );
  NAND2X0 U1433 ( .IN1(n997), .IN2(reg0[25]), .QN(n1139) );
  NAND2X0 U1434 ( .IN1(n999), .IN2(reg2[25]), .QN(n1138) );
  AO21X1 U1435 ( .IN1(n1141), .IN2(n2722), .IN3(n1136), .Q(n2013) );
  OR2X1 U1436 ( .IN1(n1206), .IN2(n2013), .Q(n1137) );
  NAND4X0 U1437 ( .IN1(n1140), .IN2(n1139), .IN3(n1138), .IN4(n1137), .QN(
        n2686) );
  NAND2X0 U1438 ( .IN1(n1412), .IN2(n2686), .QN(n1414) );
  AND2X1 U1439 ( .IN1(datai[24]), .IN2(n2520), .Q(n2452) );
  INVX0 U1440 ( .INP(n2452), .ZN(n2453) );
  NAND2X0 U1441 ( .IN1(n998), .IN2(reg1[24]), .QN(n1146) );
  NAND2X0 U1442 ( .IN1(n997), .IN2(reg0[24]), .QN(n1145) );
  NAND2X0 U1443 ( .IN1(n999), .IN2(reg2[24]), .QN(n1144) );
  OA21X1 U1444 ( .IN1(n1142), .IN2(reg3[24]), .IN3(n1141), .Q(n2455) );
  NAND2X0 U1445 ( .IN1(n2455), .IN2(n1201), .QN(n1143) );
  NAND4X0 U1446 ( .IN1(n1146), .IN2(n1145), .IN3(n1144), .IN4(n1143), .QN(
        n2685) );
  NAND2X0 U1447 ( .IN1(n2453), .IN2(n2685), .QN(n2440) );
  NAND4X0 U1448 ( .IN1(n2486), .IN2(n2463), .IN3(n1414), .IN4(n2440), .QN(
        n1248) );
  NAND2X0 U1449 ( .IN1(n2699), .IN2(n1170), .QN(n1147) );
  XNOR2X1 U1450 ( .IN1(IR[7]), .IN2(n1147), .Q(n2334) );
  MUX21X1 U1451 ( .IN1(n2334), .IN2(datai[7]), .S(n2520), .Q(n2191) );
  INVX0 U1452 ( .INP(n2191), .ZN(n1707) );
  NAND2X0 U1453 ( .IN1(n998), .IN2(reg1[7]), .QN(n1152) );
  NAND2X0 U1454 ( .IN1(n997), .IN2(reg0[7]), .QN(n1151) );
  NAND2X0 U1455 ( .IN1(n999), .IN2(reg2[7]), .QN(n1150) );
  AO21X1 U1456 ( .IN1(n1173), .IN2(n2713), .IN3(n1148), .Q(n1717) );
  OR2X1 U1457 ( .IN1(n1206), .IN2(n1717), .Q(n1149) );
  NAND4X0 U1458 ( .IN1(n1152), .IN2(n1151), .IN3(n1150), .IN4(n1149), .QN(
        n2667) );
  NAND2X0 U1459 ( .IN1(n1707), .IN2(n2667), .QN(n1372) );
  NOR2X0 U1460 ( .IN1(n1707), .IN2(n2667), .QN(n1373) );
  INVX0 U1461 ( .INP(n1373), .ZN(n1295) );
  NAND2X0 U1462 ( .IN1(n1372), .IN2(n1295), .QN(n1710) );
  INVX0 U1463 ( .INP(n1710), .ZN(n1712) );
  OA21X1 U1464 ( .IN1(n1153), .IN2(n2701), .IN3(n1186), .Q(n1342) );
  MUX21X1 U1465 ( .IN1(IR[2]), .IN2(n1342), .S(n2699), .Q(n2371) );
  MUX21X1 U1466 ( .IN1(n2371), .IN2(datai[2]), .S(n2520), .Q(n1859) );
  NAND2X0 U1467 ( .IN1(n998), .IN2(reg1[2]), .QN(n1157) );
  NAND2X0 U1468 ( .IN1(n997), .IN2(reg0[2]), .QN(n1156) );
  NAND2X0 U1469 ( .IN1(n999), .IN2(reg2[2]), .QN(n1155) );
  NAND2X0 U1470 ( .IN1(reg3[2]), .IN2(n1201), .QN(n1154) );
  NAND4X0 U1471 ( .IN1(n1157), .IN2(n1156), .IN3(n1155), .IN4(n1154), .QN(
        n2662) );
  INVX0 U1472 ( .INP(n2662), .ZN(n1858) );
  NAND2X0 U1473 ( .IN1(n1859), .IN2(n1858), .QN(n1798) );
  INVX0 U1474 ( .INP(n1798), .ZN(n1226) );
  NAND2X0 U1475 ( .IN1(n2699), .IN2(n1186), .QN(n1158) );
  XNOR2X1 U1476 ( .IN1(IR[3]), .IN2(n1158), .Q(n2358) );
  MUX21X1 U1477 ( .IN1(n2358), .IN2(datai[3]), .S(n2520), .Q(n1901) );
  INVX0 U1478 ( .INP(n1901), .ZN(n1780) );
  NAND2X0 U1479 ( .IN1(n998), .IN2(reg1[3]), .QN(n1162) );
  NAND2X0 U1480 ( .IN1(n997), .IN2(reg0[3]), .QN(n1161) );
  NAND2X0 U1481 ( .IN1(n999), .IN2(reg2[3]), .QN(n1160) );
  NAND2X0 U1482 ( .IN1(n1201), .IN2(n2698), .QN(n1159) );
  NAND4X0 U1483 ( .IN1(n1162), .IN2(n1161), .IN3(n1160), .IN4(n1159), .QN(
        n2663) );
  NOR2X0 U1484 ( .IN1(n1780), .IN2(n2663), .QN(n1281) );
  NAND2X0 U1485 ( .IN1(n2699), .IN2(n1185), .QN(n1163) );
  XNOR2X1 U1486 ( .IN1(IR[5]), .IN2(n1163), .Q(n2350) );
  MUX21X1 U1487 ( .IN1(n2350), .IN2(datai[5]), .S(n2520), .Q(n2214) );
  INVX0 U1488 ( .INP(n2214), .ZN(n1744) );
  NAND2X0 U1489 ( .IN1(n998), .IN2(reg1[5]), .QN(n1169) );
  NAND2X0 U1490 ( .IN1(reg3[3]), .IN2(reg3[4]), .QN(n1189) );
  INVX0 U1491 ( .INP(n1189), .ZN(n1165) );
  OA21X1 U1492 ( .IN1(n1165), .IN2(reg3[5]), .IN3(n1164), .Q(n2203) );
  NAND2X0 U1493 ( .IN1(n2203), .IN2(n1201), .QN(n1168) );
  NAND2X0 U1494 ( .IN1(n999), .IN2(reg2[5]), .QN(n1167) );
  NAND2X0 U1495 ( .IN1(n997), .IN2(reg0[5]), .QN(n1166) );
  NAND4X0 U1496 ( .IN1(n1169), .IN2(n1168), .IN3(n1167), .IN4(n1166), .QN(
        n2665) );
  NAND2X0 U1497 ( .IN1(n1744), .IN2(n2665), .QN(n1368) );
  INVX0 U1498 ( .INP(n1368), .ZN(n1280) );
  NOR2X0 U1499 ( .IN1(n1744), .IN2(n2665), .QN(n1369) );
  NOR2X0 U1500 ( .IN1(n1280), .IN2(n1369), .QN(n1749) );
  INVX0 U1501 ( .INP(n1749), .ZN(n1747) );
  INVX0 U1502 ( .INP(n1170), .ZN(n1172) );
  OA21X1 U1503 ( .IN1(IR[5]), .IN2(n1185), .IN3(IR[6]), .Q(n1171) );
  NOR2X0 U1504 ( .IN1(n1172), .IN2(n1171), .QN(n1346) );
  MUX21X1 U1505 ( .IN1(IR[6]), .IN2(n1346), .S(n2699), .Q(n2342) );
  MUX21X1 U1506 ( .IN1(n2342), .IN2(datai[6]), .S(n2520), .Q(n2202) );
  INVX0 U1507 ( .INP(n2202), .ZN(n1734) );
  NAND2X0 U1508 ( .IN1(n998), .IN2(reg1[6]), .QN(n1178) );
  NAND2X0 U1509 ( .IN1(n997), .IN2(reg0[6]), .QN(n1177) );
  NAND2X0 U1510 ( .IN1(n999), .IN2(reg2[6]), .QN(n1176) );
  OA21X1 U1511 ( .IN1(n1174), .IN2(reg3[6]), .IN3(n1173), .Q(n2197) );
  NAND2X0 U1512 ( .IN1(n2197), .IN2(n1201), .QN(n1175) );
  NAND4X0 U1513 ( .IN1(n1178), .IN2(n1177), .IN3(n1176), .IN4(n1175), .QN(
        n2666) );
  NAND2X0 U1514 ( .IN1(n1734), .IN2(n2666), .QN(n1370) );
  INVX0 U1515 ( .INP(n2666), .ZN(n1920) );
  NAND2X0 U1516 ( .IN1(n2202), .IN2(n1920), .QN(n1293) );
  NAND2X0 U1517 ( .IN1(n1370), .IN2(n1293), .QN(n1726) );
  INVX0 U1518 ( .INP(n1726), .ZN(n1728) );
  NAND2X0 U1519 ( .IN1(n2699), .IN2(IR[0]), .QN(n1179) );
  XNOR2X1 U1520 ( .IN1(IR[1]), .IN2(n1179), .Q(n2373) );
  MUX21X1 U1521 ( .IN1(n2373), .IN2(datai[1]), .S(n2520), .Q(n1837) );
  INVX0 U1522 ( .INP(n1837), .ZN(n1816) );
  NAND2X0 U1523 ( .IN1(reg1[1]), .IN2(n998), .QN(n1183) );
  NAND2X0 U1524 ( .IN1(reg3[1]), .IN2(n1201), .QN(n1182) );
  NAND2X0 U1525 ( .IN1(reg2[1]), .IN2(n999), .QN(n1181) );
  NAND2X0 U1526 ( .IN1(n997), .IN2(reg0[1]), .QN(n1180) );
  NAND4X0 U1527 ( .IN1(n1183), .IN2(n1182), .IN3(n1181), .IN4(n1180), .QN(
        n2661) );
  NAND2X0 U1528 ( .IN1(n1816), .IN2(n2661), .QN(n1285) );
  NOR2X0 U1529 ( .IN1(n1816), .IN2(n2661), .QN(n1283) );
  INVX0 U1530 ( .INP(n1283), .ZN(n1184) );
  NAND2X0 U1531 ( .IN1(n1285), .IN2(n1184), .QN(n1821) );
  INVX0 U1532 ( .INP(n1821), .ZN(n1819) );
  INVX0 U1533 ( .INP(n1185), .ZN(n1188) );
  OA21X1 U1534 ( .IN1(IR[3]), .IN2(n1186), .IN3(IR[4]), .Q(n1187) );
  NOR2X0 U1535 ( .IN1(n1188), .IN2(n1187), .QN(n1344) );
  MUX21X1 U1536 ( .IN1(IR[4]), .IN2(n1344), .S(n2699), .Q(n2231) );
  MUX21X1 U1537 ( .IN1(n2231), .IN2(datai[4]), .S(n2520), .Q(n2228) );
  NAND2X0 U1538 ( .IN1(n998), .IN2(reg1[4]), .QN(n1193) );
  NAND2X0 U1539 ( .IN1(n997), .IN2(reg0[4]), .QN(n1192) );
  NAND2X0 U1540 ( .IN1(n999), .IN2(reg2[4]), .QN(n1191) );
  OA21X1 U1541 ( .IN1(reg3[3]), .IN2(reg3[4]), .IN3(n1189), .Q(n2221) );
  NAND2X0 U1542 ( .IN1(n2221), .IN2(n1201), .QN(n1190) );
  NAND4X0 U1543 ( .IN1(n1193), .IN2(n1192), .IN3(n1191), .IN4(n1190), .QN(
        n2664) );
  INVX0 U1544 ( .INP(n2664), .ZN(n1922) );
  NOR2X0 U1545 ( .IN1(n2228), .IN2(n1922), .QN(n1279) );
  INVX0 U1546 ( .INP(n2228), .ZN(n1770) );
  NOR2X0 U1547 ( .IN1(n1770), .IN2(n2664), .QN(n1367) );
  NOR2X0 U1548 ( .IN1(n1279), .IN2(n1367), .QN(n1764) );
  MUX21X1 U1549 ( .IN1(IR[0]), .IN2(datai[0]), .S(n2520), .Q(n1885) );
  NAND2X0 U1550 ( .IN1(n998), .IN2(reg1[0]), .QN(n1197) );
  NAND2X0 U1551 ( .IN1(n997), .IN2(reg0[0]), .QN(n1196) );
  NAND2X0 U1552 ( .IN1(n999), .IN2(reg2[0]), .QN(n1195) );
  NAND2X0 U1553 ( .IN1(reg3[0]), .IN2(n1201), .QN(n1194) );
  NAND4X0 U1554 ( .IN1(n1197), .IN2(n1196), .IN3(n1195), .IN4(n1194), .QN(
        n2660) );
  INVX0 U1555 ( .INP(n2660), .ZN(n1838) );
  NAND2X0 U1556 ( .IN1(n1885), .IN2(n1838), .QN(n1820) );
  INVX0 U1557 ( .INP(n1885), .ZN(n2579) );
  NAND2X0 U1558 ( .IN1(n2660), .IN2(n2579), .QN(n1284) );
  AND2X1 U1559 ( .IN1(n1820), .IN2(n1284), .Q(n1873) );
  NAND4X0 U1560 ( .IN1(n1728), .IN2(n1819), .IN3(n1764), .IN4(n1873), .QN(
        n1198) );
  NOR4X0 U1561 ( .IN1(n1226), .IN2(n1281), .IN3(n1747), .IN4(n1198), .QN(n1199) );
  NAND2X0 U1562 ( .IN1(n1780), .IN2(n2663), .QN(n1782) );
  INVX0 U1563 ( .INP(n1859), .ZN(n1810) );
  NAND2X0 U1564 ( .IN1(n1810), .IN2(n2662), .QN(n1799) );
  NAND4X0 U1565 ( .IN1(n1712), .IN2(n1199), .IN3(n1782), .IN4(n1799), .QN(
        n1213) );
  AND2X1 U1566 ( .IN1(datai[28]), .IN2(n2520), .Q(n2535) );
  INVX0 U1567 ( .INP(n2535), .ZN(n2500) );
  NAND2X0 U1568 ( .IN1(n998), .IN2(reg1[28]), .QN(n1205) );
  NAND2X0 U1569 ( .IN1(n997), .IN2(reg0[28]), .QN(n1204) );
  NAND2X0 U1570 ( .IN1(n999), .IN2(reg2[28]), .QN(n1203) );
  NAND2X0 U1571 ( .IN1(n1200), .IN2(reg3[28]), .QN(n2538) );
  OA21X1 U1572 ( .IN1(n1200), .IN2(reg3[28]), .IN3(n2538), .Q(n2502) );
  NAND2X0 U1573 ( .IN1(n2502), .IN2(n1201), .QN(n1202) );
  NAND4X0 U1574 ( .IN1(n1205), .IN2(n1204), .IN3(n1203), .IN4(n1202), .QN(
        n2689) );
  NAND2X0 U1575 ( .IN1(n2500), .IN2(n2689), .QN(n2508) );
  NAND2X0 U1576 ( .IN1(datai[29]), .IN2(n2520), .QN(n2536) );
  NOR2X0 U1577 ( .IN1(n1206), .IN2(n2538), .QN(n1208) );
  AO22X1 U1578 ( .IN1(n999), .IN2(reg2[29]), .IN3(n997), .IN4(reg0[29]), .Q(
        n1207) );
  NOR2X0 U1579 ( .IN1(n1208), .IN2(n1207), .QN(n1210) );
  NAND2X0 U1580 ( .IN1(n998), .IN2(reg1[29]), .QN(n1209) );
  NAND2X0 U1581 ( .IN1(n1210), .IN2(n1209), .QN(n2690) );
  NAND2X0 U1582 ( .IN1(n2536), .IN2(n2690), .QN(n2505) );
  AO222X1 U1583 ( .IN1(n998), .IN2(reg1[31]), .IN3(n997), .IN4(reg0[31]), 
        .IN5(n999), .IN6(reg2[31]), .Q(n2692) );
  NAND2X0 U1584 ( .IN1(datai[31]), .IN2(n2520), .QN(n2550) );
  NOR2X0 U1585 ( .IN1(n2692), .IN2(n2550), .QN(n1330) );
  INVX0 U1586 ( .INP(n1330), .ZN(n1255) );
  AO222X1 U1587 ( .IN1(n998), .IN2(reg1[30]), .IN3(n999), .IN4(reg2[30]), 
        .IN5(n997), .IN6(reg0[30]), .Q(n2691) );
  INVX0 U1588 ( .INP(n2691), .ZN(n2518) );
  NAND2X0 U1589 ( .IN1(datai[30]), .IN2(n2520), .QN(n2547) );
  INVX0 U1590 ( .INP(n2547), .ZN(n2544) );
  NOR2X0 U1591 ( .IN1(n2518), .IN2(n2544), .QN(n1318) );
  INVX0 U1592 ( .INP(n1318), .ZN(n1211) );
  NAND4X0 U1593 ( .IN1(n2508), .IN2(n2505), .IN3(n1255), .IN4(n1211), .QN(
        n1269) );
  NOR2X0 U1594 ( .IN1(n1365), .IN2(n2688), .QN(n2488) );
  INVX0 U1595 ( .INP(n2687), .ZN(n1960) );
  NAND2X0 U1596 ( .IN1(n2475), .IN2(n1960), .QN(n2462) );
  INVX0 U1597 ( .INP(n2462), .ZN(n1392) );
  NOR2X0 U1598 ( .IN1(n2488), .IN2(n1392), .QN(n1249) );
  INVX0 U1599 ( .INP(n2689), .ZN(n1977) );
  NAND2X0 U1600 ( .IN1(n2535), .IN2(n1977), .QN(n2489) );
  INVX0 U1601 ( .INP(n2489), .ZN(n2510) );
  NAND2X0 U1602 ( .IN1(n2692), .IN2(n2550), .QN(n1319) );
  OA21X1 U1603 ( .IN1(n2547), .IN2(n2691), .IN3(n1319), .Q(n1267) );
  OR2X1 U1604 ( .IN1(n2536), .IN2(n2690), .Q(n2504) );
  NAND2X0 U1605 ( .IN1(n1267), .IN2(n2504), .QN(n1323) );
  NOR2X0 U1606 ( .IN1(n2510), .IN2(n1323), .QN(n1212) );
  NOR2X0 U1607 ( .IN1(n1412), .IN2(n2686), .QN(n1391) );
  INVX0 U1608 ( .INP(n1391), .ZN(n1413) );
  INVX0 U1609 ( .INP(n2685), .ZN(n1947) );
  NAND2X0 U1610 ( .IN1(n2452), .IN2(n1947), .QN(n2439) );
  NAND4X0 U1611 ( .IN1(n1249), .IN2(n1212), .IN3(n1413), .IN4(n2439), .QN(
        n1314) );
  NOR4X0 U1612 ( .IN1(n1248), .IN2(n1213), .IN3(n1269), .IN4(n1314), .QN(n1214) );
  NAND4X0 U1613 ( .IN1(n1215), .IN2(n1300), .IN3(n1311), .IN4(n1214), .QN(
        n1262) );
  AND2X1 U1614 ( .IN1(n2692), .IN2(n2691), .Q(n1218) );
  NAND2X0 U1615 ( .IN1(n2505), .IN2(n1255), .QN(n1216) );
  AO21X1 U1616 ( .IN1(n2489), .IN2(n2504), .IN3(n1216), .Q(n1270) );
  OR3X1 U1617 ( .IN1(n1218), .IN2(n2547), .IN3(n1330), .Q(n1217) );
  AO22X1 U1618 ( .IN1(n1218), .IN2(n2547), .IN3(n1270), .IN4(n1217), .Q(n1259)
         );
  NAND2X0 U1619 ( .IN1(n1218), .IN2(n2547), .QN(n1257) );
  NAND2X0 U1620 ( .IN1(n1585), .IN2(n1603), .QN(n1224) );
  NAND2X0 U1621 ( .IN1(n1667), .IN2(n1683), .QN(n1220) );
  NAND2X0 U1622 ( .IN1(n1626), .IN2(n1644), .QN(n1219) );
  AO22X1 U1623 ( .IN1(n1221), .IN2(n1220), .IN3(n1627), .IN4(n1219), .Q(n1223)
         );
  AND3X1 U1624 ( .IN1(n1545), .IN2(n1563), .IN3(n1586), .Q(n1222) );
  OA221X1 U1625 ( .IN1(n1224), .IN2(n1604), .IN3(n1224), .IN4(n1223), .IN5(
        n1222), .Q(n1236) );
  INVX0 U1626 ( .INP(n1225), .ZN(n1232) );
  NAND2X0 U1627 ( .IN1(n1295), .IN2(n1293), .QN(n1229) );
  OR2X1 U1628 ( .IN1(n1369), .IN2(n1367), .Q(n1227) );
  INVX0 U1629 ( .INP(n1279), .ZN(n1366) );
  INVX0 U1630 ( .INP(n1820), .ZN(n1822) );
  OA21X1 U1631 ( .IN1(n1283), .IN2(n1822), .IN3(n1285), .Q(n1801) );
  OA21X1 U1632 ( .IN1(n1226), .IN2(n1801), .IN3(n1799), .Q(n1788) );
  OA21X1 U1633 ( .IN1(n1788), .IN2(n1281), .IN3(n1782), .Q(n1759) );
  OA221X1 U1634 ( .IN1(n1227), .IN2(n1366), .IN3(n1227), .IN4(n1759), .IN5(
        n1368), .Q(n1228) );
  OA221X1 U1635 ( .IN1(n1229), .IN2(n1228), .IN3(n1229), .IN4(n1370), .IN5(
        n1372), .Q(n1231) );
  NAND2X0 U1636 ( .IN1(n1544), .IN2(n1562), .QN(n1230) );
  AO22X1 U1637 ( .IN1(n1232), .IN2(n1231), .IN3(n1545), .IN4(n1230), .Q(n1235)
         );
  INVX0 U1638 ( .INP(n1233), .ZN(n1234) );
  OA21X1 U1639 ( .IN1(n1236), .IN2(n1235), .IN3(n1234), .Q(n1244) );
  NAND2X0 U1640 ( .IN1(n1441), .IN2(n2393), .QN(n1242) );
  NAND2X0 U1641 ( .IN1(n1503), .IN2(n1521), .QN(n1238) );
  NAND2X0 U1642 ( .IN1(n1455), .IN2(n1480), .QN(n1237) );
  AO22X1 U1643 ( .IN1(n1239), .IN2(n1238), .IN3(n1456), .IN4(n1237), .Q(n1241)
         );
  AND3X1 U1644 ( .IN1(n1428), .IN2(n2417), .IN3(n1442), .Q(n1240) );
  OA221X1 U1645 ( .IN1(n1242), .IN2(n2394), .IN3(n1242), .IN4(n1241), .IN5(
        n1240), .Q(n1243) );
  NOR2X0 U1646 ( .IN1(n1244), .IN2(n1243), .QN(n1247) );
  NAND2X0 U1647 ( .IN1(n1427), .IN2(n2416), .QN(n1245) );
  NAND2X0 U1648 ( .IN1(n1428), .IN2(n1245), .QN(n1246) );
  NAND2X0 U1649 ( .IN1(n1247), .IN2(n1246), .QN(n1254) );
  INVX0 U1650 ( .INP(n1248), .ZN(n1253) );
  NAND2X0 U1651 ( .IN1(n1413), .IN2(n2439), .QN(n1252) );
  AND3X1 U1652 ( .IN1(n2486), .IN2(n2463), .IN3(n1414), .Q(n1251) );
  INVX0 U1653 ( .INP(n1249), .ZN(n1250) );
  AO222X1 U1654 ( .IN1(n1254), .IN2(n1253), .IN3(n1252), .IN4(n1251), .IN5(
        n1250), .IN6(n2486), .Q(n1266) );
  AND3X1 U1655 ( .IN1(n2508), .IN2(n2505), .IN3(n1255), .Q(n1256) );
  NAND3X0 U1656 ( .IN1(n1257), .IN2(n1266), .IN3(n1256), .QN(n1258) );
  AND3X1 U1657 ( .IN1(n1259), .IN2(n1258), .IN3(n1319), .Q(n1261) );
  MUX21X1 U1658 ( .IN1(IR[21]), .IN2(n2712), .S(n1260), .Q(n2645) );
  MUX21X1 U1659 ( .IN1(IR[21]), .IN2(n2645), .S(n2699), .Q(n2525) );
  MUX21X1 U1660 ( .IN1(n1262), .IN2(n1261), .S(n2525), .Q(n1263) );
  XOR2X1 U1661 ( .IN1(n1265), .IN2(n1263), .Q(n1264) );
  OA22X1 U1662 ( .IN1(n2519), .IN2(n2704), .IN3(n1363), .IN4(n1264), .Q(n1335)
         );
  INVX0 U1663 ( .INP(n2525), .ZN(n1397) );
  NAND2X0 U1664 ( .IN1(n1397), .IN2(n2555), .QN(n1396) );
  NAND2X0 U1665 ( .IN1(n1397), .IN2(n1265), .QN(n1466) );
  INVX0 U1666 ( .INP(n1266), .ZN(n1268) );
  OA222X1 U1667 ( .IN1(n1270), .IN2(n1318), .IN3(n1269), .IN4(n1268), .IN5(
        n1330), .IN6(n1267), .Q(n1271) );
  MUX21X1 U1668 ( .IN1(n1396), .IN2(n1466), .S(n1271), .Q(n1331) );
  NAND2X0 U1669 ( .IN1(n1428), .IN2(n2417), .QN(n1313) );
  NAND2X0 U1670 ( .IN1(n1586), .IN2(n1604), .QN(n1278) );
  INVX0 U1671 ( .INP(n1272), .ZN(n1275) );
  NAND2X0 U1672 ( .IN1(n1668), .IN2(n1684), .QN(n1274) );
  NAND2X0 U1673 ( .IN1(n1627), .IN2(n1645), .QN(n1273) );
  AO22X1 U1674 ( .IN1(n1275), .IN2(n1274), .IN3(n1626), .IN4(n1273), .Q(n1277)
         );
  INVX0 U1675 ( .INP(n1562), .ZN(n1380) );
  NOR3X0 U1676 ( .IN1(n1381), .IN2(n1380), .IN3(n1379), .QN(n1276) );
  OA221X1 U1677 ( .IN1(n1278), .IN2(n1603), .IN3(n1278), .IN4(n1277), .IN5(
        n1276), .Q(n1310) );
  NAND2X0 U1678 ( .IN1(n1372), .IN2(n1370), .QN(n1297) );
  NOR2X0 U1679 ( .IN1(n1280), .IN2(n1279), .QN(n1292) );
  NOR2X0 U1680 ( .IN1(n1799), .IN2(n1281), .QN(n1290) );
  INVX0 U1681 ( .INP(n1281), .ZN(n1781) );
  NAND2X0 U1682 ( .IN1(n1798), .IN2(n1781), .QN(n1282) );
  NOR2X0 U1683 ( .IN1(n1283), .IN2(n1282), .QN(n1287) );
  NAND2X0 U1684 ( .IN1(n1285), .IN2(n1284), .QN(n1286) );
  NAND2X0 U1685 ( .IN1(n1287), .IN2(n1286), .QN(n1288) );
  NAND2X0 U1686 ( .IN1(n1288), .IN2(n1782), .QN(n1289) );
  NOR2X0 U1687 ( .IN1(n1290), .IN2(n1289), .QN(n1291) );
  AO221X1 U1688 ( .IN1(n1292), .IN2(n1291), .IN3(n1292), .IN4(n1367), .IN5(
        n1369), .Q(n1294) );
  INVX0 U1689 ( .INP(n1293), .ZN(n1371) );
  NOR2X0 U1690 ( .IN1(n1294), .IN2(n1371), .QN(n1296) );
  OA21X1 U1691 ( .IN1(n1297), .IN2(n1296), .IN3(n1295), .Q(n1299) );
  NAND2X0 U1692 ( .IN1(n1545), .IN2(n1563), .QN(n1298) );
  AO22X1 U1693 ( .IN1(n1300), .IN2(n1299), .IN3(n1544), .IN4(n1298), .Q(n1309)
         );
  NAND2X0 U1694 ( .IN1(n1442), .IN2(n2394), .QN(n1307) );
  INVX0 U1695 ( .INP(n1301), .ZN(n1304) );
  NAND2X0 U1696 ( .IN1(n1504), .IN2(n1522), .QN(n1303) );
  NAND2X0 U1697 ( .IN1(n1456), .IN2(n1481), .QN(n1302) );
  AO22X1 U1698 ( .IN1(n1304), .IN2(n1303), .IN3(n1455), .IN4(n1302), .Q(n1306)
         );
  INVX0 U1699 ( .INP(n2416), .ZN(n1388) );
  NOR2X0 U1700 ( .IN1(n1388), .IN2(n1387), .QN(n1305) );
  OA221X1 U1701 ( .IN1(n1307), .IN2(n2393), .IN3(n1307), .IN4(n1306), .IN5(
        n1305), .Q(n1308) );
  AO221X1 U1702 ( .IN1(n1311), .IN2(n1310), .IN3(n1311), .IN4(n1309), .IN5(
        n1308), .Q(n1312) );
  NOR2X0 U1703 ( .IN1(n1313), .IN2(n1312), .QN(n1317) );
  INVX0 U1704 ( .INP(n1314), .ZN(n1315) );
  NAND2X0 U1705 ( .IN1(n1315), .IN2(n1427), .QN(n1316) );
  NOR2X0 U1706 ( .IN1(n1317), .IN2(n1316), .QN(n1329) );
  AND2X1 U1707 ( .IN1(n1319), .IN2(n1318), .Q(n1328) );
  NAND2X0 U1708 ( .IN1(n2508), .IN2(n2505), .QN(n1326) );
  NOR3X0 U1709 ( .IN1(n2488), .IN2(n1392), .IN3(n1391), .QN(n1322) );
  NAND2X0 U1710 ( .IN1(n1414), .IN2(n2440), .QN(n1321) );
  INVX0 U1711 ( .INP(n2488), .ZN(n1393) );
  NAND2X0 U1712 ( .IN1(n2486), .IN2(n2463), .QN(n1320) );
  AO22X1 U1713 ( .IN1(n1322), .IN2(n1321), .IN3(n1393), .IN4(n1320), .Q(n1325)
         );
  INVX0 U1714 ( .INP(n1323), .ZN(n1324) );
  OA221X1 U1715 ( .IN1(n1326), .IN2(n2489), .IN3(n1326), .IN4(n1325), .IN5(
        n1324), .Q(n1327) );
  NOR4X0 U1716 ( .IN1(n1330), .IN2(n1329), .IN3(n1328), .IN4(n1327), .QN(n1332) );
  AO221X1 U1717 ( .IN1(n1331), .IN2(n1332), .IN3(n1331), .IN4(n2555), .IN5(
        n1361), .Q(n1334) );
  NAND2X0 U1718 ( .IN1(n1363), .IN2(n2555), .QN(n1832) );
  INVX0 U1719 ( .INP(n1832), .ZN(n1840) );
  NAND3X0 U1720 ( .IN1(n1840), .IN2(n1332), .IN3(n2525), .QN(n1333) );
  NAND3X0 U1721 ( .IN1(n1335), .IN2(n1334), .IN3(n1333), .QN(n1336) );
  NAND3X0 U1722 ( .IN1(n1992), .IN2(state), .IN3(n1336), .QN(n1340) );
  NAND2X0 U1723 ( .IN1(n2525), .IN2(n1831), .QN(n1993) );
  INVX0 U1724 ( .INP(n1993), .ZN(n2529) );
  NAND2X0 U1725 ( .IN1(n1840), .IN2(n2529), .QN(n1337) );
  NOR4X0 U1726 ( .IN1(n1988), .IN2(n1996), .IN3(n1989), .IN4(n1337), .QN(n1338) );
  AO221X1 U1727 ( .IN1(state), .IN2(n1338), .IN3(state), .IN4(n1992), .IN5(
        n2704), .Q(n1339) );
  NAND2X0 U1728 ( .IN1(n1340), .IN2(n1339), .QN(n829) );
  MUX21X1 U1729 ( .IN1(datai[0]), .IN2(IR[0]), .S(state), .Q(n893) );
  MUX21X1 U1730 ( .IN1(datai[1]), .IN2(n2373), .S(state), .Q(n892) );
  NOR2X0 U1731 ( .IN1(n2703), .IN2(n2727), .QN(n2658) );
  NOR2X0 U1732 ( .IN1(n2699), .IN2(n2703), .QN(n2656) );
  AO22X1 U1733 ( .IN1(IR[2]), .IN2(n2656), .IN3(datai[2]), .IN4(n2703), .Q(
        n1341) );
  AO21X1 U1734 ( .IN1(n2658), .IN2(n1342), .IN3(n1341), .Q(n891) );
  MUX21X1 U1735 ( .IN1(datai[3]), .IN2(n2358), .S(state), .Q(n890) );
  AO22X1 U1736 ( .IN1(IR[4]), .IN2(n2656), .IN3(datai[4]), .IN4(n2703), .Q(
        n1343) );
  AO21X1 U1737 ( .IN1(n2658), .IN2(n1344), .IN3(n1343), .Q(n889) );
  MUX21X1 U1738 ( .IN1(datai[5]), .IN2(n2350), .S(state), .Q(n888) );
  AO22X1 U1739 ( .IN1(IR[6]), .IN2(n2656), .IN3(datai[6]), .IN4(n2703), .Q(
        n1345) );
  AO21X1 U1740 ( .IN1(n2658), .IN2(n1346), .IN3(n1345), .Q(n887) );
  MUX21X1 U1741 ( .IN1(datai[7]), .IN2(n2334), .S(state), .Q(n886) );
  AO22X1 U1742 ( .IN1(IR[8]), .IN2(n2656), .IN3(datai[8]), .IN4(n2703), .Q(
        n1347) );
  AO21X1 U1743 ( .IN1(n2658), .IN2(n1348), .IN3(n1347), .Q(n885) );
  MUX21X1 U1744 ( .IN1(datai[9]), .IN2(n2318), .S(state), .Q(n884) );
  AO22X1 U1745 ( .IN1(IR[10]), .IN2(n2656), .IN3(datai[10]), .IN4(n2703), .Q(
        n1349) );
  AO21X1 U1746 ( .IN1(n2658), .IN2(n1350), .IN3(n1349), .Q(n883) );
  MUX21X1 U1747 ( .IN1(datai[11]), .IN2(n2302), .S(state), .Q(n882) );
  AO22X1 U1748 ( .IN1(IR[12]), .IN2(n2656), .IN3(datai[12]), .IN4(n2703), .Q(
        n1351) );
  AO21X1 U1749 ( .IN1(n2658), .IN2(n1352), .IN3(n1351), .Q(n881) );
  MUX21X1 U1750 ( .IN1(datai[13]), .IN2(n2286), .S(state), .Q(n880) );
  AO22X1 U1751 ( .IN1(IR[14]), .IN2(n2656), .IN3(datai[14]), .IN4(n2703), .Q(
        n1353) );
  AO21X1 U1752 ( .IN1(n2658), .IN2(n1354), .IN3(n1353), .Q(n879) );
  MUX21X1 U1753 ( .IN1(datai[15]), .IN2(n2270), .S(state), .Q(n878) );
  AO22X1 U1754 ( .IN1(IR[16]), .IN2(n2656), .IN3(datai[16]), .IN4(n2703), .Q(
        n1355) );
  AO21X1 U1755 ( .IN1(n2658), .IN2(n1356), .IN3(n1355), .Q(n877) );
  MUX21X1 U1756 ( .IN1(datai[17]), .IN2(n2254), .S(state), .Q(n876) );
  AO22X1 U1757 ( .IN1(n2656), .IN2(IR[18]), .IN3(datai[18]), .IN4(n2703), .Q(
        n1357) );
  AO21X1 U1758 ( .IN1(n1358), .IN2(n2658), .IN3(n1357), .Q(n875) );
  AO22X1 U1759 ( .IN1(datai[19]), .IN2(n2703), .IN3(IR[19]), .IN4(n2656), .Q(
        n1359) );
  AO21X1 U1760 ( .IN1(n2658), .IN2(n1360), .IN3(n1359), .Q(n874) );
  NOR2X0 U1761 ( .IN1(n1361), .IN2(n1831), .QN(n2548) );
  INVX0 U1762 ( .INP(n2548), .ZN(n1467) );
  NOR2X0 U1763 ( .IN1(n2525), .IN2(n1467), .QN(n2578) );
  NAND2X0 U1764 ( .IN1(n2579), .IN2(n1816), .QN(n1813) );
  NOR2X0 U1765 ( .IN1(n1859), .IN2(n1813), .QN(n1777) );
  NAND2X0 U1766 ( .IN1(n1777), .IN2(n1780), .QN(n1776) );
  NOR2X0 U1767 ( .IN1(n2228), .IN2(n1776), .QN(n1741) );
  NAND2X0 U1768 ( .IN1(n1741), .IN2(n1744), .QN(n1740) );
  NOR2X0 U1769 ( .IN1(n2202), .IN2(n1740), .QN(n1704) );
  NAND2X0 U1770 ( .IN1(n1704), .IN2(n1707), .QN(n1703) );
  NOR2X0 U1771 ( .IN1(n2180), .IN2(n1703), .QN(n1663) );
  NAND2X0 U1772 ( .IN1(n1663), .IN2(n1666), .QN(n1662) );
  NOR2X0 U1773 ( .IN1(n2158), .IN2(n1662), .QN(n1622) );
  NAND2X0 U1774 ( .IN1(n1622), .IN2(n1625), .QN(n1621) );
  NOR2X0 U1775 ( .IN1(n2136), .IN2(n1621), .QN(n1581) );
  NAND2X0 U1776 ( .IN1(n1581), .IN2(n1584), .QN(n1580) );
  NOR2X0 U1777 ( .IN1(n2114), .IN2(n1580), .QN(n1540) );
  NAND2X0 U1778 ( .IN1(n1540), .IN2(n1543), .QN(n1539) );
  NOR2X0 U1779 ( .IN1(n2092), .IN2(n1539), .QN(n1499) );
  NAND2X0 U1780 ( .IN1(n1499), .IN2(n1502), .QN(n1498) );
  NOR2X0 U1781 ( .IN1(n2070), .IN2(n1498), .QN(n1452) );
  NAND2X0 U1782 ( .IN1(n1452), .IN2(n1454), .QN(n2405) );
  NOR2X0 U1783 ( .IN1(n2406), .IN2(n2405), .QN(n1438) );
  NAND2X0 U1784 ( .IN1(n1438), .IN2(n1440), .QN(n2428) );
  NOR2X0 U1785 ( .IN1(n2429), .IN2(n2428), .QN(n1424) );
  NAND2X0 U1786 ( .IN1(n1424), .IN2(n1426), .QN(n2451) );
  NOR2X0 U1787 ( .IN1(n2452), .IN2(n2451), .QN(n1410) );
  NAND2X0 U1788 ( .IN1(n1410), .IN2(n1412), .QN(n2474) );
  NOR2X0 U1789 ( .IN1(n2475), .IN2(n2474), .QN(n1362) );
  NAND2X0 U1790 ( .IN1(n1362), .IN2(n1365), .QN(n2534) );
  OA21X1 U1791 ( .IN1(n1362), .IN2(n1365), .IN3(n2534), .Q(n2480) );
  NOR2X0 U1792 ( .IN1(n1831), .IN2(n1363), .QN(n2554) );
  NAND2X0 U1793 ( .IN1(n1397), .IN2(n2554), .QN(n2527) );
  NAND3X0 U1794 ( .IN1(n2661), .IN2(n2660), .IN3(n2692), .QN(n1872) );
  NOR2X0 U1795 ( .IN1(n1858), .IN2(n1872), .QN(n1814) );
  NAND2X0 U1796 ( .IN1(n1814), .IN2(n2663), .QN(n1796) );
  NOR2X0 U1797 ( .IN1(n1922), .IN2(n1796), .QN(n1778) );
  NAND2X0 U1798 ( .IN1(n1778), .IN2(n2665), .QN(n1760) );
  NOR2X0 U1799 ( .IN1(n1920), .IN2(n1760), .QN(n1742) );
  NAND2X0 U1800 ( .IN1(n1742), .IN2(n2667), .QN(n1724) );
  NOR2X0 U1801 ( .IN1(n1918), .IN2(n1724), .QN(n1705) );
  NAND2X0 U1802 ( .IN1(n1705), .IN2(n2669), .QN(n1687) );
  NOR2X0 U1803 ( .IN1(n1916), .IN2(n1687), .QN(n1664) );
  NAND2X0 U1804 ( .IN1(n1664), .IN2(n2671), .QN(n1642) );
  NOR2X0 U1805 ( .IN1(n1914), .IN2(n1642), .QN(n1623) );
  NAND2X0 U1806 ( .IN1(n1623), .IN2(n2673), .QN(n1601) );
  NOR2X0 U1807 ( .IN1(n1912), .IN2(n1601), .QN(n1582) );
  NAND2X0 U1808 ( .IN1(n1582), .IN2(n2675), .QN(n1560) );
  NOR2X0 U1809 ( .IN1(n1910), .IN2(n1560), .QN(n1541) );
  NAND2X0 U1810 ( .IN1(n1541), .IN2(n2677), .QN(n1519) );
  NOR2X0 U1811 ( .IN1(n1907), .IN2(n1519), .QN(n1500) );
  NAND2X0 U1812 ( .IN1(n1500), .IN2(n2679), .QN(n1478) );
  NOR2X0 U1813 ( .IN1(n1905), .IN2(n1478), .QN(n1903) );
  NAND2X0 U1814 ( .IN1(n1903), .IN2(n2681), .QN(n1902) );
  NOR2X0 U1815 ( .IN1(n1934), .IN2(n1902), .QN(n1932) );
  NAND2X0 U1816 ( .IN1(n1932), .IN2(n2684), .QN(n1931) );
  NOR2X0 U1817 ( .IN1(n1947), .IN2(n1931), .QN(n1945) );
  NAND2X0 U1818 ( .IN1(n1945), .IN2(n2686), .QN(n1944) );
  NOR2X0 U1819 ( .IN1(n1960), .IN2(n1944), .QN(n1958) );
  NAND2X0 U1820 ( .IN1(n1958), .IN2(n2688), .QN(n1957) );
  NOR2X0 U1821 ( .IN1(n1977), .IN2(n1957), .QN(n1970) );
  AO21X1 U1822 ( .IN1(n1977), .IN2(n1957), .IN3(n1970), .Q(n1364) );
  INVX0 U1823 ( .INP(n1996), .ZN(n2528) );
  MUX21X1 U1824 ( .IN1(n1364), .IN2(n1960), .S(n2528), .Q(n2007) );
  OA22X1 U1825 ( .IN1(n2527), .IN2(n1365), .IN3(n1993), .IN4(n2007), .Q(n1403)
         );
  INVX0 U1826 ( .INP(n2439), .ZN(n1390) );
  INVX0 U1827 ( .INP(n2393), .ZN(n1386) );
  INVX0 U1828 ( .INP(n1480), .ZN(n1384) );
  INVX0 U1829 ( .INP(n1603), .ZN(n1378) );
  INVX0 U1830 ( .INP(n1644), .ZN(n1376) );
  OA21X1 U1831 ( .IN1(n1367), .IN2(n1759), .IN3(n1366), .Q(n1746) );
  OA21X1 U1832 ( .IN1(n1369), .IN2(n1746), .IN3(n1368), .Q(n1723) );
  OA21X1 U1833 ( .IN1(n1371), .IN2(n1723), .IN3(n1370), .Q(n1709) );
  OA21X1 U1834 ( .IN1(n1373), .IN2(n1709), .IN3(n1372), .Q(n1686) );
  OA21X1 U1835 ( .IN1(n1374), .IN2(n1686), .IN3(n1684), .Q(n1670) );
  OA21X1 U1836 ( .IN1(n1375), .IN2(n1670), .IN3(n1668), .Q(n1647) );
  OA21X1 U1837 ( .IN1(n1376), .IN2(n1647), .IN3(n1645), .Q(n1629) );
  OA21X1 U1838 ( .IN1(n1377), .IN2(n1629), .IN3(n1627), .Q(n1606) );
  OA21X1 U1839 ( .IN1(n1378), .IN2(n1606), .IN3(n1604), .Q(n1588) );
  OA21X1 U1840 ( .IN1(n1379), .IN2(n1588), .IN3(n1586), .Q(n1565) );
  OA21X1 U1841 ( .IN1(n1380), .IN2(n1565), .IN3(n1563), .Q(n1547) );
  OA21X1 U1842 ( .IN1(n1381), .IN2(n1547), .IN3(n1545), .Q(n1524) );
  OA21X1 U1843 ( .IN1(n1382), .IN2(n1524), .IN3(n1522), .Q(n1506) );
  OA21X1 U1844 ( .IN1(n1383), .IN2(n1506), .IN3(n1504), .Q(n1483) );
  OA21X1 U1845 ( .IN1(n1384), .IN2(n1483), .IN3(n1481), .Q(n1458) );
  OA21X1 U1846 ( .IN1(n1385), .IN2(n1458), .IN3(n1456), .Q(n2396) );
  OA21X1 U1847 ( .IN1(n1386), .IN2(n2396), .IN3(n2394), .Q(n1444) );
  OA21X1 U1848 ( .IN1(n1387), .IN2(n1444), .IN3(n1442), .Q(n2419) );
  OA21X1 U1849 ( .IN1(n1388), .IN2(n2419), .IN3(n2417), .Q(n1430) );
  OA21X1 U1850 ( .IN1(n1389), .IN2(n1430), .IN3(n1428), .Q(n2442) );
  OA21X1 U1851 ( .IN1(n1390), .IN2(n2442), .IN3(n2440), .Q(n1416) );
  OA21X1 U1852 ( .IN1(n1391), .IN2(n1416), .IN3(n1414), .Q(n2465) );
  OA21X1 U1853 ( .IN1(n1392), .IN2(n2465), .IN3(n2463), .Q(n2487) );
  NAND2X0 U1854 ( .IN1(n2486), .IN2(n1393), .QN(n1398) );
  INVX0 U1855 ( .INP(n2487), .ZN(n1395) );
  INVX0 U1856 ( .INP(n1398), .ZN(n1399) );
  INVX0 U1857 ( .INP(n2554), .ZN(n1394) );
  OA22X1 U1858 ( .IN1(n1397), .IN2(n1394), .IN3(n2519), .IN4(n1466), .Q(n2514)
         );
  AO221X1 U1859 ( .IN1(n2487), .IN2(n1398), .IN3(n1395), .IN4(n1399), .IN5(
        n2514), .Q(n1402) );
  NAND2X0 U1860 ( .IN1(n1885), .IN2(n2660), .QN(n1817) );
  INVX0 U1861 ( .INP(n1817), .ZN(n1818) );
  AO222X1 U1862 ( .IN1(n1837), .IN2(n1818), .IN3(n1837), .IN4(n2661), .IN5(
        n1818), .IN6(n2661), .Q(n1803) );
  INVX0 U1863 ( .INP(n1803), .ZN(n1805) );
  OA222X1 U1864 ( .IN1(n1810), .IN2(n1858), .IN3(n1810), .IN4(n1805), .IN5(
        n1858), .IN6(n1805), .Q(n1784) );
  INVX0 U1865 ( .INP(n1784), .ZN(n1783) );
  AO222X1 U1866 ( .IN1(n1901), .IN2(n2663), .IN3(n1901), .IN4(n1783), .IN5(
        n2663), .IN6(n1783), .Q(n1763) );
  INVX0 U1867 ( .INP(n1763), .ZN(n1765) );
  OA222X1 U1868 ( .IN1(n1770), .IN2(n1922), .IN3(n1770), .IN4(n1765), .IN5(
        n1922), .IN6(n1765), .Q(n1750) );
  INVX0 U1869 ( .INP(n1750), .ZN(n1748) );
  AO222X1 U1870 ( .IN1(n2214), .IN2(n2665), .IN3(n2214), .IN4(n1748), .IN5(
        n2665), .IN6(n1748), .Q(n1727) );
  INVX0 U1871 ( .INP(n1727), .ZN(n1729) );
  OA222X1 U1872 ( .IN1(n1734), .IN2(n1920), .IN3(n1734), .IN4(n1729), .IN5(
        n1920), .IN6(n1729), .Q(n1713) );
  INVX0 U1873 ( .INP(n1713), .ZN(n1711) );
  AO222X1 U1874 ( .IN1(n2191), .IN2(n2667), .IN3(n2191), .IN4(n1711), .IN5(
        n2667), .IN6(n1711), .Q(n1690) );
  INVX0 U1875 ( .INP(n1690), .ZN(n1692) );
  OA222X1 U1876 ( .IN1(n1697), .IN2(n1918), .IN3(n1697), .IN4(n1692), .IN5(
        n1918), .IN6(n1692), .Q(n1674) );
  INVX0 U1877 ( .INP(n1674), .ZN(n1672) );
  AO222X1 U1878 ( .IN1(n2169), .IN2(n2669), .IN3(n2169), .IN4(n1672), .IN5(
        n2669), .IN6(n1672), .Q(n1649) );
  INVX0 U1879 ( .INP(n1649), .ZN(n1651) );
  OA222X1 U1880 ( .IN1(n1656), .IN2(n1916), .IN3(n1656), .IN4(n1651), .IN5(
        n1916), .IN6(n1651), .Q(n1633) );
  INVX0 U1881 ( .INP(n1633), .ZN(n1631) );
  AO222X1 U1882 ( .IN1(n2147), .IN2(n2671), .IN3(n2147), .IN4(n1631), .IN5(
        n2671), .IN6(n1631), .Q(n1608) );
  INVX0 U1883 ( .INP(n1608), .ZN(n1610) );
  OA222X1 U1884 ( .IN1(n1615), .IN2(n1914), .IN3(n1615), .IN4(n1610), .IN5(
        n1914), .IN6(n1610), .Q(n1592) );
  INVX0 U1885 ( .INP(n1592), .ZN(n1590) );
  AO222X1 U1886 ( .IN1(n2125), .IN2(n2673), .IN3(n2125), .IN4(n1590), .IN5(
        n2673), .IN6(n1590), .Q(n1567) );
  INVX0 U1887 ( .INP(n1567), .ZN(n1569) );
  OA222X1 U1888 ( .IN1(n1574), .IN2(n1912), .IN3(n1574), .IN4(n1569), .IN5(
        n1912), .IN6(n1569), .Q(n1551) );
  INVX0 U1889 ( .INP(n1551), .ZN(n1549) );
  AO222X1 U1890 ( .IN1(n2103), .IN2(n2675), .IN3(n2103), .IN4(n1549), .IN5(
        n2675), .IN6(n1549), .Q(n1526) );
  INVX0 U1891 ( .INP(n1526), .ZN(n1528) );
  OA222X1 U1892 ( .IN1(n1533), .IN2(n1910), .IN3(n1533), .IN4(n1528), .IN5(
        n1910), .IN6(n1528), .Q(n1510) );
  INVX0 U1893 ( .INP(n1510), .ZN(n1508) );
  AO222X1 U1894 ( .IN1(n2081), .IN2(n2677), .IN3(n2081), .IN4(n1508), .IN5(
        n2677), .IN6(n1508), .Q(n1485) );
  INVX0 U1895 ( .INP(n1485), .ZN(n1487) );
  OA222X1 U1896 ( .IN1(n1492), .IN2(n1907), .IN3(n1492), .IN4(n1487), .IN5(
        n1907), .IN6(n1487), .Q(n1462) );
  INVX0 U1897 ( .INP(n1462), .ZN(n1460) );
  AO222X1 U1898 ( .IN1(n2059), .IN2(n2679), .IN3(n2059), .IN4(n1460), .IN5(
        n2679), .IN6(n1460), .Q(n2398) );
  INVX0 U1899 ( .INP(n2398), .ZN(n2400) );
  OA222X1 U1900 ( .IN1(n2407), .IN2(n1905), .IN3(n2407), .IN4(n2400), .IN5(
        n1905), .IN6(n2400), .Q(n1448) );
  INVX0 U1901 ( .INP(n1448), .ZN(n1446) );
  AO222X1 U1902 ( .IN1(n2048), .IN2(n2681), .IN3(n2048), .IN4(n1446), .IN5(
        n2681), .IN6(n1446), .Q(n2421) );
  INVX0 U1903 ( .INP(n2421), .ZN(n2423) );
  OA222X1 U1904 ( .IN1(n2430), .IN2(n1934), .IN3(n2430), .IN4(n2423), .IN5(
        n1934), .IN6(n2423), .Q(n1434) );
  INVX0 U1905 ( .INP(n1434), .ZN(n1432) );
  AO222X1 U1906 ( .IN1(n2036), .IN2(n2684), .IN3(n2036), .IN4(n1432), .IN5(
        n2684), .IN6(n1432), .Q(n2444) );
  INVX0 U1907 ( .INP(n2444), .ZN(n2446) );
  OA222X1 U1908 ( .IN1(n2453), .IN2(n1947), .IN3(n2453), .IN4(n2446), .IN5(
        n1947), .IN6(n2446), .Q(n1420) );
  INVX0 U1909 ( .INP(n1420), .ZN(n1418) );
  AO222X1 U1910 ( .IN1(n2024), .IN2(n2686), .IN3(n2024), .IN4(n1418), .IN5(
        n2686), .IN6(n1418), .Q(n2467) );
  INVX0 U1911 ( .INP(n2467), .ZN(n2469) );
  OA222X1 U1912 ( .IN1(n2476), .IN2(n1960), .IN3(n2476), .IN4(n2469), .IN5(
        n1960), .IN6(n2469), .Q(n1400) );
  INVX0 U1913 ( .INP(n1400), .ZN(n2491) );
  OA22X1 U1914 ( .IN1(n1397), .IN2(n1467), .IN3(n2519), .IN4(n1396), .Q(n2516)
         );
  AO221X1 U1915 ( .IN1(n1400), .IN2(n1399), .IN3(n2491), .IN4(n1398), .IN5(
        n2516), .Q(n1401) );
  NAND3X0 U1916 ( .IN1(n1403), .IN2(n1402), .IN3(n1401), .QN(n2483) );
  AO21X1 U1917 ( .IN1(n2578), .IN2(n2480), .IN3(n2483), .Q(n2634) );
  NOR2X0 U1918 ( .IN1(n1405), .IN2(n1404), .QN(n2575) );
  OR2X1 U1919 ( .IN1(n1405), .IN2(n1468), .Q(n2697) );
  MUX21X1 U1920 ( .IN1(n2704), .IN2(B), .S(n1404), .Q(n1406) );
  OA21X1 U1921 ( .IN1(n1468), .IN2(n1406), .IN3(n1405), .Q(n2574) );
  NAND2X0 U1922 ( .IN1(n2574), .IN2(d[0]), .QN(n1828) );
  OA22X1 U1923 ( .IN1(n2575), .IN2(n2697), .IN3(d[1]), .IN4(n1828), .Q(n1409)
         );
  NOR2X0 U1924 ( .IN1(n2525), .IN2(n1831), .QN(n1473) );
  NOR2X0 U1925 ( .IN1(n2529), .IN2(n1473), .QN(n1909) );
  NOR2X0 U1926 ( .IN1(n1840), .IN2(n1909), .QN(n1407) );
  NAND2X0 U1927 ( .IN1(n1407), .IN2(n2527), .QN(n1408) );
  NOR2X0 U1928 ( .IN1(n1988), .IN2(n1992), .QN(n2694) );
  NAND3X0 U1929 ( .IN1(n1408), .IN2(state), .IN3(n2694), .QN(n2576) );
  OR2X1 U1930 ( .IN1(n1409), .IN2(n2576), .Q(n2573) );
  INVX0 U1931 ( .INP(n2573), .ZN(n2565) );
  MUX21X1 U1932 ( .IN1(reg1[27]), .IN2(n2634), .S(n2565), .Q(n930) );
  OA21X1 U1933 ( .IN1(n1410), .IN2(n1412), .IN3(n2474), .Q(n2457) );
  AO21X1 U1934 ( .IN1(n1960), .IN2(n1944), .IN3(n1958), .Q(n1411) );
  MUX21X1 U1935 ( .IN1(n1411), .IN2(n1947), .S(n2528), .Q(n2018) );
  OA22X1 U1936 ( .IN1(n2527), .IN2(n1412), .IN3(n1993), .IN4(n2018), .Q(n1423)
         );
  NAND2X0 U1937 ( .IN1(n1414), .IN2(n1413), .QN(n1417) );
  INVX0 U1938 ( .INP(n1416), .ZN(n1415) );
  INVX0 U1939 ( .INP(n1417), .ZN(n1419) );
  AO221X1 U1940 ( .IN1(n1416), .IN2(n1417), .IN3(n1415), .IN4(n1419), .IN5(
        n2514), .Q(n1422) );
  AO221X1 U1941 ( .IN1(n1420), .IN2(n1419), .IN3(n1418), .IN4(n1417), .IN5(
        n2516), .Q(n1421) );
  NAND3X0 U1942 ( .IN1(n1423), .IN2(n1422), .IN3(n1421), .QN(n2460) );
  AO21X1 U1943 ( .IN1(n2578), .IN2(n2457), .IN3(n2460), .Q(n2630) );
  MUX21X1 U1944 ( .IN1(reg1[25]), .IN2(n2630), .S(n2565), .Q(n932) );
  OA21X1 U1945 ( .IN1(n1424), .IN2(n1426), .IN3(n2451), .Q(n2434) );
  AO21X1 U1946 ( .IN1(n1947), .IN2(n1931), .IN3(n1945), .Q(n1425) );
  MUX21X1 U1947 ( .IN1(n1425), .IN2(n1934), .S(n2528), .Q(n2030) );
  OA22X1 U1948 ( .IN1(n2527), .IN2(n1426), .IN3(n1993), .IN4(n2030), .Q(n1437)
         );
  NAND2X0 U1949 ( .IN1(n1428), .IN2(n1427), .QN(n1431) );
  INVX0 U1950 ( .INP(n1430), .ZN(n1429) );
  INVX0 U1951 ( .INP(n1431), .ZN(n1433) );
  AO221X1 U1952 ( .IN1(n1430), .IN2(n1431), .IN3(n1429), .IN4(n1433), .IN5(
        n2514), .Q(n1436) );
  AO221X1 U1953 ( .IN1(n1434), .IN2(n1433), .IN3(n1432), .IN4(n1431), .IN5(
        n2516), .Q(n1435) );
  NAND3X0 U1954 ( .IN1(n1437), .IN2(n1436), .IN3(n1435), .QN(n2437) );
  AO21X1 U1955 ( .IN1(n2578), .IN2(n2434), .IN3(n2437), .Q(n2626) );
  MUX21X1 U1956 ( .IN1(reg1[23]), .IN2(n2626), .S(n2565), .Q(n934) );
  OA21X1 U1957 ( .IN1(n1438), .IN2(n1440), .IN3(n2428), .Q(n2411) );
  AO21X1 U1958 ( .IN1(n1934), .IN2(n1902), .IN3(n1932), .Q(n1439) );
  MUX21X1 U1959 ( .IN1(n1439), .IN2(n1905), .S(n2528), .Q(n2042) );
  OA22X1 U1960 ( .IN1(n2527), .IN2(n1440), .IN3(n1993), .IN4(n2042), .Q(n1451)
         );
  NAND2X0 U1961 ( .IN1(n1442), .IN2(n1441), .QN(n1445) );
  INVX0 U1962 ( .INP(n1444), .ZN(n1443) );
  INVX0 U1963 ( .INP(n1445), .ZN(n1447) );
  AO221X1 U1964 ( .IN1(n1444), .IN2(n1445), .IN3(n1443), .IN4(n1447), .IN5(
        n2514), .Q(n1450) );
  AO221X1 U1965 ( .IN1(n1448), .IN2(n1447), .IN3(n1446), .IN4(n1445), .IN5(
        n2516), .Q(n1449) );
  NAND3X0 U1966 ( .IN1(n1451), .IN2(n1450), .IN3(n1449), .QN(n2414) );
  AO21X1 U1967 ( .IN1(n2578), .IN2(n2411), .IN3(n2414), .Q(n2622) );
  MUX21X1 U1968 ( .IN1(reg1[21]), .IN2(n2622), .S(n2565), .Q(n936) );
  OA21X1 U1969 ( .IN1(n1452), .IN2(n1454), .IN3(n2405), .Q(n1474) );
  AO21X1 U1970 ( .IN1(n1905), .IN2(n1478), .IN3(n1903), .Q(n1453) );
  MUX21X1 U1971 ( .IN1(n1453), .IN2(n1907), .S(n2528), .Q(n2054) );
  OA22X1 U1972 ( .IN1(n2527), .IN2(n1454), .IN3(n1993), .IN4(n2054), .Q(n1465)
         );
  NAND2X0 U1973 ( .IN1(n1456), .IN2(n1455), .QN(n1459) );
  INVX0 U1974 ( .INP(n1458), .ZN(n1457) );
  INVX0 U1975 ( .INP(n1459), .ZN(n1461) );
  AO221X1 U1976 ( .IN1(n1458), .IN2(n1459), .IN3(n1457), .IN4(n1461), .IN5(
        n2514), .Q(n1464) );
  AO221X1 U1977 ( .IN1(n1462), .IN2(n1461), .IN3(n1460), .IN4(n1459), .IN5(
        n2516), .Q(n1463) );
  NAND3X0 U1978 ( .IN1(n1465), .IN2(n1464), .IN3(n1463), .QN(n1477) );
  AO21X1 U1979 ( .IN1(n2578), .IN2(n1474), .IN3(n1477), .Q(n2618) );
  MUX21X1 U1980 ( .IN1(reg1[19]), .IN2(n2618), .S(n2565), .Q(n938) );
  NOR2X0 U1981 ( .IN1(n1467), .IN2(n1466), .QN(n1826) );
  INVX0 U1982 ( .INP(n2574), .ZN(n2693) );
  NOR2X0 U1983 ( .IN1(n2693), .IN2(n2709), .QN(n1469) );
  AO22X1 U1984 ( .IN1(n1469), .IN2(n2700), .IN3(n2575), .IN4(n1468), .Q(n1470)
         );
  INVX0 U1985 ( .INP(n2694), .ZN(n2391) );
  AO21X1 U1986 ( .IN1(n1832), .IN2(n2529), .IN3(n2391), .Q(n1848) );
  NOR2X0 U1987 ( .IN1(n2703), .IN2(n1848), .QN(n1472) );
  OA21X1 U1988 ( .IN1(n1826), .IN2(n1470), .IN3(n1472), .Q(n2556) );
  INVX0 U1989 ( .INP(n2556), .ZN(n2558) );
  INVX0 U1990 ( .INP(n1471), .ZN(n2049) );
  AND2X1 U1991 ( .IN1(n1826), .IN2(n1472), .Q(n2539) );
  NAND2X0 U1992 ( .IN1(n1473), .IN2(n1840), .QN(n1834) );
  NOR2X0 U1993 ( .IN1(n2558), .IN2(n1834), .QN(n2541) );
  AO22X1 U1994 ( .IN1(n2049), .IN2(n2539), .IN3(n2541), .IN4(n1474), .Q(n1475)
         );
  AO21X1 U1995 ( .IN1(reg2[19]), .IN2(n2558), .IN3(n1475), .Q(n1476) );
  AO21X1 U1996 ( .IN1(n2556), .IN2(n1477), .IN3(n1476), .Q(n970) );
  OA21X1 U1997 ( .IN1(n1500), .IN2(n2679), .IN3(n1478), .Q(n1479) );
  MUX21X1 U1998 ( .IN1(n1479), .IN2(n2677), .S(n2528), .Q(n2060) );
  NAND2X0 U1999 ( .IN1(n2529), .IN2(n2060), .QN(n1491) );
  INVX0 U2000 ( .INP(n2527), .ZN(n2485) );
  NAND2X0 U2001 ( .IN1(n2485), .IN2(n2070), .QN(n1490) );
  NAND2X0 U2002 ( .IN1(n1481), .IN2(n1480), .QN(n1484) );
  INVX0 U2003 ( .INP(n1483), .ZN(n1482) );
  INVX0 U2004 ( .INP(n1484), .ZN(n1486) );
  AO221X1 U2005 ( .IN1(n1483), .IN2(n1484), .IN3(n1482), .IN4(n1486), .IN5(
        n2514), .Q(n1489) );
  AO221X1 U2006 ( .IN1(n1487), .IN2(n1486), .IN3(n1485), .IN4(n1484), .IN5(
        n2516), .Q(n1488) );
  NAND4X0 U2007 ( .IN1(n1491), .IN2(n1490), .IN3(n1489), .IN4(n1488), .QN(
        n2617) );
  NAND2X0 U2008 ( .IN1(n2565), .IN2(n2578), .QN(n2563) );
  MUX21X1 U2009 ( .IN1(n1492), .IN2(n2070), .S(n1498), .Q(n2615) );
  NOR2X0 U2010 ( .IN1(n2563), .IN2(n2615), .QN(n1493) );
  AO21X1 U2011 ( .IN1(reg1[18]), .IN2(n2573), .IN3(n1493), .Q(n1494) );
  AO21X1 U2012 ( .IN1(n2565), .IN2(n2617), .IN3(n1494), .Q(n939) );
  INVX0 U2013 ( .INP(n2615), .ZN(n1495) );
  AO22X1 U2014 ( .IN1(n2065), .IN2(n2539), .IN3(n2541), .IN4(n1495), .Q(n1496)
         );
  AO21X1 U2015 ( .IN1(reg2[18]), .IN2(n2558), .IN3(n1496), .Q(n1497) );
  AO21X1 U2016 ( .IN1(n2556), .IN2(n2617), .IN3(n1497), .Q(n971) );
  OA21X1 U2017 ( .IN1(n1499), .IN2(n1502), .IN3(n1498), .Q(n1515) );
  AO21X1 U2018 ( .IN1(n1907), .IN2(n1519), .IN3(n1500), .Q(n1501) );
  MUX21X1 U2019 ( .IN1(n1501), .IN2(n1910), .S(n2528), .Q(n2076) );
  OA22X1 U2020 ( .IN1(n2527), .IN2(n1502), .IN3(n1993), .IN4(n2076), .Q(n1513)
         );
  NAND2X0 U2021 ( .IN1(n1504), .IN2(n1503), .QN(n1507) );
  INVX0 U2022 ( .INP(n1506), .ZN(n1505) );
  INVX0 U2023 ( .INP(n1507), .ZN(n1509) );
  AO221X1 U2024 ( .IN1(n1506), .IN2(n1507), .IN3(n1505), .IN4(n1509), .IN5(
        n2514), .Q(n1512) );
  AO221X1 U2025 ( .IN1(n1510), .IN2(n1509), .IN3(n1508), .IN4(n1507), .IN5(
        n2516), .Q(n1511) );
  NAND3X0 U2026 ( .IN1(n1513), .IN2(n1512), .IN3(n1511), .QN(n1518) );
  AO21X1 U2027 ( .IN1(n2578), .IN2(n1515), .IN3(n1518), .Q(n2614) );
  MUX21X1 U2028 ( .IN1(reg1[17]), .IN2(n2614), .S(n2565), .Q(n940) );
  INVX0 U2029 ( .INP(n1514), .ZN(n2071) );
  AO22X1 U2030 ( .IN1(n2071), .IN2(n2539), .IN3(n2541), .IN4(n1515), .Q(n1516)
         );
  AO21X1 U2031 ( .IN1(reg2[17]), .IN2(n2558), .IN3(n1516), .Q(n1517) );
  AO21X1 U2032 ( .IN1(n2556), .IN2(n1518), .IN3(n1517), .Q(n972) );
  OA21X1 U2033 ( .IN1(n1541), .IN2(n2677), .IN3(n1519), .Q(n1520) );
  MUX21X1 U2034 ( .IN1(n1520), .IN2(n2675), .S(n2528), .Q(n2082) );
  NAND2X0 U2035 ( .IN1(n2529), .IN2(n2082), .QN(n1532) );
  NAND2X0 U2036 ( .IN1(n2485), .IN2(n2092), .QN(n1531) );
  NAND2X0 U2037 ( .IN1(n1522), .IN2(n1521), .QN(n1525) );
  INVX0 U2038 ( .INP(n1524), .ZN(n1523) );
  INVX0 U2039 ( .INP(n1525), .ZN(n1527) );
  AO221X1 U2040 ( .IN1(n1524), .IN2(n1525), .IN3(n1523), .IN4(n1527), .IN5(
        n2514), .Q(n1530) );
  AO221X1 U2041 ( .IN1(n1528), .IN2(n1527), .IN3(n1526), .IN4(n1525), .IN5(
        n2516), .Q(n1529) );
  NAND4X0 U2042 ( .IN1(n1532), .IN2(n1531), .IN3(n1530), .IN4(n1529), .QN(
        n2613) );
  MUX21X1 U2043 ( .IN1(n1533), .IN2(n2092), .S(n1539), .Q(n2611) );
  NOR2X0 U2044 ( .IN1(n2563), .IN2(n2611), .QN(n1534) );
  AO21X1 U2045 ( .IN1(reg1[16]), .IN2(n2573), .IN3(n1534), .Q(n1535) );
  AO21X1 U2046 ( .IN1(n2565), .IN2(n2613), .IN3(n1535), .Q(n941) );
  INVX0 U2047 ( .INP(n2611), .ZN(n1536) );
  AO22X1 U2048 ( .IN1(n2087), .IN2(n2539), .IN3(n2541), .IN4(n1536), .Q(n1537)
         );
  AO21X1 U2049 ( .IN1(reg2[16]), .IN2(n2558), .IN3(n1537), .Q(n1538) );
  AO21X1 U2050 ( .IN1(n2556), .IN2(n2613), .IN3(n1538), .Q(n973) );
  OA21X1 U2051 ( .IN1(n1540), .IN2(n1543), .IN3(n1539), .Q(n1556) );
  AO21X1 U2052 ( .IN1(n1910), .IN2(n1560), .IN3(n1541), .Q(n1542) );
  MUX21X1 U2053 ( .IN1(n1542), .IN2(n1912), .S(n2528), .Q(n2098) );
  OA22X1 U2054 ( .IN1(n2527), .IN2(n1543), .IN3(n1993), .IN4(n2098), .Q(n1554)
         );
  NAND2X0 U2055 ( .IN1(n1545), .IN2(n1544), .QN(n1548) );
  INVX0 U2056 ( .INP(n1547), .ZN(n1546) );
  INVX0 U2057 ( .INP(n1548), .ZN(n1550) );
  AO221X1 U2058 ( .IN1(n1547), .IN2(n1548), .IN3(n1546), .IN4(n1550), .IN5(
        n2514), .Q(n1553) );
  AO221X1 U2059 ( .IN1(n1551), .IN2(n1550), .IN3(n1549), .IN4(n1548), .IN5(
        n2516), .Q(n1552) );
  NAND3X0 U2060 ( .IN1(n1554), .IN2(n1553), .IN3(n1552), .QN(n1559) );
  AO21X1 U2061 ( .IN1(n2578), .IN2(n1556), .IN3(n1559), .Q(n2610) );
  MUX21X1 U2062 ( .IN1(reg1[15]), .IN2(n2610), .S(n2565), .Q(n942) );
  INVX0 U2063 ( .INP(n1555), .ZN(n2093) );
  AO22X1 U2064 ( .IN1(n2093), .IN2(n2539), .IN3(n2541), .IN4(n1556), .Q(n1557)
         );
  AO21X1 U2065 ( .IN1(reg2[15]), .IN2(n2558), .IN3(n1557), .Q(n1558) );
  AO21X1 U2066 ( .IN1(n2556), .IN2(n1559), .IN3(n1558), .Q(n974) );
  OA21X1 U2067 ( .IN1(n1582), .IN2(n2675), .IN3(n1560), .Q(n1561) );
  MUX21X1 U2068 ( .IN1(n1561), .IN2(n2673), .S(n2528), .Q(n2104) );
  NAND2X0 U2069 ( .IN1(n2529), .IN2(n2104), .QN(n1573) );
  NAND2X0 U2070 ( .IN1(n2485), .IN2(n2114), .QN(n1572) );
  NAND2X0 U2071 ( .IN1(n1563), .IN2(n1562), .QN(n1566) );
  INVX0 U2072 ( .INP(n1565), .ZN(n1564) );
  INVX0 U2073 ( .INP(n1566), .ZN(n1568) );
  AO221X1 U2074 ( .IN1(n1565), .IN2(n1566), .IN3(n1564), .IN4(n1568), .IN5(
        n2514), .Q(n1571) );
  AO221X1 U2075 ( .IN1(n1569), .IN2(n1568), .IN3(n1567), .IN4(n1566), .IN5(
        n2516), .Q(n1570) );
  NAND4X0 U2076 ( .IN1(n1573), .IN2(n1572), .IN3(n1571), .IN4(n1570), .QN(
        n2609) );
  MUX21X1 U2077 ( .IN1(n1574), .IN2(n2114), .S(n1580), .Q(n2607) );
  NOR2X0 U2078 ( .IN1(n2563), .IN2(n2607), .QN(n1575) );
  AO21X1 U2079 ( .IN1(reg1[14]), .IN2(n2573), .IN3(n1575), .Q(n1576) );
  AO21X1 U2080 ( .IN1(n2565), .IN2(n2609), .IN3(n1576), .Q(n943) );
  INVX0 U2081 ( .INP(n2607), .ZN(n1577) );
  AO22X1 U2082 ( .IN1(n2109), .IN2(n2539), .IN3(n2541), .IN4(n1577), .Q(n1578)
         );
  AO21X1 U2083 ( .IN1(reg2[14]), .IN2(n2558), .IN3(n1578), .Q(n1579) );
  AO21X1 U2084 ( .IN1(n2556), .IN2(n2609), .IN3(n1579), .Q(n975) );
  OA21X1 U2085 ( .IN1(n1581), .IN2(n1584), .IN3(n1580), .Q(n1597) );
  AO21X1 U2086 ( .IN1(n1912), .IN2(n1601), .IN3(n1582), .Q(n1583) );
  MUX21X1 U2087 ( .IN1(n1583), .IN2(n1914), .S(n2528), .Q(n2120) );
  OA22X1 U2088 ( .IN1(n2527), .IN2(n1584), .IN3(n1993), .IN4(n2120), .Q(n1595)
         );
  NAND2X0 U2089 ( .IN1(n1586), .IN2(n1585), .QN(n1589) );
  INVX0 U2090 ( .INP(n1588), .ZN(n1587) );
  INVX0 U2091 ( .INP(n1589), .ZN(n1591) );
  AO221X1 U2092 ( .IN1(n1588), .IN2(n1589), .IN3(n1587), .IN4(n1591), .IN5(
        n2514), .Q(n1594) );
  AO221X1 U2093 ( .IN1(n1592), .IN2(n1591), .IN3(n1590), .IN4(n1589), .IN5(
        n2516), .Q(n1593) );
  NAND3X0 U2094 ( .IN1(n1595), .IN2(n1594), .IN3(n1593), .QN(n1600) );
  AO21X1 U2095 ( .IN1(n2578), .IN2(n1597), .IN3(n1600), .Q(n2606) );
  MUX21X1 U2096 ( .IN1(reg1[13]), .IN2(n2606), .S(n2565), .Q(n944) );
  INVX0 U2097 ( .INP(n1596), .ZN(n2115) );
  AO22X1 U2098 ( .IN1(n2115), .IN2(n2539), .IN3(n2541), .IN4(n1597), .Q(n1598)
         );
  AO21X1 U2099 ( .IN1(reg2[13]), .IN2(n2558), .IN3(n1598), .Q(n1599) );
  AO21X1 U2100 ( .IN1(n2556), .IN2(n1600), .IN3(n1599), .Q(n976) );
  OA21X1 U2101 ( .IN1(n1623), .IN2(n2673), .IN3(n1601), .Q(n1602) );
  MUX21X1 U2102 ( .IN1(n1602), .IN2(n2671), .S(n2528), .Q(n2126) );
  NAND2X0 U2103 ( .IN1(n2529), .IN2(n2126), .QN(n1614) );
  NAND2X0 U2104 ( .IN1(n2485), .IN2(n2136), .QN(n1613) );
  NAND2X0 U2105 ( .IN1(n1604), .IN2(n1603), .QN(n1607) );
  INVX0 U2106 ( .INP(n1606), .ZN(n1605) );
  INVX0 U2107 ( .INP(n1607), .ZN(n1609) );
  AO221X1 U2108 ( .IN1(n1606), .IN2(n1607), .IN3(n1605), .IN4(n1609), .IN5(
        n2514), .Q(n1612) );
  AO221X1 U2109 ( .IN1(n1610), .IN2(n1609), .IN3(n1608), .IN4(n1607), .IN5(
        n2516), .Q(n1611) );
  NAND4X0 U2110 ( .IN1(n1614), .IN2(n1613), .IN3(n1612), .IN4(n1611), .QN(
        n2605) );
  MUX21X1 U2111 ( .IN1(n1615), .IN2(n2136), .S(n1621), .Q(n2603) );
  NOR2X0 U2112 ( .IN1(n2563), .IN2(n2603), .QN(n1616) );
  AO21X1 U2113 ( .IN1(reg1[12]), .IN2(n2573), .IN3(n1616), .Q(n1617) );
  AO21X1 U2114 ( .IN1(n2565), .IN2(n2605), .IN3(n1617), .Q(n945) );
  INVX0 U2115 ( .INP(n2603), .ZN(n1618) );
  AO22X1 U2116 ( .IN1(n2131), .IN2(n2539), .IN3(n2541), .IN4(n1618), .Q(n1619)
         );
  AO21X1 U2117 ( .IN1(reg2[12]), .IN2(n2558), .IN3(n1619), .Q(n1620) );
  AO21X1 U2118 ( .IN1(n2556), .IN2(n2605), .IN3(n1620), .Q(n977) );
  OA21X1 U2119 ( .IN1(n1622), .IN2(n1625), .IN3(n1621), .Q(n1638) );
  AO21X1 U2120 ( .IN1(n1914), .IN2(n1642), .IN3(n1623), .Q(n1624) );
  MUX21X1 U2121 ( .IN1(n1624), .IN2(n1916), .S(n2528), .Q(n2142) );
  OA22X1 U2122 ( .IN1(n2527), .IN2(n1625), .IN3(n1993), .IN4(n2142), .Q(n1636)
         );
  NAND2X0 U2123 ( .IN1(n1627), .IN2(n1626), .QN(n1630) );
  INVX0 U2124 ( .INP(n1629), .ZN(n1628) );
  INVX0 U2125 ( .INP(n1630), .ZN(n1632) );
  AO221X1 U2126 ( .IN1(n1629), .IN2(n1630), .IN3(n1628), .IN4(n1632), .IN5(
        n2514), .Q(n1635) );
  AO221X1 U2127 ( .IN1(n1633), .IN2(n1632), .IN3(n1631), .IN4(n1630), .IN5(
        n2516), .Q(n1634) );
  NAND3X0 U2128 ( .IN1(n1636), .IN2(n1635), .IN3(n1634), .QN(n1641) );
  AO21X1 U2129 ( .IN1(n2578), .IN2(n1638), .IN3(n1641), .Q(n2602) );
  MUX21X1 U2130 ( .IN1(reg1[11]), .IN2(n2602), .S(n2565), .Q(n946) );
  INVX0 U2131 ( .INP(n1637), .ZN(n2137) );
  AO22X1 U2132 ( .IN1(n2137), .IN2(n2539), .IN3(n2541), .IN4(n1638), .Q(n1639)
         );
  AO21X1 U2133 ( .IN1(reg2[11]), .IN2(n2558), .IN3(n1639), .Q(n1640) );
  AO21X1 U2134 ( .IN1(n2556), .IN2(n1641), .IN3(n1640), .Q(n978) );
  OA21X1 U2135 ( .IN1(n1664), .IN2(n2671), .IN3(n1642), .Q(n1643) );
  MUX21X1 U2136 ( .IN1(n1643), .IN2(n2669), .S(n2528), .Q(n2148) );
  NAND2X0 U2137 ( .IN1(n2529), .IN2(n2148), .QN(n1655) );
  NAND2X0 U2138 ( .IN1(n2485), .IN2(n2158), .QN(n1654) );
  NAND2X0 U2139 ( .IN1(n1645), .IN2(n1644), .QN(n1648) );
  INVX0 U2140 ( .INP(n1647), .ZN(n1646) );
  INVX0 U2141 ( .INP(n1648), .ZN(n1650) );
  AO221X1 U2142 ( .IN1(n1647), .IN2(n1648), .IN3(n1646), .IN4(n1650), .IN5(
        n2514), .Q(n1653) );
  AO221X1 U2143 ( .IN1(n1651), .IN2(n1650), .IN3(n1649), .IN4(n1648), .IN5(
        n2516), .Q(n1652) );
  NAND4X0 U2144 ( .IN1(n1655), .IN2(n1654), .IN3(n1653), .IN4(n1652), .QN(
        n2601) );
  MUX21X1 U2145 ( .IN1(n1656), .IN2(n2158), .S(n1662), .Q(n2599) );
  NOR2X0 U2146 ( .IN1(n2563), .IN2(n2599), .QN(n1657) );
  AO21X1 U2147 ( .IN1(reg1[10]), .IN2(n2573), .IN3(n1657), .Q(n1658) );
  AO21X1 U2148 ( .IN1(n2565), .IN2(n2601), .IN3(n1658), .Q(n947) );
  INVX0 U2149 ( .INP(n2599), .ZN(n1659) );
  AO22X1 U2150 ( .IN1(n2153), .IN2(n2539), .IN3(n2541), .IN4(n1659), .Q(n1660)
         );
  AO21X1 U2151 ( .IN1(reg2[10]), .IN2(n2558), .IN3(n1660), .Q(n1661) );
  AO21X1 U2152 ( .IN1(n2556), .IN2(n2601), .IN3(n1661), .Q(n979) );
  OA21X1 U2153 ( .IN1(n1663), .IN2(n1666), .IN3(n1662), .Q(n1679) );
  AO21X1 U2154 ( .IN1(n1916), .IN2(n1687), .IN3(n1664), .Q(n1665) );
  MUX21X1 U2155 ( .IN1(n1665), .IN2(n1918), .S(n2528), .Q(n2164) );
  OA22X1 U2156 ( .IN1(n2527), .IN2(n1666), .IN3(n1993), .IN4(n2164), .Q(n1677)
         );
  NAND2X0 U2157 ( .IN1(n1668), .IN2(n1667), .QN(n1671) );
  INVX0 U2158 ( .INP(n1670), .ZN(n1669) );
  INVX0 U2159 ( .INP(n1671), .ZN(n1673) );
  AO221X1 U2160 ( .IN1(n1670), .IN2(n1671), .IN3(n1669), .IN4(n1673), .IN5(
        n2514), .Q(n1676) );
  AO221X1 U2161 ( .IN1(n1674), .IN2(n1673), .IN3(n1672), .IN4(n1671), .IN5(
        n2516), .Q(n1675) );
  NAND3X0 U2162 ( .IN1(n1677), .IN2(n1676), .IN3(n1675), .QN(n1682) );
  AO21X1 U2163 ( .IN1(n2578), .IN2(n1679), .IN3(n1682), .Q(n2598) );
  MUX21X1 U2164 ( .IN1(reg1[9]), .IN2(n2598), .S(n2565), .Q(n948) );
  INVX0 U2165 ( .INP(n1678), .ZN(n2159) );
  AO22X1 U2166 ( .IN1(n2159), .IN2(n2539), .IN3(n2541), .IN4(n1679), .Q(n1680)
         );
  AO21X1 U2167 ( .IN1(reg2[9]), .IN2(n2558), .IN3(n1680), .Q(n1681) );
  AO21X1 U2168 ( .IN1(n2556), .IN2(n1682), .IN3(n1681), .Q(n980) );
  NAND2X0 U2169 ( .IN1(n1684), .IN2(n1683), .QN(n1689) );
  INVX0 U2170 ( .INP(n1686), .ZN(n1685) );
  INVX0 U2171 ( .INP(n1689), .ZN(n1691) );
  AO221X1 U2172 ( .IN1(n1686), .IN2(n1689), .IN3(n1685), .IN4(n1691), .IN5(
        n2514), .Q(n1696) );
  NAND2X0 U2173 ( .IN1(n2485), .IN2(n2180), .QN(n1695) );
  OA21X1 U2174 ( .IN1(n1705), .IN2(n2669), .IN3(n1687), .Q(n1688) );
  MUX21X1 U2175 ( .IN1(n1688), .IN2(n2667), .S(n2528), .Q(n2170) );
  NAND2X0 U2176 ( .IN1(n2529), .IN2(n2170), .QN(n1694) );
  AO221X1 U2177 ( .IN1(n1692), .IN2(n1691), .IN3(n1690), .IN4(n1689), .IN5(
        n2516), .Q(n1693) );
  NAND4X0 U2178 ( .IN1(n1696), .IN2(n1695), .IN3(n1694), .IN4(n1693), .QN(
        n2597) );
  MUX21X1 U2179 ( .IN1(n1697), .IN2(n2180), .S(n1703), .Q(n2595) );
  NOR2X0 U2180 ( .IN1(n2563), .IN2(n2595), .QN(n1698) );
  AO21X1 U2181 ( .IN1(reg1[8]), .IN2(n2573), .IN3(n1698), .Q(n1699) );
  AO21X1 U2182 ( .IN1(n2565), .IN2(n2597), .IN3(n1699), .Q(n949) );
  INVX0 U2183 ( .INP(n2595), .ZN(n1700) );
  AO22X1 U2184 ( .IN1(n2175), .IN2(n2539), .IN3(n2541), .IN4(n1700), .Q(n1701)
         );
  AO21X1 U2185 ( .IN1(reg2[8]), .IN2(n2558), .IN3(n1701), .Q(n1702) );
  AO21X1 U2186 ( .IN1(n2556), .IN2(n2597), .IN3(n1702), .Q(n981) );
  OA21X1 U2187 ( .IN1(n1704), .IN2(n1707), .IN3(n1703), .Q(n1718) );
  AO21X1 U2188 ( .IN1(n1918), .IN2(n1724), .IN3(n1705), .Q(n1706) );
  MUX21X1 U2189 ( .IN1(n1706), .IN2(n1920), .S(n2528), .Q(n2186) );
  OA22X1 U2190 ( .IN1(n2527), .IN2(n1707), .IN3(n1993), .IN4(n2186), .Q(n1716)
         );
  INVX0 U2191 ( .INP(n1709), .ZN(n1708) );
  AO221X1 U2192 ( .IN1(n1709), .IN2(n1710), .IN3(n1708), .IN4(n1712), .IN5(
        n2514), .Q(n1715) );
  AO221X1 U2193 ( .IN1(n1713), .IN2(n1712), .IN3(n1711), .IN4(n1710), .IN5(
        n2516), .Q(n1714) );
  NAND3X0 U2194 ( .IN1(n1716), .IN2(n1715), .IN3(n1714), .QN(n1721) );
  AO21X1 U2195 ( .IN1(n2578), .IN2(n1718), .IN3(n1721), .Q(n2594) );
  MUX21X1 U2196 ( .IN1(reg1[7]), .IN2(n2594), .S(n2565), .Q(n950) );
  INVX0 U2197 ( .INP(n1717), .ZN(n2181) );
  AO22X1 U2198 ( .IN1(n2181), .IN2(n2539), .IN3(n2541), .IN4(n1718), .Q(n1719)
         );
  AO21X1 U2199 ( .IN1(reg2[7]), .IN2(n2558), .IN3(n1719), .Q(n1720) );
  AO21X1 U2200 ( .IN1(n2556), .IN2(n1721), .IN3(n1720), .Q(n982) );
  INVX0 U2201 ( .INP(n1723), .ZN(n1722) );
  AO221X1 U2202 ( .IN1(n1723), .IN2(n1726), .IN3(n1722), .IN4(n1728), .IN5(
        n2514), .Q(n1733) );
  NAND2X0 U2203 ( .IN1(n2485), .IN2(n2202), .QN(n1732) );
  OA21X1 U2204 ( .IN1(n1742), .IN2(n2667), .IN3(n1724), .Q(n1725) );
  MUX21X1 U2205 ( .IN1(n1725), .IN2(n2665), .S(n2528), .Q(n2192) );
  NAND2X0 U2206 ( .IN1(n2529), .IN2(n2192), .QN(n1731) );
  AO221X1 U2207 ( .IN1(n1729), .IN2(n1728), .IN3(n1727), .IN4(n1726), .IN5(
        n2516), .Q(n1730) );
  NAND4X0 U2208 ( .IN1(n1733), .IN2(n1732), .IN3(n1731), .IN4(n1730), .QN(
        n2593) );
  MUX21X1 U2209 ( .IN1(n1734), .IN2(n2202), .S(n1740), .Q(n2591) );
  NOR2X0 U2210 ( .IN1(n2563), .IN2(n2591), .QN(n1735) );
  AO21X1 U2211 ( .IN1(reg1[6]), .IN2(n2573), .IN3(n1735), .Q(n1736) );
  AO21X1 U2212 ( .IN1(n2565), .IN2(n2593), .IN3(n1736), .Q(n951) );
  INVX0 U2213 ( .INP(n2591), .ZN(n1737) );
  AO22X1 U2214 ( .IN1(n2197), .IN2(n2539), .IN3(n2541), .IN4(n1737), .Q(n1738)
         );
  AO21X1 U2215 ( .IN1(reg2[6]), .IN2(n2558), .IN3(n1738), .Q(n1739) );
  AO21X1 U2216 ( .IN1(n2556), .IN2(n2593), .IN3(n1739), .Q(n983) );
  OA21X1 U2217 ( .IN1(n1741), .IN2(n1744), .IN3(n1740), .Q(n1754) );
  AO21X1 U2218 ( .IN1(n1920), .IN2(n1760), .IN3(n1742), .Q(n1743) );
  MUX21X1 U2219 ( .IN1(n1743), .IN2(n1922), .S(n2528), .Q(n2208) );
  OA22X1 U2220 ( .IN1(n2527), .IN2(n1744), .IN3(n1993), .IN4(n2208), .Q(n1753)
         );
  INVX0 U2221 ( .INP(n1746), .ZN(n1745) );
  AO221X1 U2222 ( .IN1(n1746), .IN2(n1747), .IN3(n1745), .IN4(n1749), .IN5(
        n2514), .Q(n1752) );
  AO221X1 U2223 ( .IN1(n1750), .IN2(n1749), .IN3(n1748), .IN4(n1747), .IN5(
        n2516), .Q(n1751) );
  NAND3X0 U2224 ( .IN1(n1753), .IN2(n1752), .IN3(n1751), .QN(n1757) );
  AO21X1 U2225 ( .IN1(n2578), .IN2(n1754), .IN3(n1757), .Q(n2590) );
  MUX21X1 U2226 ( .IN1(reg1[5]), .IN2(n2590), .S(n2565), .Q(n952) );
  AO22X1 U2227 ( .IN1(n2203), .IN2(n2539), .IN3(n2541), .IN4(n1754), .Q(n1755)
         );
  AO21X1 U2228 ( .IN1(reg2[5]), .IN2(n2558), .IN3(n1755), .Q(n1756) );
  AO21X1 U2229 ( .IN1(n2556), .IN2(n1757), .IN3(n1756), .Q(n984) );
  INVX0 U2230 ( .INP(n1764), .ZN(n1762) );
  INVX0 U2231 ( .INP(n1759), .ZN(n1758) );
  AO221X1 U2232 ( .IN1(n1759), .IN2(n1762), .IN3(n1758), .IN4(n1764), .IN5(
        n2514), .Q(n1769) );
  NAND2X0 U2233 ( .IN1(n2485), .IN2(n2228), .QN(n1768) );
  OA21X1 U2234 ( .IN1(n1778), .IN2(n2665), .IN3(n1760), .Q(n1761) );
  MUX21X1 U2235 ( .IN1(n1761), .IN2(n2663), .S(n2528), .Q(n2215) );
  NAND2X0 U2236 ( .IN1(n2529), .IN2(n2215), .QN(n1767) );
  AO221X1 U2237 ( .IN1(n1765), .IN2(n1764), .IN3(n1763), .IN4(n1762), .IN5(
        n2516), .Q(n1766) );
  NAND4X0 U2238 ( .IN1(n1769), .IN2(n1768), .IN3(n1767), .IN4(n1766), .QN(
        n2589) );
  MUX21X1 U2239 ( .IN1(n1770), .IN2(n2228), .S(n1776), .Q(n2587) );
  NOR2X0 U2240 ( .IN1(n2563), .IN2(n2587), .QN(n1771) );
  AO21X1 U2241 ( .IN1(reg1[4]), .IN2(n2573), .IN3(n1771), .Q(n1772) );
  AO21X1 U2242 ( .IN1(n2565), .IN2(n2589), .IN3(n1772), .Q(n953) );
  INVX0 U2243 ( .INP(n2587), .ZN(n1773) );
  AO22X1 U2244 ( .IN1(n2221), .IN2(n2539), .IN3(n2541), .IN4(n1773), .Q(n1774)
         );
  AO21X1 U2245 ( .IN1(reg2[4]), .IN2(n2558), .IN3(n1774), .Q(n1775) );
  AO21X1 U2246 ( .IN1(n2556), .IN2(n2589), .IN3(n1775), .Q(n985) );
  OA21X1 U2247 ( .IN1(n1777), .IN2(n1780), .IN3(n1776), .Q(n1792) );
  AO21X1 U2248 ( .IN1(n1922), .IN2(n1796), .IN3(n1778), .Q(n1779) );
  MUX21X1 U2249 ( .IN1(n1779), .IN2(n1858), .S(n2528), .Q(n1896) );
  OA22X1 U2250 ( .IN1(n2527), .IN2(n1780), .IN3(n1993), .IN4(n1896), .Q(n1791)
         );
  NAND2X0 U2251 ( .IN1(n1782), .IN2(n1781), .QN(n1787) );
  INVX0 U2252 ( .INP(n1787), .ZN(n1785) );
  AO221X1 U2253 ( .IN1(n1784), .IN2(n1785), .IN3(n1783), .IN4(n1787), .IN5(
        n2516), .Q(n1790) );
  INVX0 U2254 ( .INP(n1788), .ZN(n1786) );
  AO221X1 U2255 ( .IN1(n1788), .IN2(n1787), .IN3(n1786), .IN4(n1785), .IN5(
        n2514), .Q(n1789) );
  NAND3X0 U2256 ( .IN1(n1791), .IN2(n1790), .IN3(n1789), .QN(n1795) );
  AO21X1 U2257 ( .IN1(n2578), .IN2(n1792), .IN3(n1795), .Q(n2586) );
  MUX21X1 U2258 ( .IN1(reg1[3]), .IN2(n2586), .S(n2565), .Q(n954) );
  AO22X1 U2259 ( .IN1(n1792), .IN2(n2541), .IN3(n2539), .IN4(n2698), .Q(n1793)
         );
  AO21X1 U2260 ( .IN1(reg2[3]), .IN2(n2558), .IN3(n1793), .Q(n1794) );
  AO21X1 U2261 ( .IN1(n2556), .IN2(n1795), .IN3(n1794), .Q(n986) );
  OA21X1 U2262 ( .IN1(n1814), .IN2(n2663), .IN3(n1796), .Q(n1797) );
  MUX21X1 U2263 ( .IN1(n2661), .IN2(n1797), .S(n1996), .Q(n1857) );
  NAND2X0 U2264 ( .IN1(n2529), .IN2(n1857), .QN(n1809) );
  NAND2X0 U2265 ( .IN1(n2485), .IN2(n1859), .QN(n1808) );
  NAND2X0 U2266 ( .IN1(n1799), .IN2(n1798), .QN(n1802) );
  INVX0 U2267 ( .INP(n1801), .ZN(n1800) );
  INVX0 U2268 ( .INP(n1802), .ZN(n1804) );
  AO221X1 U2269 ( .IN1(n1801), .IN2(n1802), .IN3(n1800), .IN4(n1804), .IN5(
        n2514), .Q(n1807) );
  AO221X1 U2270 ( .IN1(n1805), .IN2(n1804), .IN3(n1803), .IN4(n1802), .IN5(
        n2516), .Q(n1806) );
  NAND4X0 U2271 ( .IN1(n1809), .IN2(n1808), .IN3(n1807), .IN4(n1806), .QN(
        n2585) );
  MUX21X1 U2272 ( .IN1(n1810), .IN2(n1859), .S(n1813), .Q(n2583) );
  NOR2X0 U2273 ( .IN1(n2563), .IN2(n2583), .QN(n1811) );
  AO21X1 U2274 ( .IN1(reg1[2]), .IN2(n2573), .IN3(n1811), .Q(n1812) );
  AO21X1 U2275 ( .IN1(n2565), .IN2(n2585), .IN3(n1812), .Q(n955) );
  OA21X1 U2276 ( .IN1(n2579), .IN2(n1816), .IN3(n1813), .Q(n1853) );
  AO21X1 U2277 ( .IN1(n1858), .IN2(n1872), .IN3(n1814), .Q(n1815) );
  MUX21X1 U2278 ( .IN1(n1815), .IN2(n1838), .S(n2528), .Q(n1841) );
  OA22X1 U2279 ( .IN1(n2527), .IN2(n1816), .IN3(n1993), .IN4(n1841), .Q(n1825)
         );
  AO221X1 U2280 ( .IN1(n1818), .IN2(n1821), .IN3(n1817), .IN4(n1819), .IN5(
        n2516), .Q(n1824) );
  AO221X1 U2281 ( .IN1(n1822), .IN2(n1821), .IN3(n1820), .IN4(n1819), .IN5(
        n2514), .Q(n1823) );
  NAND3X0 U2282 ( .IN1(n1825), .IN2(n1824), .IN3(n1823), .QN(n1856) );
  AO21X1 U2283 ( .IN1(n2578), .IN2(n1853), .IN3(n1856), .Q(n2582) );
  MUX21X1 U2284 ( .IN1(reg1[1]), .IN2(n2582), .S(n2565), .Q(n956) );
  INVX0 U2285 ( .INP(n1826), .ZN(n1829) );
  NAND2X0 U2286 ( .IN1(n2697), .IN2(n2693), .QN(n1827) );
  OA22X1 U2287 ( .IN1(n1828), .IN2(n2709), .IN3(n2575), .IN4(n1827), .Q(n1846)
         );
  AO221X1 U2288 ( .IN1(n1829), .IN2(n2527), .IN3(n1829), .IN4(n1846), .IN5(
        n2391), .Q(n1830) );
  NOR2X0 U2289 ( .IN1(n1830), .IN2(n2703), .QN(n2229) );
  NAND2X0 U2290 ( .IN1(n2229), .IN2(n1837), .QN(n1852) );
  INVX0 U2291 ( .INP(n1909), .ZN(n2570) );
  OA21X1 U2292 ( .IN1(n1832), .IN2(n1831), .IN3(n2570), .Q(n1842) );
  INVX0 U2293 ( .INP(n2661), .ZN(n1833) );
  NOR2X0 U2294 ( .IN1(n2570), .IN2(n1833), .QN(n1862) );
  INVX0 U2295 ( .INP(n2514), .ZN(n1836) );
  INVX0 U2296 ( .INP(n1834), .ZN(n1835) );
  OR2X1 U2297 ( .IN1(n1836), .IN2(n1835), .Q(n1976) );
  XOR2X1 U2298 ( .IN1(n1976), .IN2(n1837), .Q(n1861) );
  NOR2X0 U2299 ( .IN1(n2570), .IN2(n1838), .QN(n1877) );
  XOR2X1 U2300 ( .IN1(n1976), .IN2(n1885), .Q(n1876) );
  NAND2X0 U2301 ( .IN1(n1000), .IN2(n1839), .QN(n1851) );
  NAND3X0 U2302 ( .IN1(n2694), .IN2(n1840), .IN3(n2529), .QN(n1843) );
  NOR3X0 U2303 ( .IN1(n2703), .IN2(n1843), .IN3(n1846), .QN(n2216) );
  INVX0 U2304 ( .INP(n2216), .ZN(n2209) );
  OR2X1 U2305 ( .IN1(n2209), .IN2(n1841), .Q(n1850) );
  INVX0 U2306 ( .INP(n1842), .ZN(n1845) );
  NAND2X0 U2307 ( .IN1(n2527), .IN2(n1843), .QN(n1844) );
  AO22X1 U2308 ( .IN1(n1846), .IN2(n1845), .IN3(n1846), .IN4(n1844), .Q(n1847)
         );
  NOR2X0 U2309 ( .IN1(n1848), .IN2(n1847), .QN(n1890) );
  NAND2X0 U2310 ( .IN1(state), .IN2(n1890), .QN(n1880) );
  NAND2X0 U2311 ( .IN1(n1880), .IN2(reg3[1]), .QN(n1849) );
  NAND4X0 U2312 ( .IN1(n1852), .IN2(n1851), .IN3(n1850), .IN4(n1849), .QN(n804) );
  AO22X1 U2313 ( .IN1(reg3[1]), .IN2(n2539), .IN3(n2541), .IN4(n1853), .Q(
        n1854) );
  AO21X1 U2314 ( .IN1(reg2[1]), .IN2(n2558), .IN3(n1854), .Q(n1855) );
  AO21X1 U2315 ( .IN1(n2556), .IN2(n1856), .IN3(n1855), .Q(n988) );
  NAND2X0 U2316 ( .IN1(n2216), .IN2(n1857), .QN(n1867) );
  NAND2X0 U2317 ( .IN1(n1859), .IN2(n2229), .QN(n1866) );
  NAND2X0 U2318 ( .IN1(n1880), .IN2(reg3[2]), .QN(n1865) );
  NOR2X0 U2319 ( .IN1(n2570), .IN2(n1858), .QN(n1894) );
  XOR2X1 U2320 ( .IN1(n1976), .IN2(n1859), .Q(n1893) );
  FADDX1 U2321 ( .A(n1862), .B(n1861), .CI(n1860), .CO(n1892), .S(n1839) );
  NAND2X0 U2322 ( .IN1(n1000), .IN2(n1863), .QN(n1864) );
  NAND4X0 U2323 ( .IN1(n1867), .IN2(n1866), .IN3(n1865), .IN4(n1864), .QN(n803) );
  INVX0 U2324 ( .INP(n2583), .ZN(n1868) );
  AO22X1 U2325 ( .IN1(reg3[2]), .IN2(n2539), .IN3(n2541), .IN4(n1868), .Q(
        n1869) );
  AO21X1 U2326 ( .IN1(reg2[2]), .IN2(n2558), .IN3(n1869), .Q(n1870) );
  AO21X1 U2327 ( .IN1(n2556), .IN2(n2585), .IN3(n1870), .Q(n987) );
  AO21X1 U2328 ( .IN1(n2660), .IN2(n2692), .IN3(n2661), .Q(n1871) );
  NAND3X0 U2329 ( .IN1(n1996), .IN2(n1872), .IN3(n1871), .QN(n1879) );
  OAI222X1 U2330 ( .IN1(n2579), .IN2(n2527), .IN3(n1873), .IN4(n2570), .IN5(
        n1879), .IN6(n1993), .QN(n2581) );
  INVX0 U2331 ( .INP(n2563), .ZN(n1874) );
  AO22X1 U2332 ( .IN1(reg1[0]), .IN2(n2573), .IN3(n1885), .IN4(n1874), .Q(
        n1875) );
  AO21X1 U2333 ( .IN1(n2565), .IN2(n2581), .IN3(n1875), .Q(n957) );
  NAND2X0 U2334 ( .IN1(n2229), .IN2(n1885), .QN(n1884) );
  FADDX1 U2335 ( .A(n1976), .B(n1877), .CI(n1876), .CO(n1860), .S(n1878) );
  NAND2X0 U2336 ( .IN1(n1000), .IN2(n1878), .QN(n1883) );
  OR2X1 U2337 ( .IN1(n2209), .IN2(n1879), .Q(n1882) );
  NAND2X0 U2338 ( .IN1(n1880), .IN2(reg3[0]), .QN(n1881) );
  NAND4X0 U2339 ( .IN1(n1884), .IN2(n1883), .IN3(n1882), .IN4(n1881), .QN(n805) );
  NAND2X0 U2340 ( .IN1(n2556), .IN2(n2581), .QN(n1889) );
  NAND2X0 U2341 ( .IN1(n2541), .IN2(n1885), .QN(n1888) );
  NAND2X0 U2342 ( .IN1(reg2[0]), .IN2(n2558), .QN(n1887) );
  NAND2X0 U2343 ( .IN1(reg3[0]), .IN2(n2539), .QN(n1886) );
  NAND4X0 U2344 ( .IN1(n1889), .IN2(n1888), .IN3(n1887), .IN4(n1886), .QN(n989) );
  NAND2X0 U2345 ( .IN1(reg3[3]), .IN2(n2703), .QN(n2362) );
  NOR2X0 U2346 ( .IN1(n1890), .IN2(n2703), .QN(n2222) );
  NAND2X0 U2347 ( .IN1(n2222), .IN2(n2698), .QN(n1899) );
  INVX0 U2348 ( .INP(n2663), .ZN(n1891) );
  NOR2X0 U2349 ( .IN1(n2570), .IN2(n1891), .QN(n1925) );
  XOR2X1 U2350 ( .IN1(n1976), .IN2(n1901), .Q(n1924) );
  FADDX1 U2351 ( .A(n1894), .B(n1893), .CI(n1892), .CO(n1923), .S(n1863) );
  NAND2X0 U2352 ( .IN1(n1000), .IN2(n1895), .QN(n1898) );
  OR2X1 U2353 ( .IN1(n2209), .IN2(n1896), .Q(n1897) );
  NAND4X0 U2354 ( .IN1(n2362), .IN2(n1899), .IN3(n1898), .IN4(n1897), .QN(
        n1900) );
  AO21X1 U2355 ( .IN1(n2229), .IN2(n1901), .IN3(n1900), .Q(n802) );
  AOI22X1 U2356 ( .IN1(n2409), .IN2(n2222), .IN3(reg3[20]), .IN4(n2703), .QN(
        n1930) );
  OA21X1 U2357 ( .IN1(n1903), .IN2(n2681), .IN3(n1902), .Q(n1904) );
  MUX21X1 U2358 ( .IN1(n2679), .IN2(n1904), .S(n1996), .Q(n2392) );
  NAND2X0 U2359 ( .IN1(n2216), .IN2(n2392), .QN(n1929) );
  NAND2X0 U2360 ( .IN1(n2229), .IN2(n2406), .QN(n1928) );
  NOR2X0 U2361 ( .IN1(n2570), .IN2(n1905), .QN(n1938) );
  XOR2X1 U2362 ( .IN1(n1976), .IN2(n2406), .Q(n1937) );
  INVX0 U2363 ( .INP(n2679), .ZN(n1906) );
  NOR2X0 U2364 ( .IN1(n2570), .IN2(n1906), .QN(n2052) );
  XOR2X1 U2365 ( .IN1(n1976), .IN2(n2059), .Q(n2051) );
  NOR2X0 U2366 ( .IN1(n2570), .IN2(n1907), .QN(n2063) );
  XOR2X1 U2367 ( .IN1(n1976), .IN2(n2070), .Q(n2062) );
  INVX0 U2368 ( .INP(n2677), .ZN(n1908) );
  NOR2X0 U2369 ( .IN1(n2570), .IN2(n1908), .QN(n2074) );
  XOR2X1 U2370 ( .IN1(n1976), .IN2(n2081), .Q(n2073) );
  NOR2X0 U2371 ( .IN1(n2570), .IN2(n1910), .QN(n2085) );
  XOR2X1 U2372 ( .IN1(n1976), .IN2(n2092), .Q(n2084) );
  INVX0 U2373 ( .INP(n2675), .ZN(n1911) );
  NOR2X0 U2374 ( .IN1(n2570), .IN2(n1911), .QN(n2096) );
  XOR2X1 U2375 ( .IN1(n1976), .IN2(n2103), .Q(n2095) );
  NOR2X0 U2376 ( .IN1(n2570), .IN2(n1912), .QN(n2107) );
  XOR2X1 U2377 ( .IN1(n1976), .IN2(n2114), .Q(n2106) );
  INVX0 U2378 ( .INP(n2673), .ZN(n1913) );
  NOR2X0 U2379 ( .IN1(n2570), .IN2(n1913), .QN(n2118) );
  XOR2X1 U2380 ( .IN1(n1976), .IN2(n2125), .Q(n2117) );
  NOR2X0 U2381 ( .IN1(n2570), .IN2(n1914), .QN(n2129) );
  XOR2X1 U2382 ( .IN1(n1976), .IN2(n2136), .Q(n2128) );
  INVX0 U2383 ( .INP(n2671), .ZN(n1915) );
  NOR2X0 U2384 ( .IN1(n2570), .IN2(n1915), .QN(n2140) );
  XOR2X1 U2385 ( .IN1(n1976), .IN2(n2147), .Q(n2139) );
  NOR2X0 U2386 ( .IN1(n2570), .IN2(n1916), .QN(n2151) );
  XOR2X1 U2387 ( .IN1(n1976), .IN2(n2158), .Q(n2150) );
  INVX0 U2388 ( .INP(n2669), .ZN(n1917) );
  NOR2X0 U2389 ( .IN1(n2570), .IN2(n1917), .QN(n2162) );
  XOR2X1 U2390 ( .IN1(n1976), .IN2(n2169), .Q(n2161) );
  NOR2X0 U2391 ( .IN1(n2570), .IN2(n1918), .QN(n2173) );
  XOR2X1 U2392 ( .IN1(n1976), .IN2(n2180), .Q(n2172) );
  INVX0 U2393 ( .INP(n2667), .ZN(n1919) );
  NOR2X0 U2394 ( .IN1(n2570), .IN2(n1919), .QN(n2184) );
  XOR2X1 U2395 ( .IN1(n1976), .IN2(n2191), .Q(n2183) );
  NOR2X0 U2396 ( .IN1(n2570), .IN2(n1920), .QN(n2195) );
  XOR2X1 U2397 ( .IN1(n1976), .IN2(n2202), .Q(n2194) );
  INVX0 U2398 ( .INP(n2665), .ZN(n1921) );
  NOR2X0 U2399 ( .IN1(n2570), .IN2(n1921), .QN(n2206) );
  XOR2X1 U2400 ( .IN1(n1976), .IN2(n2214), .Q(n2205) );
  NOR2X0 U2401 ( .IN1(n2570), .IN2(n1922), .QN(n2219) );
  XOR2X1 U2402 ( .IN1(n1976), .IN2(n2228), .Q(n2218) );
  FADDX1 U2403 ( .A(n1925), .B(n1924), .CI(n1923), .CO(n2217), .S(n1895) );
  NAND2X0 U2404 ( .IN1(n1000), .IN2(n1926), .QN(n1927) );
  NAND4X0 U2405 ( .IN1(n1930), .IN2(n1929), .IN3(n1928), .IN4(n1927), .QN(n785) );
  AOI22X1 U2406 ( .IN1(n2432), .IN2(n2222), .IN3(reg3[22]), .IN4(n2703), .QN(
        n1943) );
  OA21X1 U2407 ( .IN1(n1932), .IN2(n2684), .IN3(n1931), .Q(n1933) );
  MUX21X1 U2408 ( .IN1(n2681), .IN2(n1933), .S(n1996), .Q(n2415) );
  NAND2X0 U2409 ( .IN1(n2216), .IN2(n2415), .QN(n1942) );
  NAND2X0 U2410 ( .IN1(n2229), .IN2(n2429), .QN(n1941) );
  NOR2X0 U2411 ( .IN1(n2570), .IN2(n1934), .QN(n1951) );
  XOR2X1 U2412 ( .IN1(n1976), .IN2(n2429), .Q(n1950) );
  INVX0 U2413 ( .INP(n2681), .ZN(n1935) );
  NOR2X0 U2414 ( .IN1(n2570), .IN2(n1935), .QN(n2040) );
  XOR2X1 U2415 ( .IN1(n1976), .IN2(n2048), .Q(n2039) );
  FADDX1 U2416 ( .A(n1938), .B(n1937), .CI(n1936), .CO(n2038), .S(n1926) );
  NAND2X0 U2417 ( .IN1(n1000), .IN2(n1939), .QN(n1940) );
  NAND4X0 U2418 ( .IN1(n1943), .IN2(n1942), .IN3(n1941), .IN4(n1940), .QN(n783) );
  AOI22X1 U2419 ( .IN1(n2455), .IN2(n2222), .IN3(reg3[24]), .IN4(n2703), .QN(
        n1956) );
  OA21X1 U2420 ( .IN1(n1945), .IN2(n2686), .IN3(n1944), .Q(n1946) );
  MUX21X1 U2421 ( .IN1(n2684), .IN2(n1946), .S(n1996), .Q(n2438) );
  NAND2X0 U2422 ( .IN1(n2216), .IN2(n2438), .QN(n1955) );
  NAND2X0 U2423 ( .IN1(n2229), .IN2(n2452), .QN(n1954) );
  NOR2X0 U2424 ( .IN1(n2570), .IN2(n1947), .QN(n1964) );
  XOR2X1 U2425 ( .IN1(n1976), .IN2(n2452), .Q(n1963) );
  INVX0 U2426 ( .INP(n2684), .ZN(n1948) );
  NOR2X0 U2427 ( .IN1(n2570), .IN2(n1948), .QN(n2028) );
  XOR2X1 U2428 ( .IN1(n1976), .IN2(n2036), .Q(n2027) );
  FADDX1 U2429 ( .A(n1951), .B(n1950), .CI(n1949), .CO(n2026), .S(n1939) );
  NAND2X0 U2430 ( .IN1(n1000), .IN2(n1952), .QN(n1953) );
  NAND4X0 U2431 ( .IN1(n1956), .IN2(n1955), .IN3(n1954), .IN4(n1953), .QN(n781) );
  AOI22X1 U2432 ( .IN1(n2478), .IN2(n2222), .IN3(reg3[26]), .IN4(n2703), .QN(
        n1969) );
  OA21X1 U2433 ( .IN1(n1958), .IN2(n2688), .IN3(n1957), .Q(n1959) );
  MUX21X1 U2434 ( .IN1(n2686), .IN2(n1959), .S(n1996), .Q(n2461) );
  NAND2X0 U2435 ( .IN1(n2216), .IN2(n2461), .QN(n1968) );
  NAND2X0 U2436 ( .IN1(n2229), .IN2(n2475), .QN(n1967) );
  NOR2X0 U2437 ( .IN1(n2570), .IN2(n1960), .QN(n1975) );
  XOR2X1 U2438 ( .IN1(n1976), .IN2(n2475), .Q(n1974) );
  INVX0 U2439 ( .INP(n2686), .ZN(n1961) );
  NOR2X0 U2440 ( .IN1(n2570), .IN2(n1961), .QN(n2016) );
  XOR2X1 U2441 ( .IN1(n1976), .IN2(n2024), .Q(n2015) );
  FADDX1 U2442 ( .A(n1964), .B(n1963), .CI(n1962), .CO(n2014), .S(n1952) );
  NAND2X0 U2443 ( .IN1(n1000), .IN2(n1965), .QN(n1966) );
  NAND4X0 U2444 ( .IN1(n1969), .IN2(n1968), .IN3(n1967), .IN4(n1966), .QN(n779) );
  AOI22X1 U2445 ( .IN1(n2502), .IN2(n2222), .IN3(reg3[28]), .IN4(n2703), .QN(
        n1986) );
  NAND2X0 U2446 ( .IN1(n1970), .IN2(n2690), .QN(n2517) );
  OA21X1 U2447 ( .IN1(n1970), .IN2(n2690), .IN3(n2517), .Q(n1971) );
  MUX21X1 U2448 ( .IN1(n2688), .IN2(n1971), .S(n1996), .Q(n2484) );
  NAND2X0 U2449 ( .IN1(n2216), .IN2(n2484), .QN(n1985) );
  NAND2X0 U2450 ( .IN1(n2229), .IN2(n2535), .QN(n1984) );
  INVX0 U2451 ( .INP(n2688), .ZN(n1972) );
  NOR2X0 U2452 ( .IN1(n2570), .IN2(n1972), .QN(n2005) );
  XOR2X1 U2453 ( .IN1(n1976), .IN2(n2492), .Q(n2004) );
  FADDX1 U2454 ( .A(n1975), .B(n1974), .CI(n1973), .CO(n2003), .S(n1965) );
  XOR2X1 U2455 ( .IN1(n1976), .IN2(n2535), .Q(n1979) );
  NOR2X0 U2456 ( .IN1(n2570), .IN2(n1977), .QN(n1978) );
  XOR2X1 U2457 ( .IN1(n1979), .IN2(n1978), .Q(n1980) );
  XOR2X1 U2458 ( .IN1(n1981), .IN2(n1980), .Q(n1982) );
  NAND2X0 U2459 ( .IN1(n1000), .IN2(n1982), .QN(n1983) );
  NAND4X0 U2460 ( .IN1(n1986), .IN2(n1985), .IN3(n1984), .IN4(n1983), .QN(n777) );
  OA21X1 U2461 ( .IN1(n1988), .IN2(n2529), .IN3(n1987), .Q(n1995) );
  NOR4X0 U2462 ( .IN1(n1989), .IN2(n1995), .IN3(n2528), .IN4(n2703), .QN(n2384) );
  NAND2X0 U2463 ( .IN1(reg3[4]), .IN2(n2703), .QN(n2226) );
  INVX0 U2464 ( .INP(n1989), .ZN(n2233) );
  OA221X1 U2465 ( .IN1(n1989), .IN2(reg2[0]), .IN3(n2233), .IN4(reg1[0]), 
        .IN5(n2528), .Q(n1990) );
  MUX21X1 U2466 ( .IN1(IR[0]), .IN2(n2702), .S(n1990), .Q(n1991) );
  NAND2X0 U2467 ( .IN1(n2736), .IN2(n1991), .QN(n2369) );
  AOI21X1 U2468 ( .IN1(n1992), .IN2(n2520), .IN3(n2703), .QN(n2389) );
  NAND2X0 U2469 ( .IN1(n1993), .IN2(n2520), .QN(n2390) );
  AND3X1 U2470 ( .IN1(n2389), .IN2(n1994), .IN3(n2390), .Q(n2380) );
  NAND2X0 U2471 ( .IN1(addr[4]), .IN2(n2380), .QN(n2000) );
  OR2X1 U2472 ( .IN1(n1996), .IN2(n1995), .Q(n1997) );
  NOR2X0 U2473 ( .IN1(n2703), .IN2(n1997), .QN(n2383) );
  AO22X1 U2474 ( .IN1(reg1[4]), .IN2(n1989), .IN3(reg2[4]), .IN4(n2233), .Q(
        n2232) );
  AO22X1 U2475 ( .IN1(reg1[3]), .IN2(n1989), .IN3(reg2[3]), .IN4(n2233), .Q(
        n2356) );
  AO22X1 U2476 ( .IN1(reg1[2]), .IN2(n1989), .IN3(reg2[2]), .IN4(n2233), .Q(
        n2364) );
  AO22X1 U2477 ( .IN1(reg1[1]), .IN2(n1989), .IN3(reg2[1]), .IN4(n2233), .Q(
        n2374) );
  AO22X1 U2478 ( .IN1(reg1[0]), .IN2(n1989), .IN3(reg2[0]), .IN4(n2233), .Q(
        n2381) );
  NAND2X0 U2479 ( .IN1(n2383), .IN2(n1998), .QN(n1999) );
  NAND4X0 U2480 ( .IN1(n2226), .IN2(n2369), .IN3(n2000), .IN4(n1999), .QN(
        n2001) );
  AO21X1 U2481 ( .IN1(n2384), .IN2(n2231), .IN3(n2001), .Q(n822) );
  NAND2X0 U2482 ( .IN1(reg3[27]), .IN2(n2703), .QN(n2011) );
  INVX0 U2483 ( .INP(n2002), .ZN(n2481) );
  NAND2X0 U2484 ( .IN1(n2481), .IN2(n2222), .QN(n2010) );
  FADDX1 U2485 ( .A(n2005), .B(n2004), .CI(n2003), .CO(n1981), .S(n2006) );
  NAND2X0 U2486 ( .IN1(n1000), .IN2(n2006), .QN(n2009) );
  OR2X1 U2487 ( .IN1(n2209), .IN2(n2007), .Q(n2008) );
  NAND4X0 U2488 ( .IN1(n2011), .IN2(n2010), .IN3(n2009), .IN4(n2008), .QN(
        n2012) );
  AO21X1 U2489 ( .IN1(n2492), .IN2(n2229), .IN3(n2012), .Q(n778) );
  NAND2X0 U2490 ( .IN1(reg3[25]), .IN2(n2703), .QN(n2022) );
  INVX0 U2491 ( .INP(n2013), .ZN(n2458) );
  NAND2X0 U2492 ( .IN1(n2458), .IN2(n2222), .QN(n2021) );
  FADDX1 U2493 ( .A(n2016), .B(n2015), .CI(n2014), .CO(n1973), .S(n2017) );
  NAND2X0 U2494 ( .IN1(n1000), .IN2(n2017), .QN(n2020) );
  OR2X1 U2495 ( .IN1(n2209), .IN2(n2018), .Q(n2019) );
  NAND4X0 U2496 ( .IN1(n2022), .IN2(n2021), .IN3(n2020), .IN4(n2019), .QN(
        n2023) );
  AO21X1 U2497 ( .IN1(n2024), .IN2(n2229), .IN3(n2023), .Q(n780) );
  NAND2X0 U2498 ( .IN1(reg3[23]), .IN2(n2703), .QN(n2034) );
  INVX0 U2499 ( .INP(n2025), .ZN(n2435) );
  NAND2X0 U2500 ( .IN1(n2435), .IN2(n2222), .QN(n2033) );
  FADDX1 U2501 ( .A(n2028), .B(n2027), .CI(n2026), .CO(n1962), .S(n2029) );
  NAND2X0 U2502 ( .IN1(n1000), .IN2(n2029), .QN(n2032) );
  OR2X1 U2503 ( .IN1(n2209), .IN2(n2030), .Q(n2031) );
  NAND4X0 U2504 ( .IN1(n2034), .IN2(n2033), .IN3(n2032), .IN4(n2031), .QN(
        n2035) );
  AO21X1 U2505 ( .IN1(n2036), .IN2(n2229), .IN3(n2035), .Q(n782) );
  NAND2X0 U2506 ( .IN1(reg3[21]), .IN2(n2703), .QN(n2046) );
  INVX0 U2507 ( .INP(n2037), .ZN(n2412) );
  NAND2X0 U2508 ( .IN1(n2412), .IN2(n2222), .QN(n2045) );
  FADDX1 U2509 ( .A(n2040), .B(n2039), .CI(n2038), .CO(n1949), .S(n2041) );
  NAND2X0 U2510 ( .IN1(n1000), .IN2(n2041), .QN(n2044) );
  OR2X1 U2511 ( .IN1(n2209), .IN2(n2042), .Q(n2043) );
  NAND4X0 U2512 ( .IN1(n2046), .IN2(n2045), .IN3(n2044), .IN4(n2043), .QN(
        n2047) );
  AO21X1 U2513 ( .IN1(n2048), .IN2(n2229), .IN3(n2047), .Q(n784) );
  NAND2X0 U2514 ( .IN1(reg3[19]), .IN2(n2703), .QN(n2242) );
  NAND2X0 U2515 ( .IN1(n2049), .IN2(n2222), .QN(n2057) );
  FADDX1 U2516 ( .A(n2052), .B(n2051), .CI(n2050), .CO(n1936), .S(n2053) );
  NAND2X0 U2517 ( .IN1(n1000), .IN2(n2053), .QN(n2056) );
  OR2X1 U2518 ( .IN1(n2209), .IN2(n2054), .Q(n2055) );
  NAND4X0 U2519 ( .IN1(n2242), .IN2(n2057), .IN3(n2056), .IN4(n2055), .QN(
        n2058) );
  AO21X1 U2520 ( .IN1(n2059), .IN2(n2229), .IN3(n2058), .Q(n786) );
  NAND2X0 U2521 ( .IN1(reg3[18]), .IN2(n2703), .QN(n2250) );
  NAND2X0 U2522 ( .IN1(n2060), .IN2(n2216), .QN(n2068) );
  FADDX1 U2523 ( .A(n2063), .B(n2062), .CI(n2061), .CO(n2050), .S(n2064) );
  NAND2X0 U2524 ( .IN1(n1000), .IN2(n2064), .QN(n2067) );
  NAND2X0 U2525 ( .IN1(n2222), .IN2(n2065), .QN(n2066) );
  NAND4X0 U2526 ( .IN1(n2250), .IN2(n2068), .IN3(n2067), .IN4(n2066), .QN(
        n2069) );
  AO21X1 U2527 ( .IN1(n2070), .IN2(n2229), .IN3(n2069), .Q(n787) );
  NAND2X0 U2528 ( .IN1(reg3[17]), .IN2(n2703), .QN(n2258) );
  NAND2X0 U2529 ( .IN1(n2071), .IN2(n2222), .QN(n2079) );
  FADDX1 U2530 ( .A(n2074), .B(n2073), .CI(n2072), .CO(n2061), .S(n2075) );
  NAND2X0 U2531 ( .IN1(n1000), .IN2(n2075), .QN(n2078) );
  OR2X1 U2532 ( .IN1(n2209), .IN2(n2076), .Q(n2077) );
  NAND4X0 U2533 ( .IN1(n2258), .IN2(n2079), .IN3(n2078), .IN4(n2077), .QN(
        n2080) );
  AO21X1 U2534 ( .IN1(n2229), .IN2(n2081), .IN3(n2080), .Q(n788) );
  NAND2X0 U2535 ( .IN1(reg3[16]), .IN2(n2703), .QN(n2266) );
  NAND2X0 U2536 ( .IN1(n2082), .IN2(n2216), .QN(n2090) );
  FADDX1 U2537 ( .A(n2085), .B(n2084), .CI(n2083), .CO(n2072), .S(n2086) );
  NAND2X0 U2538 ( .IN1(n1000), .IN2(n2086), .QN(n2089) );
  NAND2X0 U2539 ( .IN1(n2222), .IN2(n2087), .QN(n2088) );
  NAND4X0 U2540 ( .IN1(n2266), .IN2(n2090), .IN3(n2089), .IN4(n2088), .QN(
        n2091) );
  AO21X1 U2541 ( .IN1(n2229), .IN2(n2092), .IN3(n2091), .Q(n789) );
  NAND2X0 U2542 ( .IN1(reg3[15]), .IN2(n2703), .QN(n2274) );
  NAND2X0 U2543 ( .IN1(n2093), .IN2(n2222), .QN(n2101) );
  FADDX1 U2544 ( .A(n2096), .B(n2095), .CI(n2094), .CO(n2083), .S(n2097) );
  NAND2X0 U2545 ( .IN1(n1000), .IN2(n2097), .QN(n2100) );
  OR2X1 U2546 ( .IN1(n2209), .IN2(n2098), .Q(n2099) );
  NAND4X0 U2547 ( .IN1(n2274), .IN2(n2101), .IN3(n2100), .IN4(n2099), .QN(
        n2102) );
  AO21X1 U2548 ( .IN1(n2229), .IN2(n2103), .IN3(n2102), .Q(n790) );
  NAND2X0 U2549 ( .IN1(reg3[14]), .IN2(n2703), .QN(n2282) );
  NAND2X0 U2550 ( .IN1(n2104), .IN2(n2216), .QN(n2112) );
  FADDX1 U2551 ( .A(n2107), .B(n2106), .CI(n2105), .CO(n2094), .S(n2108) );
  NAND2X0 U2552 ( .IN1(n1000), .IN2(n2108), .QN(n2111) );
  NAND2X0 U2553 ( .IN1(n2222), .IN2(n2109), .QN(n2110) );
  NAND4X0 U2554 ( .IN1(n2282), .IN2(n2112), .IN3(n2111), .IN4(n2110), .QN(
        n2113) );
  AO21X1 U2555 ( .IN1(n2229), .IN2(n2114), .IN3(n2113), .Q(n791) );
  NAND2X0 U2556 ( .IN1(reg3[13]), .IN2(n2703), .QN(n2290) );
  NAND2X0 U2557 ( .IN1(n2115), .IN2(n2222), .QN(n2123) );
  FADDX1 U2558 ( .A(n2118), .B(n2117), .CI(n2116), .CO(n2105), .S(n2119) );
  NAND2X0 U2559 ( .IN1(n1000), .IN2(n2119), .QN(n2122) );
  OR2X1 U2560 ( .IN1(n2209), .IN2(n2120), .Q(n2121) );
  NAND4X0 U2561 ( .IN1(n2290), .IN2(n2123), .IN3(n2122), .IN4(n2121), .QN(
        n2124) );
  AO21X1 U2562 ( .IN1(n2229), .IN2(n2125), .IN3(n2124), .Q(n792) );
  NAND2X0 U2563 ( .IN1(reg3[12]), .IN2(n2703), .QN(n2298) );
  NAND2X0 U2564 ( .IN1(n2126), .IN2(n2216), .QN(n2134) );
  FADDX1 U2565 ( .A(n2129), .B(n2128), .CI(n2127), .CO(n2116), .S(n2130) );
  NAND2X0 U2566 ( .IN1(n1000), .IN2(n2130), .QN(n2133) );
  NAND2X0 U2567 ( .IN1(n2222), .IN2(n2131), .QN(n2132) );
  NAND4X0 U2568 ( .IN1(n2298), .IN2(n2134), .IN3(n2133), .IN4(n2132), .QN(
        n2135) );
  AO21X1 U2569 ( .IN1(n2229), .IN2(n2136), .IN3(n2135), .Q(n793) );
  NAND2X0 U2570 ( .IN1(reg3[11]), .IN2(n2703), .QN(n2306) );
  NAND2X0 U2571 ( .IN1(n2137), .IN2(n2222), .QN(n2145) );
  FADDX1 U2572 ( .A(n2140), .B(n2139), .CI(n2138), .CO(n2127), .S(n2141) );
  NAND2X0 U2573 ( .IN1(n1000), .IN2(n2141), .QN(n2144) );
  OR2X1 U2574 ( .IN1(n2209), .IN2(n2142), .Q(n2143) );
  NAND4X0 U2575 ( .IN1(n2306), .IN2(n2145), .IN3(n2144), .IN4(n2143), .QN(
        n2146) );
  AO21X1 U2576 ( .IN1(n2229), .IN2(n2147), .IN3(n2146), .Q(n794) );
  NAND2X0 U2577 ( .IN1(reg3[10]), .IN2(n2703), .QN(n2314) );
  NAND2X0 U2578 ( .IN1(n2216), .IN2(n2148), .QN(n2156) );
  FADDX1 U2579 ( .A(n2151), .B(n2150), .CI(n2149), .CO(n2138), .S(n2152) );
  NAND2X0 U2580 ( .IN1(n1000), .IN2(n2152), .QN(n2155) );
  NAND2X0 U2581 ( .IN1(n2222), .IN2(n2153), .QN(n2154) );
  NAND4X0 U2582 ( .IN1(n2314), .IN2(n2156), .IN3(n2155), .IN4(n2154), .QN(
        n2157) );
  AO21X1 U2583 ( .IN1(n2229), .IN2(n2158), .IN3(n2157), .Q(n795) );
  NAND2X0 U2584 ( .IN1(reg3[9]), .IN2(n2703), .QN(n2322) );
  NAND2X0 U2585 ( .IN1(n2159), .IN2(n2222), .QN(n2167) );
  FADDX1 U2586 ( .A(n2162), .B(n2161), .CI(n2160), .CO(n2149), .S(n2163) );
  NAND2X0 U2587 ( .IN1(n1000), .IN2(n2163), .QN(n2166) );
  OR2X1 U2588 ( .IN1(n2209), .IN2(n2164), .Q(n2165) );
  NAND4X0 U2589 ( .IN1(n2322), .IN2(n2167), .IN3(n2166), .IN4(n2165), .QN(
        n2168) );
  AO21X1 U2590 ( .IN1(n2229), .IN2(n2169), .IN3(n2168), .Q(n796) );
  NAND2X0 U2591 ( .IN1(reg3[8]), .IN2(n2703), .QN(n2330) );
  NAND2X0 U2592 ( .IN1(n2216), .IN2(n2170), .QN(n2178) );
  FADDX1 U2593 ( .A(n2173), .B(n2172), .CI(n2171), .CO(n2160), .S(n2174) );
  NAND2X0 U2594 ( .IN1(n1000), .IN2(n2174), .QN(n2177) );
  NAND2X0 U2595 ( .IN1(n2222), .IN2(n2175), .QN(n2176) );
  NAND4X0 U2596 ( .IN1(n2330), .IN2(n2178), .IN3(n2177), .IN4(n2176), .QN(
        n2179) );
  AO21X1 U2597 ( .IN1(n2229), .IN2(n2180), .IN3(n2179), .Q(n797) );
  NAND2X0 U2598 ( .IN1(reg3[7]), .IN2(n2703), .QN(n2338) );
  NAND2X0 U2599 ( .IN1(n2181), .IN2(n2222), .QN(n2189) );
  FADDX1 U2600 ( .A(n2184), .B(n2183), .CI(n2182), .CO(n2171), .S(n2185) );
  NAND2X0 U2601 ( .IN1(n1000), .IN2(n2185), .QN(n2188) );
  OR2X1 U2602 ( .IN1(n2209), .IN2(n2186), .Q(n2187) );
  NAND4X0 U2603 ( .IN1(n2338), .IN2(n2189), .IN3(n2188), .IN4(n2187), .QN(
        n2190) );
  AO21X1 U2604 ( .IN1(n2229), .IN2(n2191), .IN3(n2190), .Q(n798) );
  NAND2X0 U2605 ( .IN1(reg3[6]), .IN2(n2703), .QN(n2346) );
  NAND2X0 U2606 ( .IN1(n2216), .IN2(n2192), .QN(n2200) );
  FADDX1 U2607 ( .A(n2195), .B(n2194), .CI(n2193), .CO(n2182), .S(n2196) );
  NAND2X0 U2608 ( .IN1(n1000), .IN2(n2196), .QN(n2199) );
  NAND2X0 U2609 ( .IN1(n2222), .IN2(n2197), .QN(n2198) );
  NAND4X0 U2610 ( .IN1(n2346), .IN2(n2200), .IN3(n2199), .IN4(n2198), .QN(
        n2201) );
  AO21X1 U2611 ( .IN1(n2229), .IN2(n2202), .IN3(n2201), .Q(n799) );
  NAND2X0 U2612 ( .IN1(reg3[5]), .IN2(n2703), .QN(n2354) );
  NAND2X0 U2613 ( .IN1(n2203), .IN2(n2222), .QN(n2212) );
  FADDX1 U2614 ( .A(n2206), .B(n2205), .CI(n2204), .CO(n2193), .S(n2207) );
  NAND2X0 U2615 ( .IN1(n1000), .IN2(n2207), .QN(n2211) );
  OR2X1 U2616 ( .IN1(n2209), .IN2(n2208), .Q(n2210) );
  NAND4X0 U2617 ( .IN1(n2354), .IN2(n2212), .IN3(n2211), .IN4(n2210), .QN(
        n2213) );
  AO21X1 U2618 ( .IN1(n2229), .IN2(n2214), .IN3(n2213), .Q(n800) );
  NAND2X0 U2619 ( .IN1(n2216), .IN2(n2215), .QN(n2225) );
  FADDX1 U2620 ( .A(n2219), .B(n2218), .CI(n2217), .CO(n2204), .S(n2220) );
  NAND2X0 U2621 ( .IN1(n1000), .IN2(n2220), .QN(n2224) );
  NAND2X0 U2622 ( .IN1(n2222), .IN2(n2221), .QN(n2223) );
  NAND4X0 U2623 ( .IN1(n2226), .IN2(n2225), .IN3(n2224), .IN4(n2223), .QN(
        n2227) );
  AO21X1 U2624 ( .IN1(n2229), .IN2(n2228), .IN3(n2227), .Q(n801) );
  NAND2X0 U2625 ( .IN1(n2380), .IN2(addr[19]), .QN(n2241) );
  AO22X1 U2626 ( .IN1(reg1[18]), .IN2(n1989), .IN3(reg2[18]), .IN4(n2233), .Q(
        n2244) );
  AO22X1 U2627 ( .IN1(reg1[17]), .IN2(n1989), .IN3(reg2[17]), .IN4(n2233), .Q(
        n2252) );
  AO22X1 U2628 ( .IN1(reg1[16]), .IN2(n1989), .IN3(reg2[16]), .IN4(n2233), .Q(
        n2260) );
  AO22X1 U2629 ( .IN1(reg1[15]), .IN2(n1989), .IN3(reg2[15]), .IN4(n2233), .Q(
        n2268) );
  AO22X1 U2630 ( .IN1(reg1[14]), .IN2(n1989), .IN3(reg2[14]), .IN4(n2233), .Q(
        n2276) );
  AO22X1 U2631 ( .IN1(reg1[13]), .IN2(n1989), .IN3(reg2[13]), .IN4(n2233), .Q(
        n2284) );
  AO22X1 U2632 ( .IN1(reg1[12]), .IN2(n1989), .IN3(reg2[12]), .IN4(n2233), .Q(
        n2292) );
  AO22X1 U2633 ( .IN1(reg1[11]), .IN2(n1989), .IN3(reg2[11]), .IN4(n2233), .Q(
        n2300) );
  AO22X1 U2634 ( .IN1(reg1[10]), .IN2(n1989), .IN3(reg2[10]), .IN4(n2233), .Q(
        n2308) );
  AO22X1 U2635 ( .IN1(reg1[9]), .IN2(n1989), .IN3(reg2[9]), .IN4(n2233), .Q(
        n2316) );
  AO22X1 U2636 ( .IN1(reg1[8]), .IN2(n1989), .IN3(reg2[8]), .IN4(n2233), .Q(
        n2324) );
  AO22X1 U2637 ( .IN1(reg1[7]), .IN2(n1989), .IN3(reg2[7]), .IN4(n2233), .Q(
        n2332) );
  AO22X1 U2638 ( .IN1(reg1[6]), .IN2(n1989), .IN3(reg2[6]), .IN4(n2233), .Q(
        n2340) );
  AO22X1 U2639 ( .IN1(reg1[5]), .IN2(n1989), .IN3(reg2[5]), .IN4(n2233), .Q(
        n2348) );
  FADDX1 U2640 ( .A(n2232), .B(n2231), .CI(n2230), .CO(n2347), .S(n1998) );
  AO22X1 U2641 ( .IN1(reg1[19]), .IN2(n1989), .IN3(reg2[19]), .IN4(n2233), .Q(
        n2234) );
  XOR2X1 U2642 ( .IN1(n2238), .IN2(n2234), .Q(n2235) );
  XOR2X1 U2643 ( .IN1(n2236), .IN2(n2235), .Q(n2237) );
  NAND2X0 U2644 ( .IN1(n2383), .IN2(n2237), .QN(n2240) );
  NAND2X0 U2645 ( .IN1(n2238), .IN2(n2384), .QN(n2239) );
  NAND4X0 U2646 ( .IN1(n2242), .IN2(n2241), .IN3(n2240), .IN4(n2239), .QN(n806) );
  NAND2X0 U2647 ( .IN1(n2380), .IN2(addr[18]), .QN(n2249) );
  FADDX1 U2648 ( .A(n2244), .B(n2246), .CI(n2243), .CO(n2236), .S(n2245) );
  NAND2X0 U2649 ( .IN1(n2383), .IN2(n2245), .QN(n2248) );
  NAND2X0 U2650 ( .IN1(n2384), .IN2(n2246), .QN(n2247) );
  NAND4X0 U2651 ( .IN1(n2250), .IN2(n2249), .IN3(n2248), .IN4(n2247), .QN(n808) );
  NAND2X0 U2652 ( .IN1(n2380), .IN2(addr[17]), .QN(n2257) );
  FADDX1 U2653 ( .A(n2252), .B(n2254), .CI(n2251), .CO(n2243), .S(n2253) );
  NAND2X0 U2654 ( .IN1(n2383), .IN2(n2253), .QN(n2256) );
  NAND2X0 U2655 ( .IN1(n2384), .IN2(n2254), .QN(n2255) );
  NAND4X0 U2656 ( .IN1(n2258), .IN2(n2257), .IN3(n2256), .IN4(n2255), .QN(n809) );
  NAND2X0 U2657 ( .IN1(n2380), .IN2(addr[16]), .QN(n2265) );
  FADDX1 U2658 ( .A(n2260), .B(n2262), .CI(n2259), .CO(n2251), .S(n2261) );
  NAND2X0 U2659 ( .IN1(n2383), .IN2(n2261), .QN(n2264) );
  NAND2X0 U2660 ( .IN1(n2384), .IN2(n2262), .QN(n2263) );
  NAND4X0 U2661 ( .IN1(n2266), .IN2(n2265), .IN3(n2264), .IN4(n2263), .QN(n810) );
  NAND2X0 U2662 ( .IN1(n2380), .IN2(addr[15]), .QN(n2273) );
  FADDX1 U2663 ( .A(n2268), .B(n2270), .CI(n2267), .CO(n2259), .S(n2269) );
  NAND2X0 U2664 ( .IN1(n2383), .IN2(n2269), .QN(n2272) );
  NAND2X0 U2665 ( .IN1(n2384), .IN2(n2270), .QN(n2271) );
  NAND4X0 U2666 ( .IN1(n2274), .IN2(n2273), .IN3(n2272), .IN4(n2271), .QN(n811) );
  NAND2X0 U2667 ( .IN1(n2380), .IN2(addr[14]), .QN(n2281) );
  FADDX1 U2668 ( .A(n2276), .B(n2278), .CI(n2275), .CO(n2267), .S(n2277) );
  NAND2X0 U2669 ( .IN1(n2383), .IN2(n2277), .QN(n2280) );
  NAND2X0 U2670 ( .IN1(n2384), .IN2(n2278), .QN(n2279) );
  NAND4X0 U2671 ( .IN1(n2282), .IN2(n2281), .IN3(n2280), .IN4(n2279), .QN(n812) );
  NAND2X0 U2672 ( .IN1(n2380), .IN2(addr[13]), .QN(n2289) );
  FADDX1 U2673 ( .A(n2284), .B(n2286), .CI(n2283), .CO(n2275), .S(n2285) );
  NAND2X0 U2674 ( .IN1(n2383), .IN2(n2285), .QN(n2288) );
  NAND2X0 U2675 ( .IN1(n2384), .IN2(n2286), .QN(n2287) );
  NAND4X0 U2676 ( .IN1(n2290), .IN2(n2289), .IN3(n2288), .IN4(n2287), .QN(n813) );
  NAND2X0 U2677 ( .IN1(n2380), .IN2(addr[12]), .QN(n2297) );
  FADDX1 U2678 ( .A(n2292), .B(n2294), .CI(n2291), .CO(n2283), .S(n2293) );
  NAND2X0 U2679 ( .IN1(n2383), .IN2(n2293), .QN(n2296) );
  NAND2X0 U2680 ( .IN1(n2384), .IN2(n2294), .QN(n2295) );
  NAND4X0 U2681 ( .IN1(n2298), .IN2(n2297), .IN3(n2296), .IN4(n2295), .QN(n814) );
  NAND2X0 U2682 ( .IN1(n2380), .IN2(addr[11]), .QN(n2305) );
  FADDX1 U2683 ( .A(n2300), .B(n2302), .CI(n2299), .CO(n2291), .S(n2301) );
  NAND2X0 U2684 ( .IN1(n2383), .IN2(n2301), .QN(n2304) );
  NAND2X0 U2685 ( .IN1(n2384), .IN2(n2302), .QN(n2303) );
  NAND4X0 U2686 ( .IN1(n2306), .IN2(n2305), .IN3(n2304), .IN4(n2303), .QN(n815) );
  NAND2X0 U2687 ( .IN1(n2380), .IN2(addr[10]), .QN(n2313) );
  FADDX1 U2688 ( .A(n2308), .B(n2310), .CI(n2307), .CO(n2299), .S(n2309) );
  NAND2X0 U2689 ( .IN1(n2383), .IN2(n2309), .QN(n2312) );
  NAND2X0 U2690 ( .IN1(n2384), .IN2(n2310), .QN(n2311) );
  NAND4X0 U2691 ( .IN1(n2314), .IN2(n2313), .IN3(n2312), .IN4(n2311), .QN(n816) );
  NAND2X0 U2692 ( .IN1(n2380), .IN2(addr[9]), .QN(n2321) );
  FADDX1 U2693 ( .A(n2316), .B(n2318), .CI(n2315), .CO(n2307), .S(n2317) );
  NAND2X0 U2694 ( .IN1(n2383), .IN2(n2317), .QN(n2320) );
  NAND2X0 U2695 ( .IN1(n2384), .IN2(n2318), .QN(n2319) );
  NAND4X0 U2696 ( .IN1(n2322), .IN2(n2321), .IN3(n2320), .IN4(n2319), .QN(n817) );
  NAND2X0 U2697 ( .IN1(n2380), .IN2(addr[8]), .QN(n2329) );
  FADDX1 U2698 ( .A(n2324), .B(n2326), .CI(n2323), .CO(n2315), .S(n2325) );
  NAND2X0 U2699 ( .IN1(n2383), .IN2(n2325), .QN(n2328) );
  NAND2X0 U2700 ( .IN1(n2384), .IN2(n2326), .QN(n2327) );
  NAND4X0 U2701 ( .IN1(n2330), .IN2(n2329), .IN3(n2328), .IN4(n2327), .QN(n818) );
  NAND2X0 U2702 ( .IN1(n2380), .IN2(addr[7]), .QN(n2337) );
  FADDX1 U2703 ( .A(n2332), .B(n2334), .CI(n2331), .CO(n2323), .S(n2333) );
  NAND2X0 U2704 ( .IN1(n2383), .IN2(n2333), .QN(n2336) );
  NAND2X0 U2705 ( .IN1(n2384), .IN2(n2334), .QN(n2335) );
  NAND4X0 U2706 ( .IN1(n2338), .IN2(n2337), .IN3(n2336), .IN4(n2335), .QN(n819) );
  NAND2X0 U2707 ( .IN1(n2380), .IN2(addr[6]), .QN(n2345) );
  FADDX1 U2708 ( .A(n2340), .B(n2342), .CI(n2339), .CO(n2331), .S(n2341) );
  NAND2X0 U2709 ( .IN1(n2383), .IN2(n2341), .QN(n2344) );
  NAND2X0 U2710 ( .IN1(n2384), .IN2(n2342), .QN(n2343) );
  NAND4X0 U2711 ( .IN1(n2346), .IN2(n2345), .IN3(n2344), .IN4(n2343), .QN(n820) );
  NAND2X0 U2712 ( .IN1(n2380), .IN2(addr[5]), .QN(n2353) );
  FADDX1 U2713 ( .A(n2348), .B(n2350), .CI(n2347), .CO(n2339), .S(n2349) );
  NAND2X0 U2714 ( .IN1(n2383), .IN2(n2349), .QN(n2352) );
  NAND2X0 U2715 ( .IN1(n2384), .IN2(n2350), .QN(n2351) );
  NAND4X0 U2716 ( .IN1(n2354), .IN2(n2353), .IN3(n2352), .IN4(n2351), .QN(n821) );
  NAND2X0 U2717 ( .IN1(n2380), .IN2(addr[3]), .QN(n2361) );
  FADDX1 U2718 ( .A(n2356), .B(n2358), .CI(n2355), .CO(n2230), .S(n2357) );
  NAND2X0 U2719 ( .IN1(n2383), .IN2(n2357), .QN(n2360) );
  NAND2X0 U2720 ( .IN1(n2384), .IN2(n2358), .QN(n2359) );
  NAND4X0 U2721 ( .IN1(n2362), .IN2(n2361), .IN3(n2360), .IN4(n2359), .QN(n823) );
  NAND2X0 U2722 ( .IN1(n2380), .IN2(addr[2]), .QN(n2368) );
  NAND2X0 U2723 ( .IN1(reg3[2]), .IN2(n2703), .QN(n2367) );
  FADDX1 U2724 ( .A(n2364), .B(n2371), .CI(n2363), .CO(n2355), .S(n2365) );
  NAND2X0 U2725 ( .IN1(n2383), .IN2(n2365), .QN(n2366) );
  NAND4X0 U2726 ( .IN1(n2369), .IN2(n2368), .IN3(n2367), .IN4(n2366), .QN(
        n2370) );
  AO21X1 U2727 ( .IN1(n2384), .IN2(n2371), .IN3(n2370), .Q(n824) );
  NAND2X0 U2728 ( .IN1(reg3[1]), .IN2(n2703), .QN(n2379) );
  NAND2X0 U2729 ( .IN1(n2380), .IN2(addr[1]), .QN(n2378) );
  NAND2X0 U2730 ( .IN1(n2384), .IN2(n2373), .QN(n2377) );
  FADDX1 U2731 ( .A(n2374), .B(n2373), .CI(n2372), .CO(n2363), .S(n2375) );
  NAND2X0 U2732 ( .IN1(n2383), .IN2(n2375), .QN(n2376) );
  NAND4X0 U2733 ( .IN1(n2379), .IN2(n2378), .IN3(n2377), .IN4(n2376), .QN(n825) );
  NAND2X0 U2734 ( .IN1(reg3[0]), .IN2(n2703), .QN(n2388) );
  NAND2X0 U2735 ( .IN1(n2380), .IN2(addr[0]), .QN(n2387) );
  HADDX1 U2736 ( .A0(IR[0]), .B0(n2381), .C1(n2372), .SO(n2382) );
  NAND2X0 U2737 ( .IN1(n2383), .IN2(n2382), .QN(n2386) );
  NAND2X0 U2738 ( .IN1(n2384), .IN2(IR[0]), .QN(n2385) );
  NAND4X0 U2739 ( .IN1(n2388), .IN2(n2387), .IN3(n2386), .IN4(n2385), .QN(n826) );
  OAI21X1 U2740 ( .IN1(n2391), .IN2(n2390), .IN3(n2389), .QN(N5560) );
  NAND2X0 U2741 ( .IN1(n2529), .IN2(n2392), .QN(n2404) );
  NAND2X0 U2742 ( .IN1(n2485), .IN2(n2406), .QN(n2403) );
  NAND2X0 U2743 ( .IN1(n2394), .IN2(n2393), .QN(n2397) );
  INVX0 U2744 ( .INP(n2396), .ZN(n2395) );
  INVX0 U2745 ( .INP(n2397), .ZN(n2399) );
  AO221X1 U2746 ( .IN1(n2396), .IN2(n2397), .IN3(n2395), .IN4(n2399), .IN5(
        n2514), .Q(n2402) );
  AO221X1 U2747 ( .IN1(n2400), .IN2(n2399), .IN3(n2398), .IN4(n2397), .IN5(
        n2516), .Q(n2401) );
  NAND4X0 U2748 ( .IN1(n2404), .IN2(n2403), .IN3(n2402), .IN4(n2401), .QN(
        n2621) );
  MUX21X1 U2749 ( .IN1(n2407), .IN2(n2406), .S(n2405), .Q(n2619) );
  INVX0 U2750 ( .INP(n2619), .ZN(n2408) );
  AO22X1 U2751 ( .IN1(n2409), .IN2(n2539), .IN3(n2541), .IN4(n2408), .Q(n2410)
         );
  AO221X1 U2752 ( .IN1(n2556), .IN2(n2621), .IN3(n2558), .IN4(reg2[20]), .IN5(
        n2410), .Q(n969) );
  AO22X1 U2753 ( .IN1(n2412), .IN2(n2539), .IN3(n2541), .IN4(n2411), .Q(n2413)
         );
  AO221X1 U2754 ( .IN1(n2556), .IN2(n2414), .IN3(n2558), .IN4(reg2[21]), .IN5(
        n2413), .Q(n968) );
  NAND2X0 U2755 ( .IN1(n2529), .IN2(n2415), .QN(n2427) );
  NAND2X0 U2756 ( .IN1(n2485), .IN2(n2429), .QN(n2426) );
  NAND2X0 U2757 ( .IN1(n2417), .IN2(n2416), .QN(n2420) );
  INVX0 U2758 ( .INP(n2419), .ZN(n2418) );
  INVX0 U2759 ( .INP(n2420), .ZN(n2422) );
  AO221X1 U2760 ( .IN1(n2419), .IN2(n2420), .IN3(n2418), .IN4(n2422), .IN5(
        n2514), .Q(n2425) );
  AO221X1 U2761 ( .IN1(n2423), .IN2(n2422), .IN3(n2421), .IN4(n2420), .IN5(
        n2516), .Q(n2424) );
  NAND4X0 U2762 ( .IN1(n2427), .IN2(n2426), .IN3(n2425), .IN4(n2424), .QN(
        n2625) );
  MUX21X1 U2763 ( .IN1(n2430), .IN2(n2429), .S(n2428), .Q(n2623) );
  INVX0 U2764 ( .INP(n2623), .ZN(n2431) );
  AO22X1 U2765 ( .IN1(n2432), .IN2(n2539), .IN3(n2541), .IN4(n2431), .Q(n2433)
         );
  AO221X1 U2766 ( .IN1(n2556), .IN2(n2625), .IN3(n2558), .IN4(reg2[22]), .IN5(
        n2433), .Q(n967) );
  AO22X1 U2767 ( .IN1(n2435), .IN2(n2539), .IN3(n2541), .IN4(n2434), .Q(n2436)
         );
  AO221X1 U2768 ( .IN1(n2556), .IN2(n2437), .IN3(n2558), .IN4(reg2[23]), .IN5(
        n2436), .Q(n966) );
  NAND2X0 U2769 ( .IN1(n2529), .IN2(n2438), .QN(n2450) );
  NAND2X0 U2770 ( .IN1(n2485), .IN2(n2452), .QN(n2449) );
  NAND2X0 U2771 ( .IN1(n2440), .IN2(n2439), .QN(n2443) );
  INVX0 U2772 ( .INP(n2442), .ZN(n2441) );
  INVX0 U2773 ( .INP(n2443), .ZN(n2445) );
  AO221X1 U2774 ( .IN1(n2442), .IN2(n2443), .IN3(n2441), .IN4(n2445), .IN5(
        n2514), .Q(n2448) );
  AO221X1 U2775 ( .IN1(n2446), .IN2(n2445), .IN3(n2444), .IN4(n2443), .IN5(
        n2516), .Q(n2447) );
  NAND4X0 U2776 ( .IN1(n2450), .IN2(n2449), .IN3(n2448), .IN4(n2447), .QN(
        n2629) );
  MUX21X1 U2777 ( .IN1(n2453), .IN2(n2452), .S(n2451), .Q(n2627) );
  INVX0 U2778 ( .INP(n2627), .ZN(n2454) );
  AO22X1 U2779 ( .IN1(n2455), .IN2(n2539), .IN3(n2541), .IN4(n2454), .Q(n2456)
         );
  AO221X1 U2780 ( .IN1(n2556), .IN2(n2629), .IN3(n2558), .IN4(reg2[24]), .IN5(
        n2456), .Q(n965) );
  AO22X1 U2781 ( .IN1(n2458), .IN2(n2539), .IN3(n2541), .IN4(n2457), .Q(n2459)
         );
  AO221X1 U2782 ( .IN1(n2556), .IN2(n2460), .IN3(n2558), .IN4(reg2[25]), .IN5(
        n2459), .Q(n964) );
  NAND2X0 U2783 ( .IN1(n2529), .IN2(n2461), .QN(n2473) );
  NAND2X0 U2784 ( .IN1(n2485), .IN2(n2475), .QN(n2472) );
  NAND2X0 U2785 ( .IN1(n2463), .IN2(n2462), .QN(n2466) );
  INVX0 U2786 ( .INP(n2465), .ZN(n2464) );
  INVX0 U2787 ( .INP(n2466), .ZN(n2468) );
  AO221X1 U2788 ( .IN1(n2465), .IN2(n2466), .IN3(n2464), .IN4(n2468), .IN5(
        n2514), .Q(n2471) );
  AO221X1 U2789 ( .IN1(n2469), .IN2(n2468), .IN3(n2467), .IN4(n2466), .IN5(
        n2516), .Q(n2470) );
  NAND4X0 U2790 ( .IN1(n2473), .IN2(n2472), .IN3(n2471), .IN4(n2470), .QN(
        n2633) );
  MUX21X1 U2791 ( .IN1(n2476), .IN2(n2475), .S(n2474), .Q(n2631) );
  INVX0 U2792 ( .INP(n2631), .ZN(n2477) );
  AO22X1 U2793 ( .IN1(n2478), .IN2(n2539), .IN3(n2541), .IN4(n2477), .Q(n2479)
         );
  AO221X1 U2794 ( .IN1(n2556), .IN2(n2633), .IN3(n2558), .IN4(reg2[26]), .IN5(
        n2479), .Q(n963) );
  AO22X1 U2795 ( .IN1(n2481), .IN2(n2539), .IN3(n2541), .IN4(n2480), .Q(n2482)
         );
  AO221X1 U2796 ( .IN1(n2556), .IN2(n2483), .IN3(n2558), .IN4(reg2[27]), .IN5(
        n2482), .Q(n962) );
  NAND2X0 U2797 ( .IN1(n2529), .IN2(n2484), .QN(n2499) );
  NAND2X0 U2798 ( .IN1(n2485), .IN2(n2535), .QN(n2498) );
  OA21X1 U2799 ( .IN1(n2488), .IN2(n2487), .IN3(n2486), .Q(n2509) );
  NAND2X0 U2800 ( .IN1(n2508), .IN2(n2489), .QN(n2493) );
  INVX0 U2801 ( .INP(n2509), .ZN(n2490) );
  INVX0 U2802 ( .INP(n2493), .ZN(n2494) );
  AO221X1 U2803 ( .IN1(n2509), .IN2(n2493), .IN3(n2490), .IN4(n2494), .IN5(
        n2514), .Q(n2497) );
  AO222X1 U2804 ( .IN1(n2492), .IN2(n2688), .IN3(n2492), .IN4(n2491), .IN5(
        n2688), .IN6(n2491), .Q(n2506) );
  INVX0 U2805 ( .INP(n2506), .ZN(n2495) );
  AO221X1 U2806 ( .IN1(n2495), .IN2(n2494), .IN3(n2506), .IN4(n2493), .IN5(
        n2516), .Q(n2496) );
  NAND4X0 U2807 ( .IN1(n2499), .IN2(n2498), .IN3(n2497), .IN4(n2496), .QN(
        n2638) );
  MUX21X1 U2808 ( .IN1(n2500), .IN2(n2535), .S(n2534), .Q(n2636) );
  INVX0 U2809 ( .INP(n2636), .ZN(n2501) );
  AO22X1 U2810 ( .IN1(n2502), .IN2(n2539), .IN3(n2541), .IN4(n2501), .Q(n2503)
         );
  AO221X1 U2811 ( .IN1(n2556), .IN2(n2638), .IN3(n2558), .IN4(reg2[28]), .IN5(
        n2503), .Q(n961) );
  NAND2X0 U2812 ( .IN1(n2505), .IN2(n2504), .QN(n2511) );
  AO222X1 U2813 ( .IN1(n2535), .IN2(n2689), .IN3(n2535), .IN4(n2506), .IN5(
        n2689), .IN6(n2506), .Q(n2507) );
  XNOR2X1 U2814 ( .IN1(n2511), .IN2(n2507), .Q(n2515) );
  OA21X1 U2815 ( .IN1(n2510), .IN2(n2509), .IN3(n2508), .Q(n2512) );
  XNOR2X1 U2816 ( .IN1(n2512), .IN2(n2511), .Q(n2513) );
  OA22X1 U2817 ( .IN1(n2516), .IN2(n2515), .IN3(n2514), .IN4(n2513), .Q(n2533)
         );
  NAND2X0 U2818 ( .IN1(n2518), .IN2(n2517), .QN(n2526) );
  NOR2X0 U2819 ( .IN1(n2518), .IN2(n2517), .QN(n2524) );
  NOR2X0 U2820 ( .IN1(n2528), .IN2(n2519), .QN(n2522) );
  NAND2X0 U2821 ( .IN1(n2520), .IN2(B), .QN(n2521) );
  NAND2X0 U2822 ( .IN1(n2522), .IN2(n2521), .QN(n2523) );
  NOR2X0 U2823 ( .IN1(n2524), .IN2(n2523), .QN(n2552) );
  NAND3X0 U2824 ( .IN1(n2526), .IN2(n2525), .IN3(n2552), .QN(n2532) );
  OR2X1 U2825 ( .IN1(n2527), .IN2(n2536), .Q(n2531) );
  NAND3X0 U2826 ( .IN1(n2529), .IN2(n2528), .IN3(n2689), .QN(n2530) );
  NAND4X0 U2827 ( .IN1(n2533), .IN2(n2532), .IN3(n2531), .IN4(n2530), .QN(
        n2566) );
  NOR2X0 U2828 ( .IN1(n2535), .IN2(n2534), .QN(n2537) );
  NAND2X0 U2829 ( .IN1(n2537), .IN2(n2536), .QN(n2543) );
  OA21X1 U2830 ( .IN1(n2537), .IN2(n2536), .IN3(n2543), .Q(n2567) );
  INVX0 U2831 ( .INP(n2538), .ZN(n2540) );
  AO22X1 U2832 ( .IN1(n2567), .IN2(n2541), .IN3(n2540), .IN4(n2539), .Q(n2542)
         );
  AO221X1 U2833 ( .IN1(n2556), .IN2(n2566), .IN3(n2558), .IN4(reg2[29]), .IN5(
        n2542), .Q(n960) );
  INVX0 U2834 ( .INP(n2543), .ZN(n2546) );
  OA221X1 U2835 ( .IN1(n2546), .IN2(n2547), .IN3(n2543), .IN4(n2544), .IN5(
        n2548), .Q(n2569) );
  AO22X1 U2836 ( .IN1(n2554), .IN2(n2544), .IN3(n2552), .IN4(n2692), .Q(n2568)
         );
  AO21X1 U2837 ( .IN1(n2555), .IN2(n2569), .IN3(n2568), .Q(n2545) );
  OA222X1 U2838 ( .IN1(n2558), .IN2(n2570), .IN3(n2558), .IN4(n2545), .IN5(
        reg2[30]), .IN6(n2556), .Q(n959) );
  NAND2X0 U2839 ( .IN1(n2547), .IN2(n2546), .QN(n2549) );
  INVX0 U2840 ( .INP(n2549), .ZN(n2551) );
  INVX0 U2841 ( .INP(n2550), .ZN(n2553) );
  OA221X1 U2842 ( .IN1(n2551), .IN2(n2550), .IN3(n2549), .IN4(n2553), .IN5(
        n2548), .Q(n2572) );
  AO22X1 U2843 ( .IN1(n2554), .IN2(n2553), .IN3(n2552), .IN4(n2692), .Q(n2571)
         );
  AO21X1 U2844 ( .IN1(n2555), .IN2(n2572), .IN3(n2571), .Q(n2557) );
  OA222X1 U2845 ( .IN1(n2558), .IN2(n2570), .IN3(n2558), .IN4(n2557), .IN5(
        reg2[31]), .IN6(n2556), .Q(n958) );
  NOR2X0 U2846 ( .IN1(n2563), .IN2(n2619), .QN(n2559) );
  AO221X1 U2847 ( .IN1(n2565), .IN2(n2621), .IN3(n2573), .IN4(reg1[20]), .IN5(
        n2559), .Q(n937) );
  NOR2X0 U2848 ( .IN1(n2563), .IN2(n2623), .QN(n2560) );
  AO221X1 U2849 ( .IN1(n2565), .IN2(n2625), .IN3(n2573), .IN4(reg1[22]), .IN5(
        n2560), .Q(n935) );
  NOR2X0 U2850 ( .IN1(n2563), .IN2(n2627), .QN(n2561) );
  AO221X1 U2851 ( .IN1(n2565), .IN2(n2629), .IN3(n2573), .IN4(reg1[24]), .IN5(
        n2561), .Q(n933) );
  NOR2X0 U2852 ( .IN1(n2563), .IN2(n2631), .QN(n2562) );
  AO221X1 U2853 ( .IN1(n2565), .IN2(n2633), .IN3(n2573), .IN4(reg1[26]), .IN5(
        n2562), .Q(n931) );
  NOR2X0 U2854 ( .IN1(n2636), .IN2(n2563), .QN(n2564) );
  AO221X1 U2855 ( .IN1(n2565), .IN2(n2638), .IN3(n2573), .IN4(reg1[28]), .IN5(
        n2564), .Q(n929) );
  AO21X1 U2856 ( .IN1(n2567), .IN2(n2578), .IN3(n2566), .Q(n2640) );
  MUX21X1 U2857 ( .IN1(n2640), .IN2(reg1[29]), .S(n2573), .Q(n928) );
  OA21X1 U2858 ( .IN1(n2569), .IN2(n2568), .IN3(n2570), .Q(n2641) );
  MUX21X1 U2859 ( .IN1(n2641), .IN2(reg1[30]), .S(n2573), .Q(n927) );
  OA21X1 U2860 ( .IN1(n2572), .IN2(n2571), .IN3(n2570), .Q(n2643) );
  MUX21X1 U2861 ( .IN1(n2643), .IN2(reg1[31]), .S(n2573), .Q(n926) );
  NAND3X0 U2862 ( .IN1(n2574), .IN2(n2700), .IN3(n2709), .QN(n2577) );
  INVX0 U2863 ( .INP(n2575), .ZN(n2695) );
  AOI221X1 U2864 ( .IN1(n2577), .IN2(n2697), .IN3(n2577), .IN4(n2695), .IN5(
        n2576), .QN(n2639) );
  INVX0 U2865 ( .INP(n2639), .ZN(n2642) );
  NAND2X0 U2866 ( .IN1(n2578), .IN2(n2639), .QN(n2635) );
  NOR2X0 U2867 ( .IN1(n2579), .IN2(n2635), .QN(n2580) );
  AO221X1 U2868 ( .IN1(n2639), .IN2(n2581), .IN3(n2642), .IN4(reg0[0]), .IN5(
        n2580), .Q(n925) );
  MUX21X1 U2869 ( .IN1(n2582), .IN2(reg0[1]), .S(n2642), .Q(n924) );
  NOR2X0 U2870 ( .IN1(n2635), .IN2(n2583), .QN(n2584) );
  AO221X1 U2871 ( .IN1(n2639), .IN2(n2585), .IN3(n2642), .IN4(reg0[2]), .IN5(
        n2584), .Q(n923) );
  MUX21X1 U2872 ( .IN1(n2586), .IN2(reg0[3]), .S(n2642), .Q(n922) );
  NOR2X0 U2873 ( .IN1(n2635), .IN2(n2587), .QN(n2588) );
  AO221X1 U2874 ( .IN1(n2639), .IN2(n2589), .IN3(n2642), .IN4(reg0[4]), .IN5(
        n2588), .Q(n921) );
  MUX21X1 U2875 ( .IN1(n2590), .IN2(reg0[5]), .S(n2642), .Q(n920) );
  NOR2X0 U2876 ( .IN1(n2635), .IN2(n2591), .QN(n2592) );
  AO221X1 U2877 ( .IN1(n2639), .IN2(n2593), .IN3(n2642), .IN4(reg0[6]), .IN5(
        n2592), .Q(n919) );
  MUX21X1 U2878 ( .IN1(n2594), .IN2(reg0[7]), .S(n2642), .Q(n918) );
  NOR2X0 U2879 ( .IN1(n2635), .IN2(n2595), .QN(n2596) );
  AO221X1 U2880 ( .IN1(n2639), .IN2(n2597), .IN3(n2642), .IN4(reg0[8]), .IN5(
        n2596), .Q(n917) );
  MUX21X1 U2881 ( .IN1(n2598), .IN2(reg0[9]), .S(n2642), .Q(n916) );
  NOR2X0 U2882 ( .IN1(n2635), .IN2(n2599), .QN(n2600) );
  AO221X1 U2883 ( .IN1(n2639), .IN2(n2601), .IN3(n2642), .IN4(reg0[10]), .IN5(
        n2600), .Q(n915) );
  MUX21X1 U2884 ( .IN1(n2602), .IN2(reg0[11]), .S(n2642), .Q(n914) );
  NOR2X0 U2885 ( .IN1(n2635), .IN2(n2603), .QN(n2604) );
  AO221X1 U2886 ( .IN1(n2639), .IN2(n2605), .IN3(n2642), .IN4(reg0[12]), .IN5(
        n2604), .Q(n913) );
  MUX21X1 U2887 ( .IN1(n2606), .IN2(reg0[13]), .S(n2642), .Q(n912) );
  NOR2X0 U2888 ( .IN1(n2635), .IN2(n2607), .QN(n2608) );
  AO221X1 U2889 ( .IN1(n2639), .IN2(n2609), .IN3(n2642), .IN4(reg0[14]), .IN5(
        n2608), .Q(n911) );
  MUX21X1 U2890 ( .IN1(n2610), .IN2(reg0[15]), .S(n2642), .Q(n910) );
  NOR2X0 U2891 ( .IN1(n2635), .IN2(n2611), .QN(n2612) );
  AO221X1 U2892 ( .IN1(n2639), .IN2(n2613), .IN3(n2642), .IN4(reg0[16]), .IN5(
        n2612), .Q(n909) );
  MUX21X1 U2893 ( .IN1(n2614), .IN2(reg0[17]), .S(n2642), .Q(n908) );
  NOR2X0 U2894 ( .IN1(n2635), .IN2(n2615), .QN(n2616) );
  AO221X1 U2895 ( .IN1(n2639), .IN2(n2617), .IN3(n2642), .IN4(reg0[18]), .IN5(
        n2616), .Q(n907) );
  MUX21X1 U2896 ( .IN1(n2618), .IN2(reg0[19]), .S(n2642), .Q(n906) );
  NOR2X0 U2897 ( .IN1(n2635), .IN2(n2619), .QN(n2620) );
  AO221X1 U2898 ( .IN1(n2639), .IN2(n2621), .IN3(n2642), .IN4(reg0[20]), .IN5(
        n2620), .Q(n905) );
  MUX21X1 U2899 ( .IN1(n2622), .IN2(reg0[21]), .S(n2642), .Q(n904) );
  NOR2X0 U2900 ( .IN1(n2635), .IN2(n2623), .QN(n2624) );
  AO221X1 U2901 ( .IN1(n2639), .IN2(n2625), .IN3(n2642), .IN4(reg0[22]), .IN5(
        n2624), .Q(n903) );
  MUX21X1 U2902 ( .IN1(n2626), .IN2(reg0[23]), .S(n2642), .Q(n902) );
  NOR2X0 U2903 ( .IN1(n2635), .IN2(n2627), .QN(n2628) );
  AO221X1 U2904 ( .IN1(n2639), .IN2(n2629), .IN3(n2642), .IN4(reg0[24]), .IN5(
        n2628), .Q(n901) );
  MUX21X1 U2905 ( .IN1(n2630), .IN2(reg0[25]), .S(n2642), .Q(n900) );
  NOR2X0 U2906 ( .IN1(n2635), .IN2(n2631), .QN(n2632) );
  AO221X1 U2907 ( .IN1(n2639), .IN2(n2633), .IN3(n2642), .IN4(reg0[26]), .IN5(
        n2632), .Q(n899) );
  MUX21X1 U2908 ( .IN1(n2634), .IN2(reg0[27]), .S(n2642), .Q(n898) );
  NOR2X0 U2909 ( .IN1(n2636), .IN2(n2635), .QN(n2637) );
  AO221X1 U2910 ( .IN1(n2639), .IN2(n2638), .IN3(n2642), .IN4(reg0[28]), .IN5(
        n2637), .Q(n897) );
  MUX21X1 U2911 ( .IN1(reg0[29]), .IN2(n2640), .S(n2639), .Q(n896) );
  MUX21X1 U2912 ( .IN1(n2641), .IN2(reg0[30]), .S(n2642), .Q(n895) );
  MUX21X1 U2913 ( .IN1(n2643), .IN2(reg0[31]), .S(n2642), .Q(n894) );
  AO222X1 U2914 ( .IN1(n2703), .IN2(datai[20]), .IN3(IR[20]), .IN4(n2656), 
        .IN5(n2658), .IN6(n2644), .Q(n873) );
  AO222X1 U2915 ( .IN1(n2703), .IN2(datai[21]), .IN3(IR[21]), .IN4(n2656), 
        .IN5(n2658), .IN6(n2645), .Q(n872) );
  AO222X1 U2916 ( .IN1(n2703), .IN2(datai[22]), .IN3(IR[22]), .IN4(n2656), 
        .IN5(n2658), .IN6(n2646), .Q(n871) );
  AO222X1 U2917 ( .IN1(n2703), .IN2(datai[23]), .IN3(IR[23]), .IN4(n2656), 
        .IN5(n2658), .IN6(n2647), .Q(n870) );
  AO222X1 U2918 ( .IN1(n2703), .IN2(datai[24]), .IN3(IR[24]), .IN4(n2656), 
        .IN5(n2658), .IN6(n2648), .Q(n869) );
  AO222X1 U2919 ( .IN1(n2703), .IN2(datai[25]), .IN3(IR[25]), .IN4(n2656), 
        .IN5(n2658), .IN6(n2649), .Q(n868) );
  AO222X1 U2920 ( .IN1(n2703), .IN2(datai[26]), .IN3(IR[26]), .IN4(n2656), 
        .IN5(n2658), .IN6(n2650), .Q(n867) );
  INVX0 U2921 ( .INP(n2651), .ZN(n2652) );
  AO222X1 U2922 ( .IN1(n2703), .IN2(datai[27]), .IN3(IR[27]), .IN4(n2656), 
        .IN5(n2658), .IN6(n2652), .Q(n866) );
  AO222X1 U2923 ( .IN1(n2703), .IN2(datai[28]), .IN3(IR[28]), .IN4(n2656), 
        .IN5(n2658), .IN6(n2653), .Q(n865) );
  AO222X1 U2924 ( .IN1(n2703), .IN2(datai[29]), .IN3(IR[29]), .IN4(n2656), 
        .IN5(n2658), .IN6(n2654), .Q(n864) );
  AO222X1 U2925 ( .IN1(n2703), .IN2(datai[30]), .IN3(IR[30]), .IN4(n2656), 
        .IN5(n2658), .IN6(n2655), .Q(n863) );
  AO22X1 U2926 ( .IN1(n2658), .IN2(n2657), .IN3(datai[31]), .IN4(n2703), .Q(
        n862) );
  INVX0 U2927 ( .INP(n2659), .ZN(n2682) );
  MUX21X1 U2928 ( .IN1(datao[0]), .IN2(n2660), .S(n2682), .Q(n861) );
  MUX21X1 U2929 ( .IN1(datao[1]), .IN2(n2661), .S(n2682), .Q(n860) );
  MUX21X1 U2930 ( .IN1(datao[2]), .IN2(n2662), .S(n2682), .Q(n859) );
  MUX21X1 U2931 ( .IN1(datao[3]), .IN2(n2663), .S(n2682), .Q(n858) );
  MUX21X1 U2932 ( .IN1(datao[4]), .IN2(n2664), .S(n2682), .Q(n857) );
  MUX21X1 U2933 ( .IN1(datao[5]), .IN2(n2665), .S(n2682), .Q(n856) );
  MUX21X1 U2934 ( .IN1(datao[6]), .IN2(n2666), .S(n2682), .Q(n855) );
  MUX21X1 U2935 ( .IN1(datao[7]), .IN2(n2667), .S(n2682), .Q(n854) );
  MUX21X1 U2936 ( .IN1(datao[8]), .IN2(n2668), .S(n2682), .Q(n853) );
  MUX21X1 U2937 ( .IN1(datao[9]), .IN2(n2669), .S(n2682), .Q(n852) );
  MUX21X1 U2938 ( .IN1(datao[10]), .IN2(n2670), .S(n2682), .Q(n851) );
  MUX21X1 U2939 ( .IN1(datao[11]), .IN2(n2671), .S(n2682), .Q(n850) );
  MUX21X1 U2940 ( .IN1(datao[12]), .IN2(n2672), .S(n2736), .Q(n849) );
  MUX21X1 U2941 ( .IN1(datao[13]), .IN2(n2673), .S(n2736), .Q(n848) );
  MUX21X1 U2942 ( .IN1(datao[14]), .IN2(n2674), .S(n2736), .Q(n847) );
  MUX21X1 U2943 ( .IN1(datao[15]), .IN2(n2675), .S(n2736), .Q(n846) );
  MUX21X1 U2944 ( .IN1(datao[16]), .IN2(n2676), .S(n2682), .Q(n845) );
  MUX21X1 U2945 ( .IN1(datao[17]), .IN2(n2677), .S(n2736), .Q(n844) );
  MUX21X1 U2946 ( .IN1(datao[18]), .IN2(n2678), .S(n2682), .Q(n843) );
  MUX21X1 U2947 ( .IN1(datao[19]), .IN2(n2679), .S(n2736), .Q(n842) );
  MUX21X1 U2948 ( .IN1(datao[20]), .IN2(n2680), .S(n2682), .Q(n841) );
  MUX21X1 U2949 ( .IN1(datao[21]), .IN2(n2681), .S(n2736), .Q(n840) );
  MUX21X1 U2950 ( .IN1(datao[22]), .IN2(n2683), .S(n2682), .Q(n839) );
  MUX21X1 U2951 ( .IN1(datao[23]), .IN2(n2684), .S(n2736), .Q(n838) );
  MUX21X1 U2952 ( .IN1(datao[24]), .IN2(n2685), .S(n2736), .Q(n837) );
  MUX21X1 U2953 ( .IN1(datao[25]), .IN2(n2686), .S(n2736), .Q(n836) );
  MUX21X1 U2954 ( .IN1(datao[26]), .IN2(n2687), .S(n2736), .Q(n835) );
  MUX21X1 U2955 ( .IN1(datao[27]), .IN2(n2688), .S(n2736), .Q(n834) );
  MUX21X1 U2956 ( .IN1(datao[28]), .IN2(n2689), .S(n2736), .Q(n833) );
  MUX21X1 U2957 ( .IN1(datao[29]), .IN2(n2690), .S(n2736), .Q(n832) );
  MUX21X1 U2958 ( .IN1(datao[30]), .IN2(n2691), .S(n2736), .Q(n831) );
  MUX21X1 U2959 ( .IN1(datao[31]), .IN2(n2692), .S(n2736), .Q(n830) );
  NAND3X0 U2960 ( .IN1(n2694), .IN2(state), .IN3(n2693), .QN(n2696) );
  MUX21X1 U2961 ( .IN1(n2695), .IN2(d[0]), .S(n2696), .Q(n828) );
  MUX21X1 U2962 ( .IN1(n2697), .IN2(d[1]), .S(n2696), .Q(n827) );
endmodule

