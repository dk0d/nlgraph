
module divider ( in, out, N, reset );
  input [5:0] N;
  input in, reset;
  output out;
  wire   \even_0/out_counter , \odd_0/rst_pulse , \odd_0/out_counter ,
         \odd_0/out_counter2 , n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303;
  wire   [5:0] \even_0/counter ;
  wire   [5:0] \odd_0/old_N ;
  wire   [5:0] \odd_0/initial_begin ;
  wire   [5:0] \odd_0/counter2 ;
  wire   [5:0] \odd_0/counter ;

  DFFARX1 \even_0/counter_reg[5]  ( .D(n117), .CLK(in), .RSTB(n111), .Q(
        \even_0/counter [5]) );
  DFFARX1 \even_0/counter_reg[1]  ( .D(n116), .CLK(in), .RSTB(n111), .Q(
        \even_0/counter [1]), .QN(n298) );
  DFFARX1 \even_0/counter_reg[2]  ( .D(n115), .CLK(in), .RSTB(n111), .Q(
        \even_0/counter [2]) );
  DFFARX1 \even_0/counter_reg[3]  ( .D(n114), .CLK(in), .RSTB(n111), .Q(
        \even_0/counter [3]) );
  DFFARX1 \even_0/counter_reg[4]  ( .D(n113), .CLK(in), .RSTB(n111), .Q(
        \even_0/counter [4]), .QN(n296) );
  DFFASX1 \even_0/counter_reg[0]  ( .D(n112), .CLK(in), .SETB(n111), .Q(
        \even_0/counter [0]), .QN(n295) );
  DFFASX1 \even_0/out_counter_reg  ( .D(n139), .CLK(in), .SETB(n111), .Q(
        \even_0/out_counter ) );
  DFFX1 \odd_0/old_N_reg[0]  ( .D(N[0]), .CLK(in), .Q(\odd_0/old_N [0]) );
  DFFX1 \odd_0/old_N_reg[1]  ( .D(N[1]), .CLK(in), .Q(\odd_0/old_N [1]) );
  DFFX1 \odd_0/old_N_reg[2]  ( .D(N[2]), .CLK(in), .Q(\odd_0/old_N [2]) );
  DFFX1 \odd_0/old_N_reg[3]  ( .D(N[3]), .CLK(in), .Q(\odd_0/old_N [3]) );
  DFFX1 \odd_0/old_N_reg[4]  ( .D(N[4]), .CLK(in), .Q(\odd_0/old_N [4]) );
  DFFX1 \odd_0/old_N_reg[5]  ( .D(N[5]), .CLK(in), .Q(\odd_0/old_N [5]) );
  DFFX1 \odd_0/counter_reg[5]  ( .D(n124), .CLK(in), .Q(\odd_0/counter [5]), 
        .QN(n301) );
  DFFX1 \odd_0/counter_reg[3]  ( .D(n118), .CLK(in), .QN(n299) );
  DFFX1 \odd_0/out_counter_reg  ( .D(n122), .CLK(in), .Q(\odd_0/out_counter ), 
        .QN(n291) );
  DFFX1 \odd_0/counter_reg[0]  ( .D(n121), .CLK(in), .Q(\odd_0/counter [0]), 
        .QN(n303) );
  DFFX1 \odd_0/counter_reg[2]  ( .D(n119), .CLK(in), .Q(\odd_0/counter [2]) );
  DFFX1 \odd_0/counter_reg[1]  ( .D(n120), .CLK(in), .Q(\odd_0/counter [1]) );
  DFFX1 \odd_0/counter_reg[4]  ( .D(n123), .CLK(in), .Q(\odd_0/counter [4]) );
  DFFARX1 \odd_0/rst_pulse_reg  ( .D(n138), .CLK(in), .RSTB(n111), .Q(
        \odd_0/rst_pulse ) );
  DFFNX1 \odd_0/initial_begin_reg[5]  ( .D(n137), .CLK(in), .Q(
        \odd_0/initial_begin [5]) );
  DFFNX1 \odd_0/initial_begin_reg[1]  ( .D(n133), .CLK(in), .Q(
        \odd_0/initial_begin [1]) );
  DFFNX1 \odd_0/initial_begin_reg[4]  ( .D(n135), .CLK(in), .Q(
        \odd_0/initial_begin [4]), .QN(n293) );
  DFFNX1 \odd_0/initial_begin_reg[2]  ( .D(n132), .CLK(in), .Q(
        \odd_0/initial_begin [2]), .QN(n297) );
  DFFNX1 \odd_0/initial_begin_reg[3]  ( .D(n131), .CLK(in), .Q(
        \odd_0/initial_begin [3]) );
  DFFNX1 \odd_0/initial_begin_reg[0]  ( .D(n134), .CLK(in), .Q(
        \odd_0/initial_begin [0]), .QN(n302) );
  DFFNX1 \odd_0/counter2_reg[4]  ( .D(n125), .CLK(in), .Q(\odd_0/counter2 [4])
         );
  DFFNX1 \odd_0/counter2_reg[0]  ( .D(n129), .CLK(in), .Q(\odd_0/counter2 [0]), 
        .QN(n292) );
  DFFNX1 \odd_0/out_counter2_reg  ( .D(n136), .CLK(in), .Q(
        \odd_0/out_counter2 ), .QN(n294) );
  DFFNX1 \odd_0/counter2_reg[5]  ( .D(n130), .CLK(in), .Q(\odd_0/counter2 [5])
         );
  DFFNX1 \odd_0/counter2_reg[1]  ( .D(n128), .CLK(in), .Q(\odd_0/counter2 [1])
         );
  DFFNX1 \odd_0/counter2_reg[2]  ( .D(n127), .CLK(in), .Q(\odd_0/counter2 [2]), 
        .QN(n300) );
  DFFNX1 \odd_0/counter2_reg[3]  ( .D(n126), .CLK(in), .Q(\odd_0/counter2 [3])
         );
  INVX0 U141 ( .INP(reset), .ZN(n111) );
  INVX0 U142 ( .INP(N[1]), .ZN(n214) );
  OR3X1 U143 ( .IN1(\even_0/counter [1]), .IN2(\even_0/counter [3]), .IN3(
        \even_0/counter [2]), .Q(n143) );
  OR4X1 U144 ( .IN1(\even_0/counter [5]), .IN2(\even_0/counter [4]), .IN3(n143), .IN4(n295), .Q(n145) );
  NOR2X0 U145 ( .IN1(n214), .IN2(n145), .QN(n140) );
  INVX0 U146 ( .INP(N[0]), .ZN(n272) );
  NAND2X0 U147 ( .IN1(n272), .IN2(n295), .QN(n284) );
  INVX0 U148 ( .INP(n284), .ZN(n285) );
  NOR2X0 U149 ( .IN1(n140), .IN2(n285), .QN(n142) );
  NAND2X0 U150 ( .IN1(\even_0/counter [0]), .IN2(N[0]), .QN(n141) );
  NAND2X0 U151 ( .IN1(n142), .IN2(n141), .QN(n112) );
  NOR2X0 U152 ( .IN1(n284), .IN2(n143), .QN(n289) );
  NAND2X0 U153 ( .IN1(n285), .IN2(n298), .QN(n287) );
  OA21X1 U154 ( .IN1(\even_0/counter [2]), .IN2(n287), .IN3(
        \even_0/counter [3]), .Q(n144) );
  NOR2X0 U155 ( .IN1(n289), .IN2(n144), .QN(n147) );
  NOR2X0 U156 ( .IN1(N[0]), .IN2(n145), .QN(n288) );
  NAND2X0 U157 ( .IN1(n288), .IN2(N[4]), .QN(n146) );
  NAND2X0 U158 ( .IN1(n147), .IN2(n146), .QN(n114) );
  NOR2X0 U159 ( .IN1(reset), .IN2(\odd_0/rst_pulse ), .QN(n255) );
  INVX0 U160 ( .INP(N[5]), .ZN(n201) );
  INVX0 U161 ( .INP(N[4]), .ZN(n256) );
  INVX0 U162 ( .INP(N[3]), .ZN(n279) );
  NAND4X0 U163 ( .IN1(n201), .IN2(n214), .IN3(n256), .IN4(n279), .QN(n200) );
  OR2X1 U164 ( .IN1(n200), .IN2(N[2]), .Q(n190) );
  NAND2X0 U165 ( .IN1(N[0]), .IN2(n190), .QN(n236) );
  INVX0 U166 ( .INP(n236), .ZN(n264) );
  NOR4X0 U167 ( .IN1(\odd_0/counter [5]), .IN2(\odd_0/counter [4]), .IN3(
        \odd_0/counter [2]), .IN4(\odd_0/counter [1]), .QN(n148) );
  AND3X1 U168 ( .IN1(\odd_0/counter [0]), .IN2(n148), .IN3(n299), .Q(n262) );
  NAND2X0 U169 ( .IN1(n264), .IN2(n262), .QN(n149) );
  MUX21X1 U170 ( .IN1(\odd_0/out_counter ), .IN2(n291), .S(n149), .Q(n150) );
  NAND2X0 U171 ( .IN1(n255), .IN2(n150), .QN(n122) );
  OR4X1 U172 ( .IN1(\odd_0/initial_begin [4]), .IN2(\odd_0/initial_begin [5]), 
        .IN3(\odd_0/initial_begin [3]), .IN4(\odd_0/initial_begin [1]), .Q(
        n151) );
  NOR2X0 U173 ( .IN1(\odd_0/initial_begin [2]), .IN2(n151), .QN(n237) );
  NAND2X0 U174 ( .IN1(n255), .IN2(n237), .QN(n213) );
  NOR2X0 U175 ( .IN1(n236), .IN2(n213), .QN(n230) );
  INVX0 U176 ( .INP(n255), .ZN(n261) );
  NOR2X0 U177 ( .IN1(n261), .IN2(n264), .QN(n267) );
  INVX0 U178 ( .INP(n267), .ZN(n275) );
  INVX0 U179 ( .INP(n237), .ZN(n235) );
  NAND2X0 U180 ( .IN1(n255), .IN2(n235), .QN(n157) );
  NAND2X0 U181 ( .IN1(n275), .IN2(n157), .QN(n228) );
  AO221X1 U182 ( .IN1(n230), .IN2(\odd_0/counter2 [0]), .IN3(n230), .IN4(
        \odd_0/counter2 [1]), .IN5(n228), .Q(n247) );
  OA221X1 U183 ( .IN1(n247), .IN2(\odd_0/counter2 [2]), .IN3(n247), .IN4(n230), 
        .IN5(\odd_0/counter2 [3]), .Q(n152) );
  OR4X1 U184 ( .IN1(\odd_0/counter2 [0]), .IN2(\odd_0/counter2 [1]), .IN3(
        \odd_0/counter2 [3]), .IN4(\odd_0/counter2 [2]), .Q(n229) );
  INVX0 U185 ( .INP(n230), .ZN(n186) );
  NOR2X0 U186 ( .IN1(n229), .IN2(n186), .QN(n178) );
  NOR2X0 U187 ( .IN1(n152), .IN2(n178), .QN(n156) );
  OR3X1 U188 ( .IN1(\odd_0/counter2 [1]), .IN2(\odd_0/counter2 [3]), .IN3(
        \odd_0/counter2 [2]), .Q(n153) );
  NOR4X0 U189 ( .IN1(\odd_0/counter2 [4]), .IN2(\odd_0/counter2 [5]), .IN3(
        n153), .IN4(n292), .QN(n238) );
  NAND3X0 U190 ( .IN1(N[0]), .IN2(n238), .IN3(n237), .QN(n154) );
  NAND2X0 U191 ( .IN1(n154), .IN2(n255), .QN(n234) );
  NAND2X0 U192 ( .IN1(N[3]), .IN2(n234), .QN(n155) );
  NAND2X0 U193 ( .IN1(n156), .IN2(n155), .QN(n126) );
  NOR2X0 U194 ( .IN1(\odd_0/initial_begin [1]), .IN2(\odd_0/initial_begin [0]), 
        .QN(n223) );
  NOR2X0 U195 ( .IN1(n236), .IN2(n157), .QN(n216) );
  OA221X1 U196 ( .IN1(n223), .IN2(\odd_0/initial_begin [1]), .IN3(n223), .IN4(
        \odd_0/initial_begin [0]), .IN5(n216), .Q(n162) );
  NAND2X0 U197 ( .IN1(n272), .IN2(n214), .QN(n158) );
  NOR2X0 U198 ( .IN1(n158), .IN2(N[2]), .QN(n160) );
  NAND2X0 U199 ( .IN1(N[2]), .IN2(n158), .QN(n219) );
  NAND2X0 U200 ( .IN1(n261), .IN2(n219), .QN(n159) );
  NOR2X0 U201 ( .IN1(n160), .IN2(n159), .QN(n161) );
  NOR2X0 U202 ( .IN1(n162), .IN2(n161), .QN(n164) );
  NAND2X0 U203 ( .IN1(n267), .IN2(\odd_0/initial_begin [1]), .QN(n163) );
  NAND2X0 U204 ( .IN1(n164), .IN2(n163), .QN(n133) );
  NAND2X0 U205 ( .IN1(n223), .IN2(n297), .QN(n224) );
  NOR2X0 U206 ( .IN1(\odd_0/initial_begin [3]), .IN2(n224), .QN(n170) );
  NAND2X0 U207 ( .IN1(n170), .IN2(n293), .QN(n208) );
  OA21X1 U208 ( .IN1(n170), .IN2(n293), .IN3(n208), .Q(n165) );
  INVX0 U209 ( .INP(n216), .ZN(n222) );
  OA22X1 U210 ( .IN1(n165), .IN2(n222), .IN3(n293), .IN4(n275), .Q(n169) );
  NOR2X0 U211 ( .IN1(n279), .IN2(n219), .QN(n218) );
  NAND2X0 U212 ( .IN1(N[4]), .IN2(n218), .QN(n171) );
  NOR2X0 U213 ( .IN1(n201), .IN2(n171), .QN(n212) );
  NOR2X0 U214 ( .IN1(n212), .IN2(n255), .QN(n167) );
  NAND2X0 U215 ( .IN1(n201), .IN2(n171), .QN(n166) );
  NAND2X0 U216 ( .IN1(n167), .IN2(n166), .QN(n168) );
  NAND2X0 U217 ( .IN1(n169), .IN2(n168), .QN(n135) );
  OA221X1 U218 ( .IN1(n170), .IN2(\odd_0/initial_begin [3]), .IN3(n170), .IN4(
        n224), .IN5(n216), .Q(n175) );
  NOR2X0 U219 ( .IN1(n218), .IN2(N[4]), .QN(n173) );
  NAND2X0 U220 ( .IN1(n261), .IN2(n171), .QN(n172) );
  NOR2X0 U221 ( .IN1(n173), .IN2(n172), .QN(n174) );
  NOR2X0 U222 ( .IN1(n175), .IN2(n174), .QN(n177) );
  NAND2X0 U223 ( .IN1(n267), .IN2(\odd_0/initial_begin [3]), .QN(n176) );
  NAND2X0 U224 ( .IN1(n177), .IN2(n176), .QN(n131) );
  INVX0 U225 ( .INP(n178), .ZN(n179) );
  NOR2X0 U226 ( .IN1(\odd_0/counter2 [4]), .IN2(n179), .QN(n232) );
  INVX0 U227 ( .INP(n234), .ZN(n244) );
  NOR2X0 U228 ( .IN1(n244), .IN2(n256), .QN(n180) );
  NOR2X0 U229 ( .IN1(n232), .IN2(n180), .QN(n183) );
  AO21X1 U230 ( .IN1(n230), .IN2(n229), .IN3(n228), .Q(n181) );
  NAND2X0 U231 ( .IN1(\odd_0/counter2 [4]), .IN2(n181), .QN(n182) );
  NAND2X0 U232 ( .IN1(n183), .IN2(n182), .QN(n125) );
  NAND3X0 U233 ( .IN1(n264), .IN2(n237), .IN3(n238), .QN(n184) );
  MUX21X1 U234 ( .IN1(\odd_0/out_counter2 ), .IN2(n294), .S(n184), .Q(n185) );
  NAND2X0 U235 ( .IN1(n255), .IN2(n185), .QN(n136) );
  NOR3X0 U236 ( .IN1(\odd_0/counter2 [0]), .IN2(\odd_0/counter2 [1]), .IN3(
        n186), .QN(n246) );
  OA221X1 U237 ( .IN1(n228), .IN2(\odd_0/counter2 [0]), .IN3(n228), .IN4(n230), 
        .IN5(\odd_0/counter2 [1]), .Q(n187) );
  NOR2X0 U238 ( .IN1(n246), .IN2(n187), .QN(n189) );
  NAND2X0 U239 ( .IN1(N[1]), .IN2(n234), .QN(n188) );
  NAND2X0 U240 ( .IN1(n189), .IN2(n188), .QN(n128) );
  MUX21X1 U241 ( .IN1(n294), .IN2(\odd_0/out_counter2 ), .S(n291), .Q(n192) );
  MUX21X1 U242 ( .IN1(in), .IN2(\even_0/out_counter ), .S(n190), .Q(n191) );
  AO22X1 U243 ( .IN1(n192), .IN2(n264), .IN3(n191), .IN4(n272), .Q(out) );
  INVX0 U244 ( .INP(n288), .ZN(n193) );
  MUX21X1 U245 ( .IN1(n288), .IN2(n193), .S(\even_0/out_counter ), .Q(n139) );
  OA22X1 U246 ( .IN1(\odd_0/old_N [3]), .IN2(n279), .IN3(\odd_0/old_N [1]), 
        .IN4(n214), .Q(n199) );
  NAND2X0 U247 ( .IN1(n256), .IN2(\odd_0/old_N [4]), .QN(n195) );
  NOR4X0 U248 ( .IN1(N[2]), .IN2(N[5]), .IN3(N[1]), .IN4(N[3]), .QN(n257) );
  INVX0 U249 ( .INP(N[2]), .ZN(n243) );
  OA22X1 U250 ( .IN1(\odd_0/old_N [2]), .IN2(n243), .IN3(\odd_0/old_N [5]), 
        .IN4(n201), .Q(n194) );
  OA221X1 U251 ( .IN1(n195), .IN2(n257), .IN3(n256), .IN4(\odd_0/old_N [4]), 
        .IN5(n194), .Q(n198) );
  NAND4X0 U252 ( .IN1(n243), .IN2(n201), .IN3(n256), .IN4(n279), .QN(n196) );
  NAND3X0 U253 ( .IN1(\odd_0/old_N [1]), .IN2(n214), .IN3(n196), .QN(n197) );
  AND3X1 U254 ( .IN1(n199), .IN2(n198), .IN3(n197), .Q(n205) );
  NAND3X0 U255 ( .IN1(\odd_0/old_N [2]), .IN2(n243), .IN3(n200), .QN(n204) );
  NAND4X0 U256 ( .IN1(n243), .IN2(n214), .IN3(n256), .IN4(n279), .QN(n250) );
  NAND3X0 U257 ( .IN1(\odd_0/old_N [5]), .IN2(n201), .IN3(n250), .QN(n203) );
  NAND4X0 U258 ( .IN1(n243), .IN2(n201), .IN3(n214), .IN4(n256), .QN(n271) );
  NAND3X0 U259 ( .IN1(\odd_0/old_N [3]), .IN2(n279), .IN3(n271), .QN(n202) );
  NAND4X0 U260 ( .IN1(n205), .IN2(n204), .IN3(n203), .IN4(n202), .QN(n206) );
  AOI22X1 U261 ( .IN1(N[0]), .IN2(n206), .IN3(\odd_0/rst_pulse ), .IN4(n236), 
        .QN(n207) );
  OAI21X1 U262 ( .IN1(\odd_0/old_N [0]), .IN2(n236), .IN3(n207), .QN(n138) );
  NOR2X0 U263 ( .IN1(n208), .IN2(n236), .QN(n210) );
  NAND2X0 U264 ( .IN1(n255), .IN2(\odd_0/initial_begin [5]), .QN(n209) );
  NOR2X0 U265 ( .IN1(n210), .IN2(n209), .QN(n211) );
  AO21X1 U266 ( .IN1(n212), .IN2(n261), .IN3(n211), .Q(n137) );
  NAND2X0 U267 ( .IN1(n213), .IN2(n275), .QN(n217) );
  OA221X1 U268 ( .IN1(N[1]), .IN2(n272), .IN3(n214), .IN4(N[0]), .IN5(n261), 
        .Q(n215) );
  AO221X1 U269 ( .IN1(\odd_0/initial_begin [0]), .IN2(n217), .IN3(n302), .IN4(
        n216), .IN5(n215), .Q(n134) );
  NAND2X0 U270 ( .IN1(\odd_0/initial_begin [2]), .IN2(n267), .QN(n227) );
  NOR2X0 U271 ( .IN1(n218), .IN2(n255), .QN(n221) );
  NAND2X0 U272 ( .IN1(n279), .IN2(n219), .QN(n220) );
  NAND2X0 U273 ( .IN1(n221), .IN2(n220), .QN(n226) );
  AO221X1 U274 ( .IN1(n224), .IN2(n223), .IN3(n224), .IN4(n297), .IN5(n222), 
        .Q(n225) );
  NAND3X0 U275 ( .IN1(n227), .IN2(n226), .IN3(n225), .QN(n132) );
  AO221X1 U276 ( .IN1(n230), .IN2(\odd_0/counter2 [4]), .IN3(n230), .IN4(n229), 
        .IN5(n228), .Q(n231) );
  MUX21X1 U277 ( .IN1(n232), .IN2(n231), .S(\odd_0/counter2 [5]), .Q(n233) );
  AO21X1 U278 ( .IN1(N[5]), .IN2(n234), .IN3(n233), .Q(n130) );
  NOR2X0 U279 ( .IN1(n236), .IN2(n235), .QN(n242) );
  NOR2X0 U280 ( .IN1(n237), .IN2(n292), .QN(n239) );
  NOR3X0 U281 ( .IN1(n239), .IN2(n238), .IN3(n261), .QN(n240) );
  NOR2X0 U282 ( .IN1(n240), .IN2(n272), .QN(n241) );
  AO221X1 U283 ( .IN1(\odd_0/counter2 [0]), .IN2(n267), .IN3(n292), .IN4(n242), 
        .IN5(n241), .Q(n129) );
  NOR2X0 U284 ( .IN1(n244), .IN2(n243), .QN(n245) );
  AO221X1 U285 ( .IN1(\odd_0/counter2 [2]), .IN2(n247), .IN3(n300), .IN4(n246), 
        .IN5(n245), .Q(n127) );
  NAND2X0 U286 ( .IN1(N[0]), .IN2(n262), .QN(n248) );
  NAND2X0 U287 ( .IN1(n255), .IN2(n248), .QN(n277) );
  NOR2X0 U288 ( .IN1(\odd_0/counter [1]), .IN2(\odd_0/counter [0]), .QN(n265)
         );
  INVX0 U289 ( .INP(n265), .ZN(n268) );
  NOR2X0 U290 ( .IN1(\odd_0/counter [2]), .IN2(n268), .QN(n276) );
  NAND2X0 U291 ( .IN1(n276), .IN2(n299), .QN(n281) );
  NOR2X0 U292 ( .IN1(\odd_0/counter [4]), .IN2(n281), .QN(n249) );
  MUX21X1 U293 ( .IN1(\odd_0/counter [5]), .IN2(n301), .S(n249), .Q(n253) );
  NOR2X0 U294 ( .IN1(n250), .IN2(N[5]), .QN(n252) );
  NAND2X0 U295 ( .IN1(N[0]), .IN2(n255), .QN(n251) );
  NOR2X0 U296 ( .IN1(n252), .IN2(n251), .QN(n269) );
  AO22X1 U297 ( .IN1(N[5]), .IN2(n277), .IN3(n253), .IN4(n269), .Q(n254) );
  AO21X1 U298 ( .IN1(n267), .IN2(\odd_0/counter [5]), .IN3(n254), .Q(n124) );
  NAND2X0 U299 ( .IN1(N[0]), .IN2(n255), .QN(n273) );
  OAI22X1 U300 ( .IN1(n257), .IN2(n273), .IN3(n272), .IN4(n256), .QN(n259) );
  XNOR2X1 U301 ( .IN1(\odd_0/counter [4]), .IN2(n281), .Q(n258) );
  AO22X1 U302 ( .IN1(\odd_0/counter [4]), .IN2(n267), .IN3(n259), .IN4(n258), 
        .Q(n260) );
  AO21X1 U303 ( .IN1(N[4]), .IN2(n277), .IN3(n260), .Q(n123) );
  OA21X1 U304 ( .IN1(n262), .IN2(n261), .IN3(N[0]), .Q(n263) );
  AO221X1 U305 ( .IN1(\odd_0/counter [0]), .IN2(n267), .IN3(n303), .IN4(n264), 
        .IN5(n263), .Q(n121) );
  AO21X1 U306 ( .IN1(\odd_0/counter [0]), .IN2(n269), .IN3(n267), .Q(n266) );
  AO222X1 U307 ( .IN1(n266), .IN2(\odd_0/counter [1]), .IN3(n269), .IN4(n265), 
        .IN5(n277), .IN6(N[1]), .Q(n120) );
  AO21X1 U308 ( .IN1(n268), .IN2(n269), .IN3(n267), .Q(n270) );
  AO222X1 U309 ( .IN1(n270), .IN2(\odd_0/counter [2]), .IN3(n269), .IN4(n276), 
        .IN5(n277), .IN6(N[2]), .Q(n119) );
  INVX0 U310 ( .INP(n271), .ZN(n274) );
  OA22X1 U311 ( .IN1(n274), .IN2(n273), .IN3(n272), .IN4(n279), .Q(n280) );
  OA21X1 U312 ( .IN1(n276), .IN2(n280), .IN3(n275), .Q(n282) );
  INVX0 U313 ( .INP(n277), .ZN(n278) );
  OAI222X1 U314 ( .IN1(n299), .IN2(n282), .IN3(n281), .IN4(n280), .IN5(n279), 
        .IN6(n278), .QN(n118) );
  NAND2X0 U315 ( .IN1(n289), .IN2(n296), .QN(n283) );
  XNOR2X1 U316 ( .IN1(\even_0/counter [5]), .IN2(n283), .Q(n117) );
  AO222X1 U317 ( .IN1(n285), .IN2(n298), .IN3(n284), .IN4(\even_0/counter [1]), 
        .IN5(N[2]), .IN6(n288), .Q(n116) );
  NOR2X0 U318 ( .IN1(n287), .IN2(\even_0/counter [2]), .QN(n286) );
  AO221X1 U319 ( .IN1(n288), .IN2(N[3]), .IN3(n287), .IN4(\even_0/counter [2]), 
        .IN5(n286), .Q(n115) );
  INVX0 U320 ( .INP(n289), .ZN(n290) );
  AO222X1 U321 ( .IN1(\even_0/counter [4]), .IN2(n290), .IN3(n296), .IN4(n289), 
        .IN5(N[5]), .IN6(n288), .Q(n113) );
endmodule

