
module top ( enable, degrees, data1, rst, actv, clock );
  input [31:0] degrees;
  output [63:0] data1;
  input [2:0] actv;
  input enable, rst, clock;
  wire   N324, N325, N326, N327, N328, N329, N330, N331, N332, N334, N356,
         N357, N386, N387, N388, N389, N390, N391, N392, N393, N394, N395,
         N396, N397, N398, N399, N400, N401, N402, N403, N404, N405, N406,
         N407, N408, N409, N410, N411, N412, N413, N414, N415, N416, N417,
         N418, N419, N420, N421, N422, N423, N424, N425, N426, N427, N428,
         N429, N430, N431, N432, N433, N434, N435, N436, N437, N438, N439,
         N440, N441, N442, N443, N444, N445, N446, N447, N448, N449, \a1/N491 ,
         \a1/N490 , \a1/N489 , \a1/N488 , \a1/N487 , \a1/N486 , \a1/N485 ,
         \a1/N484 , \a1/N483 , \a1/N482 , \a1/N481 , \a1/N480 , \a1/N479 ,
         \a1/N478 , \a1/N477 , \a1/N476 , \a1/N475 , \a1/N474 , \a1/N473 ,
         \a1/N472 , \a1/N471 , \a1/N470 , \a1/N469 , \a1/N468 , \a1/N467 ,
         \a1/N466 , \a1/N465 , \a1/N464 , \a1/N463 , \a1/N462 , \a1/N461 ,
         \a1/N460 , \a1/N459 , \a1/N458 , \a1/N457 , \a1/N456 , \a1/N455 ,
         \a1/N454 , \a1/N453 , \a1/N452 , \a1/N451 , \a1/N450 , \a1/N449 ,
         \a1/N448 , \a1/N447 , \a1/N446 , \a1/N445 , \a1/N444 , \a1/N443 ,
         \a1/N442 , \a1/N441 , \a1/N440 , \a1/N439 , \a1/N438 , \a1/N437 ,
         \a1/N436 , \a1/N435 , \a2/N491 , \a2/N490 , \a2/N489 , \a2/N488 ,
         \a2/N487 , \a2/N486 , \a2/N485 , \a2/N484 , \a2/N483 , \a2/N482 ,
         \a2/N481 , \a2/N480 , \a2/N479 , \a2/N478 , \a2/N477 , \a2/N476 ,
         \a2/N475 , \a2/N474 , \a2/N473 , \a2/N472 , \a2/N471 , \a2/N470 ,
         \a2/N469 , \a2/N468 , \a2/N467 , \a2/N466 , \a2/N465 , \a2/N464 ,
         \a2/N463 , \a2/N462 , \a2/N461 , \a2/N460 , \a2/N459 , \a2/N458 ,
         \a2/N457 , \a2/N456 , \a2/N455 , \a2/N454 , \a2/N453 , \a2/N452 ,
         \a2/N451 , \a2/N450 , \a2/N449 , \a2/N448 , \a2/N447 , \a2/N446 ,
         \a2/N445 , \a2/N444 , \a2/N443 , \a2/N442 , \a2/N441 , \a2/N440 ,
         \a2/N439 , \a2/N438 , \a2/N437 , \a2/N436 , \a2/N435 , \a3/N493 ,
         \a3/N492 , \a3/N491 , \a3/N490 , \a3/N489 , \a3/N488 , \a3/N487 ,
         \a3/N486 , \a3/N485 , \a3/N484 , \a3/N483 , \a3/N482 , \a3/N481 ,
         \a3/N480 , \a3/N479 , \a3/N478 , \a3/N477 , \a3/N476 , \a3/N475 ,
         \a3/N474 , \a3/N473 , \a3/N472 , \a3/N471 , \a3/N470 , \a3/N469 ,
         \a3/N468 , \a3/N467 , \a3/N466 , \a3/N465 , \a3/N464 , \a3/N463 ,
         \a3/N462 , \a3/N461 , \a3/N460 , \a3/N459 , \a3/N458 , \a3/N457 ,
         \a3/N456 , \a3/N455 , \a3/N454 , \a3/N453 , \a3/N452 , \a3/N451 ,
         \a3/N450 , \a3/N449 , \a3/N448 , \a3/N447 , \a3/N446 , \a3/N445 ,
         \a3/N444 , \a3/N443 , \a3/N442 , \a3/N441 , \a3/N440 , \a3/N439 ,
         \a3/N438 , \a3/N437 , \a3/N436 , \a4/N492 , \a4/N491 , \a4/N490 ,
         \a4/N489 , \a4/N488 , \a4/N487 , \a4/N486 , \a4/N485 , \a4/N484 ,
         \a4/N483 , \a4/N482 , \a4/N481 , \a4/N480 , \a4/N479 , \a4/N478 ,
         \a4/N477 , \a4/N476 , \a4/N475 , \a4/N474 , \a4/N473 , \a4/N472 ,
         \a4/N471 , \a4/N470 , \a4/N469 , \a4/N468 , \a4/N467 , \a4/N466 ,
         \a4/N465 , \a4/N464 , \a4/N463 , \a4/N462 , \a4/N461 , \a4/N460 ,
         \a4/N459 , \a4/N458 , \a4/N457 , \a4/N456 , \a4/N455 , \a4/N454 ,
         \a4/N453 , \a4/N452 , \a4/N451 , \a4/N450 , \a4/N449 , \a4/N448 ,
         \a4/N447 , \a4/N446 , \a4/N445 , \a4/N444 , \a4/N443 , \a4/N442 ,
         \a4/N441 , \a4/N440 , \a4/N439 , \a4/N438 , \a4/N437 , \a4/N436 ,
         \a5/N492 , \a5/N491 , \a5/N490 , \a5/N489 , \a5/N488 , \a5/N487 ,
         \a5/N486 , \a5/N485 , \a5/N484 , \a5/N483 , \a5/N482 , \a5/N481 ,
         \a5/N480 , \a5/N479 , \a5/N478 , \a5/N477 , \a5/N476 , \a5/N475 ,
         \a5/N474 , \a5/N473 , \a5/N472 , \a5/N471 , \a5/N470 , \a5/N469 ,
         \a5/N468 , \a5/N467 , \a5/N466 , \a5/N465 , \a5/N464 , \a5/N463 ,
         \a5/N462 , \a5/N461 , \a5/N460 , \a5/N459 , \a5/N458 , \a5/N457 ,
         \a5/N456 , \a5/N455 , \a5/N454 , \a5/N453 , \a5/N452 , \a5/N451 ,
         \a5/N450 , \a5/N449 , \a5/N448 , \a5/N447 , \a5/N446 , \a5/N445 ,
         \a5/N444 , \a5/N443 , \a5/N442 , \a5/N441 , \a5/N440 , \a5/N439 ,
         \a5/N438 , \a5/N437 , \a5/N436 , \a6/N492 , \a6/N491 , \a6/N490 ,
         \a6/N489 , \a6/N488 , \a6/N487 , \a6/N486 , \a6/N485 , \a6/N484 ,
         \a6/N483 , \a6/N482 , \a6/N481 , \a6/N480 , \a6/N479 , \a6/N478 ,
         \a6/N477 , \a6/N476 , \a6/N475 , \a6/N474 , \a6/N473 , \a6/N472 ,
         \a6/N471 , \a6/N470 , \a6/N469 , \a6/N468 , \a6/N467 , \a6/N466 ,
         \a6/N465 , \a6/N464 , \a6/N463 , \a6/N462 , \a6/N461 , \a6/N460 ,
         \a6/N459 , \a6/N458 , \a6/N457 , \a6/N456 , \a6/N455 , \a6/N454 ,
         \a6/N453 , \a6/N452 , \a6/N451 , \a6/N450 , \a6/N449 , \a6/N448 ,
         \a6/N447 , \a6/N446 , \a6/N445 , \a6/N444 , \a6/N443 , \a6/N442 ,
         \a6/N441 , \a6/N440 , \a6/N439 , \a6/N438 , \a6/N437 , \a6/N436 ,
         \a7/N43 , \a7/N42 , \a7/N41 , \a7/N40 , \a7/N39 , \a7/N38 , \a7/N37 ,
         \a7/N36 , \a7/N35 , \a7/N2 , \a7/N1 , \a7/N0 , n4520, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445;
  wire   [1:0] quad;
  wire   [31:0] degrees_tmp2;
  wire   [63:0] data_sin;
  wire   [63:0] data_cos;
  wire   [63:0] data_tan;
  wire   [63:0] data_csc;
  wire   [63:0] data_sec;
  wire   [63:0] data_cot;
  wire   [31:0] divider_out;
  wire   [31:0] degrees_tmp1;
  assign \a7/N2  = degrees[2];
  assign \a7/N1  = degrees[1];
  assign \a7/N0  = degrees[0];

  DFFX1 \degrees_tmp1_reg[7]  ( .D(n4528), .CLK(clock), .Q(degrees_tmp1[7]) );
  DFFX1 \degrees_tmp1_reg[6]  ( .D(n4527), .CLK(clock), .Q(degrees_tmp1[6]) );
  DFFX1 \degrees_tmp1_reg[5]  ( .D(n4526), .CLK(clock), .Q(degrees_tmp1[5]) );
  DFFX1 \degrees_tmp1_reg[4]  ( .D(n4525), .CLK(clock), .Q(degrees_tmp1[4]) );
  DFFX1 \degrees_tmp1_reg[3]  ( .D(n4524), .CLK(clock), .Q(degrees_tmp1[3]) );
  DFFX1 \degrees_tmp1_reg[2]  ( .D(n4523), .CLK(clock), .Q(degrees_tmp1[2]) );
  DFFX1 \degrees_tmp1_reg[1]  ( .D(n4522), .CLK(clock), .Q(degrees_tmp1[1]) );
  DFFX1 \degrees_tmp1_reg[0]  ( .D(n4520), .CLK(clock), .Q(degrees_tmp1[0]) );
  DFFX1 \data1_reg[63]  ( .D(N449), .CLK(clock), .Q(data1[63]) );
  DFFX1 \data1_reg[62]  ( .D(N448), .CLK(clock), .Q(data1[62]) );
  DFFX1 \data1_reg[61]  ( .D(N447), .CLK(clock), .Q(data1[61]) );
  DFFX1 \data1_reg[60]  ( .D(N446), .CLK(clock), .Q(data1[60]) );
  DFFX1 \data1_reg[59]  ( .D(N445), .CLK(clock), .Q(data1[59]) );
  DFFX1 \data1_reg[58]  ( .D(N444), .CLK(clock), .Q(data1[58]) );
  DFFX1 \data1_reg[57]  ( .D(N443), .CLK(clock), .Q(data1[57]) );
  DFFX1 \data1_reg[56]  ( .D(N442), .CLK(clock), .Q(data1[56]) );
  DFFX1 \data1_reg[55]  ( .D(N441), .CLK(clock), .Q(data1[55]) );
  DFFX1 \data1_reg[54]  ( .D(N440), .CLK(clock), .Q(data1[54]) );
  DFFX1 \data1_reg[53]  ( .D(N439), .CLK(clock), .Q(data1[53]) );
  DFFX1 \data1_reg[52]  ( .D(N438), .CLK(clock), .Q(data1[52]) );
  DFFX1 \data1_reg[51]  ( .D(N437), .CLK(clock), .Q(data1[51]) );
  DFFX1 \data1_reg[50]  ( .D(N436), .CLK(clock), .Q(data1[50]) );
  DFFX1 \data1_reg[49]  ( .D(N435), .CLK(clock), .Q(data1[49]) );
  DFFX1 \data1_reg[48]  ( .D(N434), .CLK(clock), .Q(data1[48]) );
  DFFX1 \data1_reg[47]  ( .D(N433), .CLK(clock), .Q(data1[47]) );
  DFFX1 \data1_reg[46]  ( .D(N432), .CLK(clock), .Q(data1[46]) );
  DFFX1 \data1_reg[45]  ( .D(N431), .CLK(clock), .Q(data1[45]) );
  DFFX1 \data1_reg[44]  ( .D(N430), .CLK(clock), .Q(data1[44]) );
  DFFX1 \data1_reg[43]  ( .D(N429), .CLK(clock), .Q(data1[43]) );
  DFFX1 \data1_reg[42]  ( .D(N428), .CLK(clock), .Q(data1[42]) );
  DFFX1 \data1_reg[41]  ( .D(N427), .CLK(clock), .Q(data1[41]) );
  DFFX1 \data1_reg[40]  ( .D(N426), .CLK(clock), .Q(data1[40]) );
  DFFX1 \data1_reg[39]  ( .D(N425), .CLK(clock), .Q(data1[39]) );
  DFFX1 \data1_reg[38]  ( .D(N424), .CLK(clock), .Q(data1[38]) );
  DFFX1 \data1_reg[37]  ( .D(N423), .CLK(clock), .Q(data1[37]) );
  DFFX1 \data1_reg[36]  ( .D(N422), .CLK(clock), .Q(data1[36]) );
  DFFX1 \data1_reg[35]  ( .D(N421), .CLK(clock), .Q(data1[35]) );
  DFFX1 \data1_reg[34]  ( .D(N420), .CLK(clock), .Q(data1[34]) );
  DFFX1 \data1_reg[33]  ( .D(N419), .CLK(clock), .Q(data1[33]) );
  DFFX1 \data1_reg[32]  ( .D(N418), .CLK(clock), .Q(data1[32]) );
  DFFX1 \data1_reg[31]  ( .D(N417), .CLK(clock), .Q(data1[31]) );
  DFFX1 \data1_reg[30]  ( .D(N416), .CLK(clock), .Q(data1[30]) );
  DFFX1 \data1_reg[29]  ( .D(N415), .CLK(clock), .Q(data1[29]) );
  DFFX1 \data1_reg[28]  ( .D(N414), .CLK(clock), .Q(data1[28]) );
  DFFX1 \data1_reg[27]  ( .D(N413), .CLK(clock), .Q(data1[27]) );
  DFFX1 \data1_reg[26]  ( .D(N412), .CLK(clock), .Q(data1[26]) );
  DFFX1 \data1_reg[25]  ( .D(N411), .CLK(clock), .Q(data1[25]) );
  DFFX1 \data1_reg[24]  ( .D(N410), .CLK(clock), .Q(data1[24]) );
  DFFX1 \data1_reg[23]  ( .D(N409), .CLK(clock), .Q(data1[23]) );
  DFFX1 \data1_reg[22]  ( .D(N408), .CLK(clock), .Q(data1[22]) );
  DFFX1 \data1_reg[21]  ( .D(N407), .CLK(clock), .Q(data1[21]) );
  DFFX1 \data1_reg[20]  ( .D(N406), .CLK(clock), .Q(data1[20]) );
  DFFX1 \data1_reg[19]  ( .D(N405), .CLK(clock), .Q(data1[19]) );
  DFFX1 \data1_reg[18]  ( .D(N404), .CLK(clock), .Q(data1[18]) );
  DFFX1 \data1_reg[17]  ( .D(N403), .CLK(clock), .Q(data1[17]) );
  DFFX1 \data1_reg[16]  ( .D(N402), .CLK(clock), .Q(data1[16]) );
  DFFX1 \data1_reg[15]  ( .D(N401), .CLK(clock), .Q(data1[15]) );
  DFFX1 \data1_reg[14]  ( .D(N400), .CLK(clock), .Q(data1[14]) );
  DFFX1 \data1_reg[13]  ( .D(N399), .CLK(clock), .Q(data1[13]) );
  DFFX1 \data1_reg[12]  ( .D(N398), .CLK(clock), .Q(data1[12]) );
  DFFX1 \data1_reg[11]  ( .D(N397), .CLK(clock), .Q(data1[11]) );
  DFFX1 \data1_reg[10]  ( .D(N396), .CLK(clock), .Q(data1[10]) );
  DFFX1 \data1_reg[9]  ( .D(N395), .CLK(clock), .Q(data1[9]) );
  DFFX1 \data1_reg[8]  ( .D(N394), .CLK(clock), .Q(data1[8]) );
  DFFX1 \data1_reg[7]  ( .D(N393), .CLK(clock), .Q(data1[7]) );
  DFFX1 \data1_reg[6]  ( .D(N392), .CLK(clock), .Q(data1[6]) );
  DFFX1 \data1_reg[5]  ( .D(N391), .CLK(clock), .Q(data1[5]) );
  DFFX1 \data1_reg[4]  ( .D(N390), .CLK(clock), .Q(data1[4]) );
  DFFX1 \data1_reg[3]  ( .D(N389), .CLK(clock), .Q(data1[3]) );
  DFFX1 \data1_reg[2]  ( .D(N388), .CLK(clock), .Q(data1[2]) );
  DFFX1 \data1_reg[1]  ( .D(N387), .CLK(clock), .Q(data1[1]) );
  DFFX1 \data1_reg[0]  ( .D(N386), .CLK(clock), .Q(data1[0]) );
  DFFX1 \a7/out_reg[0]  ( .D(\a7/N35 ), .CLK(clock), .Q(divider_out[0]) );
  DFFX1 \a7/out_reg[1]  ( .D(\a7/N36 ), .CLK(clock), .Q(divider_out[1]) );
  DFFX1 \a7/out_reg[2]  ( .D(\a7/N37 ), .CLK(clock), .Q(divider_out[2]) );
  DFFX1 \a7/out_reg[3]  ( .D(\a7/N38 ), .CLK(clock), .Q(divider_out[3]) );
  DFFX1 \a7/out_reg[4]  ( .D(\a7/N39 ), .CLK(clock), .Q(divider_out[4]) );
  DFFX1 \a7/out_reg[5]  ( .D(\a7/N40 ), .CLK(clock), .Q(divider_out[5]) );
  DFFX1 \a7/out_reg[6]  ( .D(\a7/N41 ), .CLK(clock), .Q(divider_out[6]), .QN(
        n9443) );
  DFFX1 \a7/out_reg[7]  ( .D(\a7/N42 ), .CLK(clock), .Q(divider_out[7]), .QN(
        n9439) );
  DFFX1 \a7/out_reg[8]  ( .D(\a7/N43 ), .CLK(clock), .Q(divider_out[8]), .QN(
        n9444) );
  DFFX1 \quad_reg[0]  ( .D(N356), .CLK(clock), .Q(quad[0]) );
  DFFX1 \degrees_tmp2_reg[2]  ( .D(N326), .CLK(clock), .Q(degrees_tmp2[2]), .QN(
        n9445) );
  DFFX1 \degrees_tmp2_reg[4]  ( .D(N328), .CLK(clock), .Q(n9434), .QN(n9440) );
  DFFX1 \degrees_tmp2_reg[5]  ( .D(N329), .CLK(clock), .Q(degrees_tmp2[5]), .QN(
        n9438) );
  DFFX1 \degrees_tmp2_reg[7]  ( .D(N331), .CLK(clock), .Q(degrees_tmp2[7]) );
  DFFX1 \degrees_tmp2_reg[0]  ( .D(N324), .CLK(clock), .Q(degrees_tmp2[0]), .QN(
        n9436) );
  DFFX1 \degrees_tmp2_reg[1]  ( .D(N325), .CLK(clock), .Q(n9435), .QN(n9442) );
  DFFX1 \degrees_tmp2_reg[3]  ( .D(N327), .CLK(clock), .Q(degrees_tmp2[3]), .QN(
        n9433) );
  DFFX1 \degrees_tmp2_reg[6]  ( .D(N330), .CLK(clock), .Q(n9437), .QN(n9441) );
  DFFX1 \degrees_tmp2_reg[8]  ( .D(N332), .CLK(clock), .Q(degrees_tmp2[8]) );
  DFFX1 \degrees_tmp2_reg[9]  ( .D(N334), .CLK(clock), .Q(degrees_tmp2[9]) );
  DFFX1 \degrees_tmp2_reg[10]  ( .D(N334), .CLK(clock), .Q(degrees_tmp2[10]) );
  DFFX1 \degrees_tmp2_reg[11]  ( .D(N334), .CLK(clock), .Q(degrees_tmp2[11]) );
  DFFX1 \degrees_tmp2_reg[12]  ( .D(N334), .CLK(clock), .Q(degrees_tmp2[12]) );
  DFFX1 \degrees_tmp2_reg[13]  ( .D(N334), .CLK(clock), .Q(degrees_tmp2[13]) );
  DFFX1 \degrees_tmp2_reg[14]  ( .D(N334), .CLK(clock), .Q(degrees_tmp2[14]) );
  DFFX1 \degrees_tmp2_reg[15]  ( .D(N334), .CLK(clock), .Q(degrees_tmp2[15]) );
  DFFX1 \degrees_tmp2_reg[16]  ( .D(N334), .CLK(clock), .Q(degrees_tmp2[16]) );
  DFFX1 \degrees_tmp2_reg[17]  ( .D(N334), .CLK(clock), .Q(degrees_tmp2[17]) );
  DFFX1 \degrees_tmp2_reg[18]  ( .D(N334), .CLK(clock), .Q(degrees_tmp2[18]) );
  DFFX1 \degrees_tmp2_reg[19]  ( .D(N334), .CLK(clock), .Q(degrees_tmp2[19]) );
  DFFX1 \degrees_tmp2_reg[20]  ( .D(N334), .CLK(clock), .Q(degrees_tmp2[20]) );
  DFFX1 \degrees_tmp2_reg[21]  ( .D(N334), .CLK(clock), .Q(degrees_tmp2[21]) );
  DFFX1 \degrees_tmp2_reg[22]  ( .D(N334), .CLK(clock), .Q(degrees_tmp2[22]) );
  DFFX1 \degrees_tmp2_reg[23]  ( .D(N334), .CLK(clock), .Q(degrees_tmp2[23]) );
  DFFX1 \degrees_tmp2_reg[24]  ( .D(N334), .CLK(clock), .Q(degrees_tmp2[24]) );
  DFFX1 \degrees_tmp2_reg[25]  ( .D(N334), .CLK(clock), .Q(degrees_tmp2[25]) );
  DFFX1 \degrees_tmp2_reg[26]  ( .D(N334), .CLK(clock), .Q(degrees_tmp2[26]) );
  DFFX1 \degrees_tmp2_reg[27]  ( .D(N334), .CLK(clock), .Q(degrees_tmp2[27]) );
  DFFX1 \degrees_tmp2_reg[28]  ( .D(N334), .CLK(clock), .Q(degrees_tmp2[28]) );
  DFFX1 \degrees_tmp2_reg[29]  ( .D(N334), .CLK(clock), .Q(degrees_tmp2[29]) );
  DFFX1 \degrees_tmp2_reg[30]  ( .D(N334), .CLK(clock), .Q(degrees_tmp2[30]) );
  DFFX1 \degrees_tmp2_reg[31]  ( .D(N334), .CLK(clock), .Q(degrees_tmp2[31]) );
  DFFX1 \a6/data_reg[62]  ( .D(\a6/N492 ), .CLK(clock), .Q(data_cot[62]) );
  DFFX1 \a4/data_reg[62]  ( .D(\a4/N492 ), .CLK(clock), .Q(data_csc[62]) );
  DFFX1 \a4/data_reg[51]  ( .D(\a4/N487 ), .CLK(clock), .Q(data_csc[51]) );
  DFFX1 \a4/data_reg[49]  ( .D(\a4/N485 ), .CLK(clock), .Q(data_csc[49]) );
  DFFX1 \a4/data_reg[50]  ( .D(\a4/N486 ), .CLK(clock), .Q(data_csc[50]) );
  DFFX1 \a5/data_reg[55]  ( .D(\a5/N491 ), .CLK(clock), .Q(data_sec[55]) );
  DFFX1 \a5/data_reg[56]  ( .D(\a5/N491 ), .CLK(clock), .Q(data_sec[56]) );
  DFFX1 \a5/data_reg[57]  ( .D(\a5/N491 ), .CLK(clock), .Q(data_sec[57]) );
  DFFX1 \a5/data_reg[58]  ( .D(\a5/N491 ), .CLK(clock), .Q(data_sec[58]) );
  DFFX1 \a5/data_reg[59]  ( .D(\a5/N491 ), .CLK(clock), .Q(data_sec[59]) );
  DFFX1 \a5/data_reg[60]  ( .D(\a5/N491 ), .CLK(clock), .Q(data_sec[60]) );
  DFFX1 \a5/data_reg[61]  ( .D(\a5/N491 ), .CLK(clock), .Q(data_sec[61]) );
  DFFX1 \a3/data_reg[55]  ( .D(\a3/N491 ), .CLK(clock), .Q(data_tan[55]) );
  DFFX1 \a3/data_reg[56]  ( .D(\a3/N491 ), .CLK(clock), .Q(data_tan[56]) );
  DFFX1 \a3/data_reg[57]  ( .D(\a3/N491 ), .CLK(clock), .Q(data_tan[57]) );
  DFFX1 \a3/data_reg[58]  ( .D(\a3/N491 ), .CLK(clock), .Q(data_tan[58]) );
  DFFX1 \a3/data_reg[59]  ( .D(\a3/N491 ), .CLK(clock), .Q(data_tan[59]) );
  DFFX1 \a3/data_reg[60]  ( .D(\a3/N491 ), .CLK(clock), .Q(data_tan[60]) );
  DFFX1 \a3/data_reg[61]  ( .D(\a3/N491 ), .CLK(clock), .Q(data_tan[61]) );
  DFFX1 \a3/data_reg[35]  ( .D(\a3/N471 ), .CLK(clock), .Q(data_tan[35]) );
  DFFX1 \a5/data_reg[54]  ( .D(\a5/N490 ), .CLK(clock), .Q(data_sec[54]) );
  DFFX1 \a3/data_reg[54]  ( .D(\a3/N490 ), .CLK(clock), .Q(data_tan[54]) );
  DFFX1 \a2/data_reg[55]  ( .D(\a2/N490 ), .CLK(clock), .Q(data_cos[55]) );
  DFFX1 \a2/data_reg[56]  ( .D(\a2/N490 ), .CLK(clock), .Q(data_cos[56]) );
  DFFX1 \a2/data_reg[57]  ( .D(\a2/N490 ), .CLK(clock), .Q(data_cos[57]) );
  DFFX1 \a2/data_reg[58]  ( .D(\a2/N490 ), .CLK(clock), .Q(data_cos[58]) );
  DFFX1 \a2/data_reg[59]  ( .D(\a2/N490 ), .CLK(clock), .Q(data_cos[59]) );
  DFFX1 \a2/data_reg[60]  ( .D(\a2/N490 ), .CLK(clock), .Q(data_cos[60]) );
  DFFX1 \a2/data_reg[61]  ( .D(\a2/N490 ), .CLK(clock), .Q(data_cos[61]) );
  DFFX1 \a3/data_reg[9]  ( .D(\a3/N445 ), .CLK(clock), .Q(data_tan[9]) );
  DFFX1 \a6/data_reg[0]  ( .D(\a6/N436 ), .CLK(clock), .Q(data_cot[0]) );
  DFFX1 \a2/data_reg[40]  ( .D(\a2/N475 ), .CLK(clock), .Q(data_cos[40]) );
  DFFX1 \a2/data_reg[21]  ( .D(\a2/N456 ), .CLK(clock), .Q(data_cos[21]) );
  DFFX1 \a3/data_reg[44]  ( .D(\a3/N480 ), .CLK(clock), .Q(data_tan[44]) );
  DFFX1 \a6/data_reg[36]  ( .D(\a6/N472 ), .CLK(clock), .Q(data_cot[36]) );
  DFFX1 \a4/data_reg[15]  ( .D(\a4/N451 ), .CLK(clock), .Q(data_csc[15]) );
  DFFX1 \a2/data_reg[34]  ( .D(\a2/N469 ), .CLK(clock), .Q(data_cos[34]) );
  DFFX1 \a3/data_reg[34]  ( .D(\a3/N470 ), .CLK(clock), .Q(data_tan[34]) );
  DFFX1 \a2/data_reg[10]  ( .D(\a2/N445 ), .CLK(clock), .Q(data_cos[10]) );
  DFFX1 \a6/data_reg[33]  ( .D(\a6/N469 ), .CLK(clock), .Q(data_cot[33]) );
  DFFX1 \a6/data_reg[44]  ( .D(\a6/N480 ), .CLK(clock), .Q(data_cot[44]) );
  DFFX1 \a2/data_reg[9]  ( .D(\a2/N444 ), .CLK(clock), .Q(data_cos[9]) );
  DFFX1 \a2/data_reg[20]  ( .D(\a2/N455 ), .CLK(clock), .Q(data_cos[20]) );
  DFFX1 \a6/data_reg[13]  ( .D(\a6/N449 ), .CLK(clock), .Q(data_cot[13]) );
  DFFX1 \a2/data_reg[33]  ( .D(\a2/N468 ), .CLK(clock), .Q(data_cos[33]) );
  DFFX1 \a6/data_reg[51]  ( .D(\a6/N487 ), .CLK(clock), .Q(data_cot[51]) );
  DFFX1 \a4/data_reg[10]  ( .D(\a4/N446 ), .CLK(clock), .Q(data_csc[10]) );
  DFFX1 \a3/data_reg[4]  ( .D(\a3/N440 ), .CLK(clock), .Q(data_tan[4]) );
  DFFX1 \a6/data_reg[15]  ( .D(\a6/N451 ), .CLK(clock), .Q(data_cot[15]) );
  DFFX1 \a5/data_reg[15]  ( .D(\a5/N451 ), .CLK(clock), .Q(data_sec[15]) );
  DFFX1 \a4/data_reg[30]  ( .D(\a4/N466 ), .CLK(clock), .Q(data_csc[30]) );
  DFFX1 \a2/data_reg[6]  ( .D(\a2/N441 ), .CLK(clock), .Q(data_cos[6]) );
  DFFX1 \a5/data_reg[14]  ( .D(\a5/N450 ), .CLK(clock), .Q(data_sec[14]) );
  DFFX1 \a5/data_reg[52]  ( .D(\a5/N488 ), .CLK(clock), .Q(data_sec[52]) );
  DFFX1 \a3/data_reg[52]  ( .D(\a3/N488 ), .CLK(clock), .Q(data_tan[52]) );
  DFFX1 \a2/data_reg[2]  ( .D(\a2/N437 ), .CLK(clock), .Q(data_cos[2]) );
  DFFX1 \a2/data_reg[23]  ( .D(\a2/N458 ), .CLK(clock), .Q(data_cos[23]) );
  DFFX1 \a1/data_reg[16]  ( .D(\a1/N451 ), .CLK(clock), .Q(data_sin[16]) );
  DFFX1 \a1/data_reg[52]  ( .D(\a1/N487 ), .CLK(clock), .Q(data_sin[52]) );
  DFFX1 \a3/data_reg[36]  ( .D(\a3/N472 ), .CLK(clock), .Q(data_tan[36]) );
  DFFX1 \a6/data_reg[22]  ( .D(\a6/N458 ), .CLK(clock), .Q(data_cot[22]) );
  DFFX1 \a5/data_reg[26]  ( .D(\a5/N462 ), .CLK(clock), .Q(data_sec[26]) );
  DFFX1 \a4/data_reg[8]  ( .D(\a4/N444 ), .CLK(clock), .Q(data_csc[8]) );
  DFFX1 \a6/data_reg[53]  ( .D(\a6/N489 ), .CLK(clock), .Q(data_cot[53]) );
  DFFX1 \a1/data_reg[30]  ( .D(\a1/N465 ), .CLK(clock), .Q(data_sin[30]) );
  DFFX1 \a3/data_reg[45]  ( .D(\a3/N481 ), .CLK(clock), .Q(data_tan[45]) );
  DFFX1 \a1/data_reg[31]  ( .D(\a1/N466 ), .CLK(clock), .Q(data_sin[31]) );
  DFFX1 \a5/data_reg[42]  ( .D(\a5/N478 ), .CLK(clock), .Q(data_sec[42]) );
  DFFX1 \a5/data_reg[4]  ( .D(\a5/N440 ), .CLK(clock), .Q(data_sec[4]) );
  DFFX1 \a4/data_reg[11]  ( .D(\a4/N447 ), .CLK(clock), .Q(data_csc[11]) );
  DFFX1 \a4/data_reg[48]  ( .D(\a4/N484 ), .CLK(clock), .Q(data_csc[48]) );
  DFFX1 \a2/data_reg[11]  ( .D(\a2/N446 ), .CLK(clock), .Q(data_cos[11]) );
  DFFX1 \a6/data_reg[54]  ( .D(\a6/N490 ), .CLK(clock), .Q(data_cot[54]) );
  DFFX1 \a3/data_reg[5]  ( .D(\a3/N441 ), .CLK(clock), .Q(data_tan[5]) );
  DFFX1 \a3/data_reg[32]  ( .D(\a3/N468 ), .CLK(clock), .Q(data_tan[32]) );
  DFFX1 \a2/data_reg[38]  ( .D(\a2/N473 ), .CLK(clock), .Q(data_cos[38]) );
  DFFX1 \a5/data_reg[0]  ( .D(\a5/N436 ), .CLK(clock), .Q(data_sec[0]) );
  DFFX1 \a2/data_reg[45]  ( .D(\a2/N480 ), .CLK(clock), .Q(data_cos[45]) );
  DFFX1 \a4/data_reg[43]  ( .D(\a4/N479 ), .CLK(clock), .Q(data_csc[43]) );
  DFFX1 \a2/data_reg[50]  ( .D(\a2/N485 ), .CLK(clock), .Q(data_cos[50]) );
  DFFX1 \a5/data_reg[21]  ( .D(\a5/N457 ), .CLK(clock), .Q(data_sec[21]) );
  DFFX1 \a5/data_reg[44]  ( .D(\a5/N480 ), .CLK(clock), .Q(data_sec[44]) );
  DFFX1 \a4/data_reg[38]  ( .D(\a4/N474 ), .CLK(clock), .Q(data_csc[38]) );
  DFFX1 \a6/data_reg[1]  ( .D(\a6/N437 ), .CLK(clock), .Q(data_cot[1]) );
  DFFX1 \a5/data_reg[35]  ( .D(\a5/N471 ), .CLK(clock), .Q(data_sec[35]) );
  DFFX1 \a4/data_reg[21]  ( .D(\a4/N457 ), .CLK(clock), .Q(data_csc[21]) );
  DFFX1 \a3/data_reg[11]  ( .D(\a3/N447 ), .CLK(clock), .Q(data_tan[11]) );
  DFFX1 \a2/data_reg[22]  ( .D(\a2/N457 ), .CLK(clock), .Q(data_cos[22]) );
  DFFX1 \a2/data_reg[41]  ( .D(\a2/N476 ), .CLK(clock), .Q(data_cos[41]) );
  DFFX1 \a6/data_reg[42]  ( .D(\a6/N478 ), .CLK(clock), .Q(data_cot[42]) );
  DFFX1 \a4/data_reg[33]  ( .D(\a4/N469 ), .CLK(clock), .Q(data_csc[33]) );
  DFFX1 \a4/data_reg[35]  ( .D(\a4/N471 ), .CLK(clock), .Q(data_csc[35]) );
  DFFX1 \a4/data_reg[44]  ( .D(\a4/N480 ), .CLK(clock), .Q(data_csc[44]) );
  DFFX1 \a6/data_reg[7]  ( .D(\a6/N443 ), .CLK(clock), .Q(data_cot[7]) );
  DFFX1 \a6/data_reg[8]  ( .D(\a6/N444 ), .CLK(clock), .Q(data_cot[8]) );
  DFFX1 \a3/data_reg[16]  ( .D(\a3/N452 ), .CLK(clock), .Q(data_tan[16]) );
  DFFX1 \a6/data_reg[18]  ( .D(\a6/N454 ), .CLK(clock), .Q(data_cot[18]) );
  DFFX1 \a5/data_reg[20]  ( .D(\a5/N456 ), .CLK(clock), .Q(data_sec[20]) );
  DFFX1 \a6/data_reg[31]  ( .D(\a6/N467 ), .CLK(clock), .Q(data_cot[31]) );
  DFFX1 \a6/data_reg[38]  ( .D(\a6/N474 ), .CLK(clock), .Q(data_cot[38]) );
  DFFX1 \a1/data_reg[22]  ( .D(\a1/N457 ), .CLK(clock), .Q(data_sin[22]) );
  DFFX1 \a3/data_reg[51]  ( .D(\a3/N487 ), .CLK(clock), .Q(data_tan[51]) );
  DFFX1 \a5/data_reg[9]  ( .D(\a5/N445 ), .CLK(clock), .Q(data_sec[9]) );
  DFFX1 \a5/data_reg[30]  ( .D(\a5/N466 ), .CLK(clock), .Q(data_sec[30]) );
  DFFX1 \a4/data_reg[19]  ( .D(\a4/N455 ), .CLK(clock), .Q(data_csc[19]) );
  DFFX1 \a6/data_reg[10]  ( .D(\a6/N446 ), .CLK(clock), .Q(data_cot[10]) );
  DFFX1 \a1/data_reg[2]  ( .D(\a1/N437 ), .CLK(clock), .Q(data_sin[2]) );
  DFFX1 \a6/data_reg[9]  ( .D(\a6/N445 ), .CLK(clock), .Q(data_cot[9]) );
  DFFX1 \a3/data_reg[50]  ( .D(\a3/N486 ), .CLK(clock), .Q(data_tan[50]) );
  DFFX1 \a1/data_reg[32]  ( .D(\a1/N467 ), .CLK(clock), .Q(data_sin[32]) );
  DFFX1 \a6/data_reg[20]  ( .D(\a6/N456 ), .CLK(clock), .Q(data_cot[20]) );
  DFFX1 \a4/data_reg[45]  ( .D(\a4/N481 ), .CLK(clock), .Q(data_csc[45]) );
  DFFX1 \a2/data_reg[4]  ( .D(\a2/N439 ), .CLK(clock), .Q(data_cos[4]) );
  DFFX1 \a2/data_reg[7]  ( .D(\a2/N442 ), .CLK(clock), .Q(data_cos[7]) );
  DFFX1 \a2/data_reg[13]  ( .D(\a2/N448 ), .CLK(clock), .Q(data_cos[13]) );
  DFFX1 \a6/data_reg[37]  ( .D(\a6/N473 ), .CLK(clock), .Q(data_cot[37]) );
  DFFX1 \a4/data_reg[16]  ( .D(\a4/N452 ), .CLK(clock), .Q(data_csc[16]) );
  DFFX1 \a3/data_reg[15]  ( .D(\a3/N451 ), .CLK(clock), .Q(data_tan[15]) );
  DFFX1 \a3/data_reg[48]  ( .D(\a3/N484 ), .CLK(clock), .Q(data_tan[48]) );
  DFFX1 \a3/data_reg[7]  ( .D(\a3/N443 ), .CLK(clock), .Q(data_tan[7]) );
  DFFX1 \a5/data_reg[12]  ( .D(\a5/N448 ), .CLK(clock), .Q(data_sec[12]) );
  DFFX1 \a4/data_reg[6]  ( .D(\a4/N442 ), .CLK(clock), .Q(data_csc[6]) );
  DFFX1 \a4/data_reg[13]  ( .D(\a4/N449 ), .CLK(clock), .Q(data_csc[13]) );
  DFFX1 \a4/data_reg[12]  ( .D(\a4/N448 ), .CLK(clock), .Q(data_csc[12]) );
  DFFX1 \a4/data_reg[24]  ( .D(\a4/N460 ), .CLK(clock), .Q(data_csc[24]) );
  DFFX1 \a3/data_reg[10]  ( .D(\a3/N446 ), .CLK(clock), .Q(data_tan[10]) );
  DFFX1 \a3/data_reg[13]  ( .D(\a3/N449 ), .CLK(clock), .Q(data_tan[13]) );
  DFFX1 \a3/data_reg[29]  ( .D(\a3/N465 ), .CLK(clock), .Q(data_tan[29]) );
  DFFX1 \a5/data_reg[19]  ( .D(\a5/N455 ), .CLK(clock), .Q(data_sec[19]) );
  DFFX1 \a3/data_reg[24]  ( .D(\a3/N460 ), .CLK(clock), .Q(data_tan[24]) );
  DFFX1 \a2/data_reg[1]  ( .D(\a2/N436 ), .CLK(clock), .Q(data_cos[1]) );
  DFFX1 \a2/data_reg[30]  ( .D(\a2/N465 ), .CLK(clock), .Q(data_cos[30]) );
  DFFX1 \a6/data_reg[4]  ( .D(\a6/N440 ), .CLK(clock), .Q(data_cot[4]) );
  DFFX1 \a2/data_reg[36]  ( .D(\a2/N471 ), .CLK(clock), .Q(data_cos[36]) );
  DFFX1 \a2/data_reg[51]  ( .D(\a2/N486 ), .CLK(clock), .Q(data_cos[51]) );
  DFFX1 \a1/data_reg[38]  ( .D(\a1/N473 ), .CLK(clock), .Q(data_sin[38]) );
  DFFX1 \a6/data_reg[2]  ( .D(\a6/N438 ), .CLK(clock), .Q(data_cot[2]) );
  DFFX1 \a4/data_reg[0]  ( .D(\a4/N436 ), .CLK(clock), .Q(data_csc[0]) );
  DFFX1 \a4/data_reg[28]  ( .D(\a4/N464 ), .CLK(clock), .Q(data_csc[28]) );
  DFFX1 \a3/data_reg[20]  ( .D(\a3/N456 ), .CLK(clock), .Q(data_tan[20]) );
  DFFX1 \a2/data_reg[19]  ( .D(\a2/N454 ), .CLK(clock), .Q(data_cos[19]) );
  DFFX1 \a1/data_reg[1]  ( .D(\a1/N436 ), .CLK(clock), .Q(data_sin[1]) );
  DFFX1 \a5/data_reg[23]  ( .D(\a5/N459 ), .CLK(clock), .Q(data_sec[23]) );
  DFFX1 \a6/data_reg[27]  ( .D(\a6/N463 ), .CLK(clock), .Q(data_cot[27]) );
  DFFX1 \a4/data_reg[22]  ( .D(\a4/N458 ), .CLK(clock), .Q(data_csc[22]) );
  DFFX1 \a4/data_reg[39]  ( .D(\a4/N475 ), .CLK(clock), .Q(data_csc[39]) );
  DFFX1 \a2/data_reg[46]  ( .D(\a2/N481 ), .CLK(clock), .Q(data_cos[46]) );
  DFFX1 \a2/data_reg[48]  ( .D(\a2/N483 ), .CLK(clock), .Q(data_cos[48]) );
  DFFX1 \a1/data_reg[12]  ( .D(\a1/N447 ), .CLK(clock), .Q(data_sin[12]) );
  DFFX1 \a5/data_reg[43]  ( .D(\a5/N479 ), .CLK(clock), .Q(data_sec[43]) );
  DFFX1 \a2/data_reg[25]  ( .D(\a2/N460 ), .CLK(clock), .Q(data_cos[25]) );
  DFFX1 \a3/data_reg[33]  ( .D(\a3/N469 ), .CLK(clock), .Q(data_tan[33]) );
  DFFX1 \a2/data_reg[0]  ( .D(\a2/N435 ), .CLK(clock), .Q(data_cos[0]) );
  DFFX1 \a2/data_reg[26]  ( .D(\a2/N461 ), .CLK(clock), .Q(data_cos[26]) );
  DFFX1 \a6/data_reg[47]  ( .D(\a6/N483 ), .CLK(clock), .Q(data_cot[47]) );
  DFFX1 \a5/data_reg[11]  ( .D(\a5/N447 ), .CLK(clock), .Q(data_sec[11]) );
  DFFX1 \a2/data_reg[12]  ( .D(\a2/N447 ), .CLK(clock), .Q(data_cos[12]) );
  DFFX1 \a1/data_reg[42]  ( .D(\a1/N477 ), .CLK(clock), .Q(data_sin[42]) );
  DFFX1 \a4/data_reg[5]  ( .D(\a4/N441 ), .CLK(clock), .Q(data_csc[5]) );
  DFFX1 \a4/data_reg[29]  ( .D(\a4/N465 ), .CLK(clock), .Q(data_csc[29]) );
  DFFX1 \a3/data_reg[14]  ( .D(\a3/N450 ), .CLK(clock), .Q(data_tan[14]) );
  DFFX1 \a3/data_reg[38]  ( .D(\a3/N474 ), .CLK(clock), .Q(data_tan[38]) );
  DFFX1 \a4/data_reg[9]  ( .D(\a4/N445 ), .CLK(clock), .Q(data_csc[9]) );
  DFFX1 \a6/data_reg[52]  ( .D(\a6/N488 ), .CLK(clock), .Q(data_cot[52]) );
  DFFX1 \a2/data_reg[52]  ( .D(\a2/N487 ), .CLK(clock), .Q(data_cos[52]) );
  DFFX1 \a6/data_reg[41]  ( .D(\a6/N477 ), .CLK(clock), .Q(data_cot[41]) );
  DFFX1 \a5/data_reg[8]  ( .D(\a5/N444 ), .CLK(clock), .Q(data_sec[8]) );
  DFFX1 \a5/data_reg[13]  ( .D(\a5/N449 ), .CLK(clock), .Q(data_sec[13]) );
  DFFX1 \a5/data_reg[24]  ( .D(\a5/N460 ), .CLK(clock), .Q(data_sec[24]) );
  DFFX1 \a5/data_reg[27]  ( .D(\a5/N463 ), .CLK(clock), .Q(data_sec[27]) );
  DFFX1 \a5/data_reg[34]  ( .D(\a5/N470 ), .CLK(clock), .Q(data_sec[34]) );
  DFFX1 \a4/data_reg[4]  ( .D(\a4/N440 ), .CLK(clock), .Q(data_csc[4]) );
  DFFX1 \a2/data_reg[3]  ( .D(\a2/N438 ), .CLK(clock), .Q(data_cos[3]) );
  DFFX1 \a2/data_reg[39]  ( .D(\a2/N474 ), .CLK(clock), .Q(data_cos[39]) );
  DFFX1 \a1/data_reg[14]  ( .D(\a1/N449 ), .CLK(clock), .Q(data_sin[14]) );
  DFFX1 \a6/data_reg[26]  ( .D(\a6/N462 ), .CLK(clock), .Q(data_cot[26]) );
  DFFX1 \a1/data_reg[29]  ( .D(\a1/N464 ), .CLK(clock), .Q(data_sin[29]) );
  DFFX1 \a3/data_reg[43]  ( .D(\a3/N479 ), .CLK(clock), .Q(data_tan[43]) );
  DFFX1 \a1/data_reg[34]  ( .D(\a1/N469 ), .CLK(clock), .Q(data_sin[34]) );
  DFFX1 \a3/data_reg[8]  ( .D(\a3/N444 ), .CLK(clock), .Q(data_tan[8]) );
  DFFX1 \a1/data_reg[4]  ( .D(\a1/N439 ), .CLK(clock), .Q(data_sin[4]) );
  DFFX1 \a1/data_reg[27]  ( .D(\a1/N462 ), .CLK(clock), .Q(data_sin[27]) );
  DFFX1 \a6/data_reg[17]  ( .D(\a6/N453 ), .CLK(clock), .Q(data_cot[17]) );
  DFFX1 \a6/data_reg[29]  ( .D(\a6/N465 ), .CLK(clock), .Q(data_cot[29]) );
  DFFX1 \a4/data_reg[31]  ( .D(\a4/N467 ), .CLK(clock), .Q(data_csc[31]) );
  DFFX1 \a3/data_reg[2]  ( .D(\a3/N438 ), .CLK(clock), .Q(data_tan[2]) );
  DFFX1 \a3/data_reg[19]  ( .D(\a3/N455 ), .CLK(clock), .Q(data_tan[19]) );
  DFFX1 \a3/data_reg[22]  ( .D(\a3/N458 ), .CLK(clock), .Q(data_tan[22]) );
  DFFX1 \a3/data_reg[27]  ( .D(\a3/N463 ), .CLK(clock), .Q(data_tan[27]) );
  DFFX1 \a3/data_reg[39]  ( .D(\a3/N475 ), .CLK(clock), .Q(data_tan[39]) );
  DFFX1 \a1/data_reg[7]  ( .D(\a1/N442 ), .CLK(clock), .Q(data_sin[7]) );
  DFFX1 \a6/data_reg[35]  ( .D(\a6/N471 ), .CLK(clock), .Q(data_cot[35]) );
  DFFX1 \a2/data_reg[35]  ( .D(\a2/N470 ), .CLK(clock), .Q(data_cos[35]) );
  DFFX1 \a1/data_reg[25]  ( .D(\a1/N460 ), .CLK(clock), .Q(data_sin[25]) );
  DFFX1 \a6/data_reg[43]  ( .D(\a6/N479 ), .CLK(clock), .Q(data_cot[43]) );
  DFFX1 \a2/data_reg[31]  ( .D(\a2/N466 ), .CLK(clock), .Q(data_cos[31]) );
  DFFX1 \a6/data_reg[32]  ( .D(\a6/N468 ), .CLK(clock), .Q(data_cot[32]) );
  DFFX1 \a5/data_reg[51]  ( .D(\a5/N487 ), .CLK(clock), .Q(data_sec[51]) );
  DFFX1 \a3/data_reg[26]  ( .D(\a3/N462 ), .CLK(clock), .Q(data_tan[26]) );
  DFFX1 \a2/data_reg[37]  ( .D(\a2/N472 ), .CLK(clock), .Q(data_cos[37]) );
  DFFX1 \a2/data_reg[44]  ( .D(\a2/N479 ), .CLK(clock), .Q(data_cos[44]) );
  DFFX1 \a2/data_reg[47]  ( .D(\a2/N482 ), .CLK(clock), .Q(data_cos[47]) );
  DFFX1 \a5/data_reg[2]  ( .D(\a5/N438 ), .CLK(clock), .Q(data_sec[2]) );
  DFFX1 \a5/data_reg[5]  ( .D(\a5/N441 ), .CLK(clock), .Q(data_sec[5]) );
  DFFX1 \a5/data_reg[18]  ( .D(\a5/N454 ), .CLK(clock), .Q(data_sec[18]) );
  DFFX1 \a5/data_reg[40]  ( .D(\a5/N476 ), .CLK(clock), .Q(data_sec[40]) );
  DFFX1 \a5/data_reg[47]  ( .D(\a5/N483 ), .CLK(clock), .Q(data_sec[47]) );
  DFFX1 \a1/data_reg[6]  ( .D(\a1/N441 ), .CLK(clock), .Q(data_sin[6]) );
  DFFX1 \a1/data_reg[8]  ( .D(\a1/N443 ), .CLK(clock), .Q(data_sin[8]) );
  DFFX1 \a5/data_reg[50]  ( .D(\a5/N486 ), .CLK(clock), .Q(data_sec[50]) );
  DFFX1 \a4/data_reg[25]  ( .D(\a4/N461 ), .CLK(clock), .Q(data_csc[25]) );
  DFFX1 \a4/data_reg[32]  ( .D(\a4/N468 ), .CLK(clock), .Q(data_csc[32]) );
  DFFX1 \a2/data_reg[5]  ( .D(\a2/N440 ), .CLK(clock), .Q(data_cos[5]) );
  DFFX1 \a6/data_reg[6]  ( .D(\a6/N442 ), .CLK(clock), .Q(data_cot[6]) );
  DFFX1 \a6/data_reg[48]  ( .D(\a6/N484 ), .CLK(clock), .Q(data_cot[48]) );
  DFFX1 \a5/data_reg[31]  ( .D(\a5/N467 ), .CLK(clock), .Q(data_sec[31]) );
  DFFX1 \a3/data_reg[30]  ( .D(\a3/N466 ), .CLK(clock), .Q(data_tan[30]) );
  DFFX1 \a5/data_reg[1]  ( .D(\a5/N437 ), .CLK(clock), .Q(data_sec[1]) );
  DFFX1 \a6/data_reg[24]  ( .D(\a6/N460 ), .CLK(clock), .Q(data_cot[24]) );
  DFFX1 \a6/data_reg[30]  ( .D(\a6/N466 ), .CLK(clock), .Q(data_cot[30]) );
  DFFX1 \a5/data_reg[3]  ( .D(\a5/N439 ), .CLK(clock), .Q(data_sec[3]) );
  DFFX1 \a4/data_reg[7]  ( .D(\a4/N443 ), .CLK(clock), .Q(data_csc[7]) );
  DFFX1 \a4/data_reg[36]  ( .D(\a4/N472 ), .CLK(clock), .Q(data_csc[36]) );
  DFFX1 \a4/data_reg[40]  ( .D(\a4/N476 ), .CLK(clock), .Q(data_csc[40]) );
  DFFX1 \a4/data_reg[46]  ( .D(\a4/N482 ), .CLK(clock), .Q(data_csc[46]) );
  DFFX1 \a2/data_reg[28]  ( .D(\a2/N463 ), .CLK(clock), .Q(data_cos[28]) );
  DFFX1 \a2/data_reg[29]  ( .D(\a2/N464 ), .CLK(clock), .Q(data_cos[29]) );
  DFFX1 \a2/data_reg[32]  ( .D(\a2/N467 ), .CLK(clock), .Q(data_cos[32]) );
  DFFX1 \a2/data_reg[43]  ( .D(\a2/N478 ), .CLK(clock), .Q(data_cos[43]) );
  DFFX1 \a1/data_reg[11]  ( .D(\a1/N446 ), .CLK(clock), .Q(data_sin[11]) );
  DFFX1 \a1/data_reg[24]  ( .D(\a1/N459 ), .CLK(clock), .Q(data_sin[24]) );
  DFFX1 \a5/data_reg[37]  ( .D(\a5/N473 ), .CLK(clock), .Q(data_sec[37]) );
  DFFX1 \a5/data_reg[41]  ( .D(\a5/N477 ), .CLK(clock), .Q(data_sec[41]) );
  DFFX1 \a2/data_reg[42]  ( .D(\a2/N477 ), .CLK(clock), .Q(data_cos[42]) );
  DFFX1 \a1/data_reg[18]  ( .D(\a1/N453 ), .CLK(clock), .Q(data_sin[18]) );
  DFFX1 \a1/data_reg[41]  ( .D(\a1/N476 ), .CLK(clock), .Q(data_sin[41]) );
  DFFX1 \a6/data_reg[49]  ( .D(\a6/N485 ), .CLK(clock), .Q(data_cot[49]) );
  DFFX1 \a5/data_reg[16]  ( .D(\a5/N452 ), .CLK(clock), .Q(data_sec[16]) );
  DFFX1 \a3/data_reg[41]  ( .D(\a3/N477 ), .CLK(clock), .Q(data_tan[41]) );
  DFFX1 \a1/data_reg[13]  ( .D(\a1/N448 ), .CLK(clock), .Q(data_sin[13]) );
  DFFX1 \a6/data_reg[23]  ( .D(\a6/N459 ), .CLK(clock), .Q(data_cot[23]) );
  DFFX1 \a5/data_reg[33]  ( .D(\a5/N469 ), .CLK(clock), .Q(data_sec[33]) );
  DFFX1 \a3/data_reg[53]  ( .D(\a3/N489 ), .CLK(clock), .Q(data_tan[53]) );
  DFFX1 \a2/data_reg[15]  ( .D(\a2/N450 ), .CLK(clock), .Q(data_cos[15]) );
  DFFX1 \a3/data_reg[17]  ( .D(\a3/N453 ), .CLK(clock), .Q(data_tan[17]) );
  DFFX1 \a3/data_reg[47]  ( .D(\a3/N483 ), .CLK(clock), .Q(data_tan[47]) );
  DFFX1 \a5/data_reg[25]  ( .D(\a5/N461 ), .CLK(clock), .Q(data_sec[25]) );
  DFFX1 \a4/data_reg[3]  ( .D(\a4/N439 ), .CLK(clock), .Q(data_csc[3]) );
  DFFX1 \a1/data_reg[5]  ( .D(\a1/N440 ), .CLK(clock), .Q(data_sin[5]) );
  DFFX1 \a1/data_reg[33]  ( .D(\a1/N468 ), .CLK(clock), .Q(data_sin[33]) );
  DFFX1 \a1/data_reg[45]  ( .D(\a1/N480 ), .CLK(clock), .Q(data_sin[45]) );
  DFFX1 \a1/data_reg[17]  ( .D(\a1/N452 ), .CLK(clock), .Q(data_sin[17]) );
  DFFX1 \a1/data_reg[37]  ( .D(\a1/N472 ), .CLK(clock), .Q(data_sin[37]) );
  DFFX1 \a5/data_reg[6]  ( .D(\a5/N442 ), .CLK(clock), .Q(data_sec[6]) );
  DFFX1 \a4/data_reg[27]  ( .D(\a4/N463 ), .CLK(clock), .Q(data_csc[27]) );
  DFFX1 \a3/data_reg[21]  ( .D(\a3/N457 ), .CLK(clock), .Q(data_tan[21]) );
  DFFX1 \a3/data_reg[23]  ( .D(\a3/N459 ), .CLK(clock), .Q(data_tan[23]) );
  DFFX1 \a2/data_reg[8]  ( .D(\a2/N443 ), .CLK(clock), .Q(data_cos[8]) );
  DFFX1 \a2/data_reg[49]  ( .D(\a2/N484 ), .CLK(clock), .Q(data_cos[49]) );
  DFFX1 \a1/data_reg[26]  ( .D(\a1/N461 ), .CLK(clock), .Q(data_sin[26]) );
  DFFX1 \a1/data_reg[28]  ( .D(\a1/N463 ), .CLK(clock), .Q(data_sin[28]) );
  DFFX1 \a3/data_reg[25]  ( .D(\a3/N461 ), .CLK(clock), .Q(data_tan[25]) );
  DFFX1 \a2/data_reg[14]  ( .D(\a2/N449 ), .CLK(clock), .Q(data_cos[14]) );
  DFFX1 \a2/data_reg[16]  ( .D(\a2/N451 ), .CLK(clock), .Q(data_cos[16]) );
  DFFX1 \a1/data_reg[46]  ( .D(\a1/N481 ), .CLK(clock), .Q(data_sin[46]) );
  DFFX1 \a1/data_reg[23]  ( .D(\a1/N458 ), .CLK(clock), .Q(data_sin[23]) );
  DFFX1 \a6/data_reg[28]  ( .D(\a6/N464 ), .CLK(clock), .Q(data_cot[28]) );
  DFFX1 \a6/data_reg[45]  ( .D(\a6/N481 ), .CLK(clock), .Q(data_cot[45]) );
  DFFX1 \a5/data_reg[39]  ( .D(\a5/N475 ), .CLK(clock), .Q(data_sec[39]) );
  DFFX1 \a5/data_reg[48]  ( .D(\a5/N484 ), .CLK(clock), .Q(data_sec[48]) );
  DFFX1 \a5/data_reg[49]  ( .D(\a5/N485 ), .CLK(clock), .Q(data_sec[49]) );
  DFFX1 \a4/data_reg[23]  ( .D(\a4/N459 ), .CLK(clock), .Q(data_csc[23]) );
  DFFX1 \a4/data_reg[34]  ( .D(\a4/N470 ), .CLK(clock), .Q(data_csc[34]) );
  DFFX1 \a3/data_reg[42]  ( .D(\a3/N478 ), .CLK(clock), .Q(data_tan[42]) );
  DFFX1 \a2/data_reg[27]  ( .D(\a2/N462 ), .CLK(clock), .Q(data_cos[27]) );
  DFFX1 \a1/data_reg[36]  ( .D(\a1/N471 ), .CLK(clock), .Q(data_sin[36]) );
  DFFX1 \a1/data_reg[40]  ( .D(\a1/N475 ), .CLK(clock), .Q(data_sin[40]) );
  DFFX1 \a1/data_reg[10]  ( .D(\a1/N445 ), .CLK(clock), .Q(data_sin[10]) );
  DFFX1 \a1/data_reg[47]  ( .D(\a1/N482 ), .CLK(clock), .Q(data_sin[47]) );
  DFFX1 \a1/data_reg[48]  ( .D(\a1/N483 ), .CLK(clock), .Q(data_sin[48]) );
  DFFX1 \a6/data_reg[11]  ( .D(\a6/N447 ), .CLK(clock), .Q(data_cot[11]) );
  DFFX1 \a5/data_reg[22]  ( .D(\a5/N458 ), .CLK(clock), .Q(data_sec[22]) );
  DFFX1 \a1/data_reg[49]  ( .D(\a1/N484 ), .CLK(clock), .Q(data_sin[49]) );
  DFFX1 \a3/data_reg[12]  ( .D(\a3/N448 ), .CLK(clock), .Q(data_tan[12]) );
  DFFX1 \a3/data_reg[46]  ( .D(\a3/N482 ), .CLK(clock), .Q(data_tan[46]) );
  DFFX1 \a1/data_reg[20]  ( .D(\a1/N455 ), .CLK(clock), .Q(data_sin[20]) );
  DFFX1 \a3/data_reg[62]  ( .D(\a3/N492 ), .CLK(clock), .Q(data_tan[62]) );
  DFFX1 \a5/data_reg[62]  ( .D(\a5/N492 ), .CLK(clock), .Q(data_sec[62]) );
  DFFX1 \a4/data_reg[52]  ( .D(\a4/N488 ), .CLK(clock), .Q(data_csc[52]) );
  DFFX1 \a4/data_reg[53]  ( .D(\a4/N489 ), .CLK(clock), .Q(data_csc[53]) );
  DFFX1 \a4/data_reg[54]  ( .D(\a4/N490 ), .CLK(clock), .Q(data_csc[54]) );
  DFFX1 \a4/data_reg[55]  ( .D(\a4/N491 ), .CLK(clock), .Q(data_csc[55]) );
  DFFX1 \a4/data_reg[56]  ( .D(\a4/N491 ), .CLK(clock), .Q(data_csc[56]) );
  DFFX1 \a4/data_reg[57]  ( .D(\a4/N491 ), .CLK(clock), .Q(data_csc[57]) );
  DFFX1 \a4/data_reg[58]  ( .D(\a4/N491 ), .CLK(clock), .Q(data_csc[58]) );
  DFFX1 \a4/data_reg[59]  ( .D(\a4/N491 ), .CLK(clock), .Q(data_csc[59]) );
  DFFX1 \a4/data_reg[60]  ( .D(\a4/N491 ), .CLK(clock), .Q(data_csc[60]) );
  DFFX1 \a4/data_reg[61]  ( .D(\a4/N491 ), .CLK(clock), .Q(data_csc[61]) );
  DFFX1 \a1/data_reg[53]  ( .D(\a1/N488 ), .CLK(clock), .Q(data_sin[53]) );
  DFFX1 \a6/data_reg[40]  ( .D(\a6/N476 ), .CLK(clock), .Q(data_cot[40]) );
  DFFX1 \a6/data_reg[46]  ( .D(\a6/N482 ), .CLK(clock), .Q(data_cot[46]) );
  DFFX1 \a5/data_reg[10]  ( .D(\a5/N446 ), .CLK(clock), .Q(data_sec[10]) );
  DFFX1 \a5/data_reg[38]  ( .D(\a5/N474 ), .CLK(clock), .Q(data_sec[38]) );
  DFFX1 \a4/data_reg[1]  ( .D(\a4/N437 ), .CLK(clock), .Q(data_csc[1]) );
  DFFX1 \a3/data_reg[0]  ( .D(\a3/N436 ), .CLK(clock), .Q(data_tan[0]) );
  DFFX1 \a6/data_reg[14]  ( .D(\a6/N450 ), .CLK(clock), .Q(data_cot[14]) );
  DFFX1 \a6/data_reg[21]  ( .D(\a6/N457 ), .CLK(clock), .Q(data_cot[21]) );
  DFFX1 \a5/data_reg[36]  ( .D(\a5/N472 ), .CLK(clock), .Q(data_sec[36]) );
  DFFX1 \a4/data_reg[18]  ( .D(\a4/N454 ), .CLK(clock), .Q(data_csc[18]) );
  DFFX1 \a4/data_reg[20]  ( .D(\a4/N456 ), .CLK(clock), .Q(data_csc[20]) );
  DFFX1 \a6/data_reg[5]  ( .D(\a6/N441 ), .CLK(clock), .Q(data_cot[5]) );
  DFFX1 \a4/data_reg[42]  ( .D(\a4/N478 ), .CLK(clock), .Q(data_csc[42]) );
  DFFX1 \a3/data_reg[28]  ( .D(\a3/N464 ), .CLK(clock), .Q(data_tan[28]) );
  DFFX1 \a2/data_reg[17]  ( .D(\a2/N452 ), .CLK(clock), .Q(data_cos[17]) );
  DFFX1 \a2/data_reg[24]  ( .D(\a2/N459 ), .CLK(clock), .Q(data_cos[24]) );
  DFFX1 \a4/data_reg[37]  ( .D(\a4/N473 ), .CLK(clock), .Q(data_csc[37]) );
  DFFX1 \a3/data_reg[1]  ( .D(\a3/N437 ), .CLK(clock), .Q(data_tan[1]) );
  DFFX1 \a3/data_reg[37]  ( .D(\a3/N473 ), .CLK(clock), .Q(data_tan[37]) );
  DFFX1 \a1/data_reg[0]  ( .D(\a1/N435 ), .CLK(clock), .Q(data_sin[0]) );
  DFFX1 \a1/data_reg[3]  ( .D(\a1/N438 ), .CLK(clock), .Q(data_sin[3]) );
  DFFX1 \a1/data_reg[21]  ( .D(\a1/N456 ), .CLK(clock), .Q(data_sin[21]) );
  DFFX1 \a1/data_reg[39]  ( .D(\a1/N474 ), .CLK(clock), .Q(data_sin[39]) );
  DFFX1 \a4/data_reg[26]  ( .D(\a4/N462 ), .CLK(clock), .Q(data_csc[26]) );
  DFFX1 \a1/data_reg[19]  ( .D(\a1/N454 ), .CLK(clock), .Q(data_sin[19]) );
  DFFX1 \a1/data_reg[44]  ( .D(\a1/N479 ), .CLK(clock), .Q(data_sin[44]) );
  DFFX1 \a6/data_reg[55]  ( .D(\a6/N491 ), .CLK(clock), .Q(data_cot[55]) );
  DFFX1 \a6/data_reg[56]  ( .D(\a6/N491 ), .CLK(clock), .Q(data_cot[56]) );
  DFFX1 \a6/data_reg[57]  ( .D(\a6/N491 ), .CLK(clock), .Q(data_cot[57]) );
  DFFX1 \a6/data_reg[58]  ( .D(\a6/N491 ), .CLK(clock), .Q(data_cot[58]) );
  DFFX1 \a6/data_reg[59]  ( .D(\a6/N491 ), .CLK(clock), .Q(data_cot[59]) );
  DFFX1 \a6/data_reg[60]  ( .D(\a6/N491 ), .CLK(clock), .Q(data_cot[60]) );
  DFFX1 \a6/data_reg[61]  ( .D(\a6/N491 ), .CLK(clock), .Q(data_cot[61]) );
  DFFX1 \a1/data_reg[50]  ( .D(\a1/N485 ), .CLK(clock), .Q(data_sin[50]) );
  DFFX1 \a1/data_reg[51]  ( .D(\a1/N486 ), .CLK(clock), .Q(data_sin[51]) );
  DFFX1 \a6/data_reg[16]  ( .D(\a6/N452 ), .CLK(clock), .Q(data_cot[16]) );
  DFFX1 \a6/data_reg[25]  ( .D(\a6/N461 ), .CLK(clock), .Q(data_cot[25]) );
  DFFX1 \a3/data_reg[49]  ( .D(\a3/N485 ), .CLK(clock), .Q(data_tan[49]) );
  DFFX1 \a6/data_reg[3]  ( .D(\a6/N439 ), .CLK(clock), .Q(data_cot[3]) );
  DFFX1 \a5/data_reg[29]  ( .D(\a5/N465 ), .CLK(clock), .Q(data_sec[29]) );
  DFFX1 \a5/data_reg[32]  ( .D(\a5/N468 ), .CLK(clock), .Q(data_sec[32]) );
  DFFX1 \a3/data_reg[3]  ( .D(\a3/N439 ), .CLK(clock), .Q(data_tan[3]) );
  DFFX1 \a6/data_reg[12]  ( .D(\a6/N448 ), .CLK(clock), .Q(data_cot[12]) );
  DFFX1 \a5/data_reg[53]  ( .D(\a5/N489 ), .CLK(clock), .Q(data_sec[53]) );
  DFFX1 \a2/data_reg[53]  ( .D(\a2/N488 ), .CLK(clock), .Q(data_cos[53]) );
  DFFX1 \a1/data_reg[15]  ( .D(\a1/N450 ), .CLK(clock), .Q(data_sin[15]) );
  DFFX1 \a6/data_reg[34]  ( .D(\a6/N470 ), .CLK(clock), .Q(data_cot[34]) );
  DFFX1 \a6/data_reg[39]  ( .D(\a6/N475 ), .CLK(clock), .Q(data_cot[39]) );
  DFFX1 \a4/data_reg[14]  ( .D(\a4/N450 ), .CLK(clock), .Q(data_csc[14]) );
  DFFX1 \a4/data_reg[41]  ( .D(\a4/N477 ), .CLK(clock), .Q(data_csc[41]) );
  DFFX1 \a3/data_reg[31]  ( .D(\a3/N467 ), .CLK(clock), .Q(data_tan[31]) );
  DFFX1 \a3/data_reg[40]  ( .D(\a3/N476 ), .CLK(clock), .Q(data_tan[40]) );
  DFFX1 \a1/data_reg[54]  ( .D(\a1/N489 ), .CLK(clock), .Q(data_sin[54]) );
  DFFX1 \a2/data_reg[54]  ( .D(\a2/N489 ), .CLK(clock), .Q(data_cos[54]) );
  DFFX1 \a1/data_reg[9]  ( .D(\a1/N444 ), .CLK(clock), .Q(data_sin[9]) );
  DFFX1 \a6/data_reg[19]  ( .D(\a6/N455 ), .CLK(clock), .Q(data_cot[19]) );
  DFFX1 \a5/data_reg[17]  ( .D(\a5/N453 ), .CLK(clock), .Q(data_sec[17]) );
  DFFX1 \a5/data_reg[28]  ( .D(\a5/N464 ), .CLK(clock), .Q(data_sec[28]) );
  DFFX1 \a4/data_reg[17]  ( .D(\a4/N453 ), .CLK(clock), .Q(data_csc[17]) );
  DFFX1 \a4/data_reg[47]  ( .D(\a4/N483 ), .CLK(clock), .Q(data_csc[47]) );
  DFFX1 \a3/data_reg[6]  ( .D(\a3/N442 ), .CLK(clock), .Q(data_tan[6]) );
  DFFX1 \a5/data_reg[7]  ( .D(\a5/N443 ), .CLK(clock), .Q(data_sec[7]) );
  DFFX1 \a6/data_reg[50]  ( .D(\a6/N486 ), .CLK(clock), .Q(data_cot[50]) );
  DFFX1 \a5/data_reg[45]  ( .D(\a5/N481 ), .CLK(clock), .Q(data_sec[45]) );
  DFFX1 \a3/data_reg[18]  ( .D(\a3/N454 ), .CLK(clock), .Q(data_tan[18]) );
  DFFX1 \a2/data_reg[18]  ( .D(\a2/N453 ), .CLK(clock), .Q(data_cos[18]) );
  DFFX1 \a5/data_reg[46]  ( .D(\a5/N482 ), .CLK(clock), .Q(data_sec[46]) );
  DFFX1 \a4/data_reg[2]  ( .D(\a4/N438 ), .CLK(clock), .Q(data_csc[2]) );
  DFFX1 \a1/data_reg[35]  ( .D(\a1/N470 ), .CLK(clock), .Q(data_sin[35]) );
  DFFX1 \a1/data_reg[43]  ( .D(\a1/N478 ), .CLK(clock), .Q(data_sin[43]) );
  DFFX1 \a1/data_reg[55]  ( .D(\a1/N490 ), .CLK(clock), .Q(data_sin[55]) );
  DFFX1 \a1/data_reg[56]  ( .D(\a1/N490 ), .CLK(clock), .Q(data_sin[56]) );
  DFFX1 \a1/data_reg[57]  ( .D(\a1/N490 ), .CLK(clock), .Q(data_sin[57]) );
  DFFX1 \a1/data_reg[58]  ( .D(\a1/N490 ), .CLK(clock), .Q(data_sin[58]) );
  DFFX1 \a1/data_reg[59]  ( .D(\a1/N490 ), .CLK(clock), .Q(data_sin[59]) );
  DFFX1 \a1/data_reg[60]  ( .D(\a1/N490 ), .CLK(clock), .Q(data_sin[60]) );
  DFFX1 \a1/data_reg[61]  ( .D(\a1/N490 ), .CLK(clock), .Q(data_sin[61]) );
  DFFX1 \a3/data_reg[63]  ( .D(\a3/N493 ), .CLK(clock), .Q(data_tan[63]) );
  DFFX1 \a6/data_reg[63]  ( .D(\a3/N493 ), .CLK(clock), .Q(data_cot[63]) );
  DFFX1 \quad_reg[1]  ( .D(N357), .CLK(clock), .Q(quad[1]) );
  DFFX1 \a2/data_reg[63]  ( .D(\a2/N491 ), .CLK(clock), .Q(data_cos[63]) );
  DFFX1 \a5/data_reg[63]  ( .D(\a2/N491 ), .CLK(clock), .Q(data_sec[63]) );
  DFFX1 \a1/data_reg[63]  ( .D(\a1/N491 ), .CLK(clock), .Q(data_sin[63]) );
  DFFX1 \a4/data_reg[63]  ( .D(\a1/N491 ), .CLK(clock), .Q(data_csc[63]) );
  INVX0 U5034 ( .INP(n4562), .ZN(n4557) );
  INVX0 U5035 ( .INP(n4557), .ZN(n4558) );
  INVX0 U5036 ( .INP(n4557), .ZN(n4559) );
  INVX0 U5037 ( .INP(n4557), .ZN(n4560) );
  INVX0 U5038 ( .INP(n4557), .ZN(n4561) );
  NOR3X0 U5039 ( .IN1(actv[2]), .IN2(actv[0]), .IN3(n9225), .QN(n4562) );
  NOR4X0 U5040 ( .IN1(divider_out[6]), .IN2(divider_out[7]), .IN3(
        divider_out[5]), .IN4(divider_out[4]), .QN(n4563) );
  INVX0 U5041 ( .INP(n4563), .ZN(n4566) );
  NAND3X0 U5042 ( .IN1(divider_out[1]), .IN2(divider_out[3]), .IN3(
        divider_out[2]), .QN(n4564) );
  NAND2X0 U5043 ( .IN1(n4564), .IN2(n4563), .QN(n4565) );
  AND2X1 U5044 ( .IN1(divider_out[8]), .IN2(n4565), .Q(n4581) );
  OA21X1 U5045 ( .IN1(divider_out[0]), .IN2(n4566), .IN3(n4581), .Q(n4666) );
  INVX0 U5046 ( .INP(degrees[22]), .ZN(n4859) );
  INVX0 U5047 ( .INP(degrees[21]), .ZN(n4876) );
  INVX0 U5048 ( .INP(degrees[20]), .ZN(n4896) );
  INVX0 U5049 ( .INP(degrees[18]), .ZN(n4952) );
  NAND4X0 U5050 ( .IN1(n4859), .IN2(n4876), .IN3(n4896), .IN4(n4952), .QN(
        n4569) );
  INVX0 U5051 ( .INP(degrees[28]), .ZN(n4792) );
  INVX0 U5052 ( .INP(degrees[26]), .ZN(n4789) );
  INVX0 U5053 ( .INP(degrees[25]), .ZN(n4802) );
  INVX0 U5054 ( .INP(degrees[19]), .ZN(n4921) );
  NAND4X0 U5055 ( .IN1(n4792), .IN2(n4789), .IN3(n4802), .IN4(n4921), .QN(
        n4568) );
  INVX0 U5056 ( .INP(degrees[12]), .ZN(n5058) );
  INVX0 U5057 ( .INP(degrees[23]), .ZN(n4835) );
  INVX0 U5058 ( .INP(degrees[11]), .ZN(n5086) );
  INVX0 U5059 ( .INP(degrees[10]), .ZN(n5101) );
  NAND4X0 U5060 ( .IN1(n5058), .IN2(n4835), .IN3(n5086), .IN4(n5101), .QN(
        n4567) );
  NOR3X0 U5061 ( .IN1(n4569), .IN2(n4568), .IN3(n4567), .QN(n4570) );
  INVX0 U5062 ( .INP(degrees[24]), .ZN(n4816) );
  INVX0 U5063 ( .INP(degrees[27]), .ZN(n4787) );
  INVX0 U5064 ( .INP(degrees[9]), .ZN(n5126) );
  NAND4X0 U5065 ( .IN1(n4570), .IN2(n4816), .IN3(n4787), .IN4(n5126), .QN(
        n4573) );
  NOR4X0 U5066 ( .IN1(degrees[14]), .IN2(degrees[31]), .IN3(degrees[29]), 
        .IN4(degrees[30]), .QN(n4571) );
  INVX0 U5067 ( .INP(degrees[17]), .ZN(n4963) );
  INVX0 U5068 ( .INP(degrees[16]), .ZN(n4977) );
  NAND3X0 U5069 ( .IN1(n4571), .IN2(n4963), .IN3(n4977), .QN(n4572) );
  NOR2X0 U5070 ( .IN1(n4573), .IN2(n4572), .QN(n4574) );
  INVX0 U5071 ( .INP(degrees[15]), .ZN(n5000) );
  INVX0 U5072 ( .INP(degrees[13]), .ZN(n5051) );
  NAND3X0 U5073 ( .IN1(n4574), .IN2(n5000), .IN3(n5051), .QN(n4607) );
  INVX0 U5074 ( .INP(degrees[7]), .ZN(n5244) );
  INVX0 U5075 ( .INP(degrees[4]), .ZN(n5218) );
  INVX0 U5076 ( .INP(\a7/N2 ), .ZN(n5330) );
  NAND3X0 U5077 ( .IN1(n5244), .IN2(n5218), .IN3(n5330), .QN(n4608) );
  NOR2X0 U5078 ( .IN1(\a7/N1 ), .IN2(\a7/N0 ), .QN(n4605) );
  INVX0 U5079 ( .INP(n4605), .ZN(n4609) );
  INVX0 U5080 ( .INP(degrees[8]), .ZN(n5139) );
  INVX0 U5081 ( .INP(degrees[6]), .ZN(n5251) );
  INVX0 U5082 ( .INP(degrees[5]), .ZN(n5256) );
  OA21X1 U5083 ( .IN1(n5251), .IN2(n5256), .IN3(n5244), .Q(n4587) );
  INVX0 U5084 ( .INP(degrees[3]), .ZN(n5247) );
  AND3X1 U5085 ( .IN1(n5244), .IN2(n5218), .IN3(n5247), .Q(n4575) );
  NOR3X0 U5086 ( .IN1(n5139), .IN2(n4587), .IN3(n4575), .QN(n4610) );
  OA21X1 U5087 ( .IN1(n4608), .IN2(n4609), .IN3(n4610), .Q(n4576) );
  OR2X1 U5088 ( .IN1(n4607), .IN2(n4576), .Q(n5308) );
  AND2X1 U5089 ( .IN1(n4666), .IN2(n5308), .Q(n9218) );
  NAND3X0 U5090 ( .IN1(divider_out[7]), .IN2(divider_out[5]), .IN3(
        divider_out[4]), .QN(n4594) );
  NOR2X0 U5091 ( .IN1(divider_out[3]), .IN2(divider_out[2]), .QN(n4577) );
  OA21X1 U5092 ( .IN1(n4594), .IN2(n4577), .IN3(n9444), .Q(n4592) );
  NOR4X0 U5093 ( .IN1(divider_out[1]), .IN2(divider_out[3]), .IN3(
        divider_out[0]), .IN4(divider_out[8]), .QN(n4578) );
  NOR2X0 U5094 ( .IN1(n4592), .IN2(n4578), .QN(n4584) );
  NAND2X0 U5095 ( .IN1(divider_out[7]), .IN2(divider_out[6]), .QN(n4593) );
  INVX0 U5096 ( .INP(n4593), .ZN(n4583) );
  NOR3X0 U5097 ( .IN1(divider_out[7]), .IN2(divider_out[5]), .IN3(
        divider_out[4]), .QN(n4579) );
  NOR2X0 U5098 ( .IN1(divider_out[6]), .IN2(divider_out[0]), .QN(n4598) );
  NAND2X0 U5099 ( .IN1(n4579), .IN2(n4598), .QN(n4580) );
  NAND2X0 U5100 ( .IN1(n4581), .IN2(n4580), .QN(n4582) );
  OA21X1 U5101 ( .IN1(n4584), .IN2(n4583), .IN3(n4582), .Q(n4667) );
  AND2X1 U5102 ( .IN1(n4667), .IN2(n5308), .Q(n4616) );
  NOR2X0 U5103 ( .IN1(n9218), .IN2(n4616), .QN(n4635) );
  INVX0 U5104 ( .INP(n4635), .ZN(n5295) );
  AND2X1 U5105 ( .IN1(divider_out[8]), .IN2(n5295), .Q(n5275) );
  INVX0 U5106 ( .INP(n9218), .ZN(n5274) );
  NOR2X0 U5107 ( .IN1(degrees[8]), .IN2(n4607), .QN(n4606) );
  NAND2X0 U5108 ( .IN1(n5247), .IN2(n5330), .QN(n5253) );
  NAND3X0 U5109 ( .IN1(degrees[4]), .IN2(degrees[5]), .IN3(n5253), .QN(n5257)
         );
  NAND2X0 U5110 ( .IN1(n5251), .IN2(n5257), .QN(n5245) );
  NAND2X0 U5111 ( .IN1(degrees[7]), .IN2(n5245), .QN(n4585) );
  NAND2X0 U5112 ( .IN1(n4606), .IN2(n4585), .QN(n4613) );
  OA221X1 U5113 ( .IN1(\a7/N2 ), .IN2(\a7/N1 ), .IN3(\a7/N2 ), .IN4(\a7/N0 ), 
        .IN5(degrees[3]), .Q(n4586) );
  NAND3X0 U5114 ( .IN1(n4586), .IN2(degrees[6]), .IN3(degrees[4]), .QN(n4588)
         );
  NAND2X0 U5115 ( .IN1(n4588), .IN2(n4587), .QN(n5306) );
  INVX0 U5116 ( .INP(n5306), .ZN(n5331) );
  NOR2X0 U5117 ( .IN1(n4613), .IN2(n5331), .QN(n9216) );
  INVX0 U5118 ( .INP(n9216), .ZN(n4615) );
  INVX0 U5119 ( .INP(n5308), .ZN(n4743) );
  OA221X1 U5120 ( .IN1(divider_out[2]), .IN2(divider_out[1]), .IN3(
        divider_out[2]), .IN4(divider_out[0]), .IN5(divider_out[3]), .Q(n4589)
         );
  OA221X1 U5121 ( .IN1(divider_out[5]), .IN2(divider_out[4]), .IN3(
        divider_out[5]), .IN4(n4589), .IN5(divider_out[6]), .Q(n4590) );
  NOR2X0 U5122 ( .IN1(divider_out[7]), .IN2(n4590), .QN(n4591) );
  NAND2X0 U5123 ( .IN1(n4591), .IN2(n9444), .QN(n5307) );
  NAND3X0 U5124 ( .IN1(n4593), .IN2(n5307), .IN3(n4592), .QN(n4668) );
  OR2X1 U5125 ( .IN1(n4743), .IN2(n4668), .Q(n4600) );
  NAND2X0 U5126 ( .IN1(divider_out[2]), .IN2(n5308), .QN(n5332) );
  NOR2X0 U5127 ( .IN1(n4594), .IN2(n5332), .QN(n4596) );
  NOR2X0 U5128 ( .IN1(divider_out[3]), .IN2(divider_out[1]), .QN(n4595) );
  AND3X1 U5129 ( .IN1(n4596), .IN2(n9444), .IN3(n4595), .Q(n4597) );
  NAND2X0 U5130 ( .IN1(n4598), .IN2(n4597), .QN(n4599) );
  NAND2X0 U5131 ( .IN1(n4600), .IN2(n4599), .QN(n9217) );
  INVX0 U5132 ( .INP(n9217), .ZN(n4614) );
  AO21X1 U5133 ( .IN1(degrees_tmp1[1]), .IN2(degrees_tmp1[0]), .IN3(
        degrees_tmp1[2]), .Q(n4601) );
  AND4X1 U5134 ( .IN1(degrees_tmp1[3]), .IN2(degrees_tmp1[6]), .IN3(
        degrees_tmp1[4]), .IN4(n4601), .Q(n4602) );
  NOR2X0 U5135 ( .IN1(n4602), .IN2(degrees_tmp1[7]), .QN(n4604) );
  NAND2X0 U5136 ( .IN1(degrees_tmp1[6]), .IN2(degrees_tmp1[5]), .QN(n4603) );
  AND2X1 U5137 ( .IN1(n4604), .IN2(n4603), .Q(n5280) );
  NAND4X0 U5138 ( .IN1(n4606), .IN2(n4605), .IN3(n5251), .IN4(n5247), .QN(
        n4612) );
  AOI221X1 U5139 ( .IN1(n4610), .IN2(n4609), .IN3(n4610), .IN4(n4608), .IN5(
        n4607), .QN(n4611) );
  AND3X1 U5140 ( .IN1(n4613), .IN2(n4612), .IN3(n4611), .Q(n5281) );
  INVX0 U5141 ( .INP(n5281), .ZN(n4745) );
  OR2X1 U5142 ( .IN1(n5280), .IN2(n4745), .Q(n4617) );
  NAND3X0 U5143 ( .IN1(n4615), .IN2(n4614), .IN3(n4617), .QN(n4631) );
  AO21X1 U5144 ( .IN1(divider_out[7]), .IN2(n5295), .IN3(n4631), .Q(n5272) );
  INVX0 U5145 ( .INP(n4616), .ZN(n4627) );
  NAND2X0 U5146 ( .IN1(divider_out[7]), .IN2(n9217), .QN(n4620) );
  INVX0 U5147 ( .INP(n4617), .ZN(n9215) );
  NAND2X0 U5148 ( .IN1(n9215), .IN2(degrees_tmp1[7]), .QN(n4619) );
  NAND2X0 U5149 ( .IN1(degrees[7]), .IN2(n9216), .QN(n4618) );
  AND4X1 U5150 ( .IN1(n4627), .IN2(n4620), .IN3(n4619), .IN4(n4618), .Q(n5271)
         );
  NOR2X0 U5151 ( .IN1(n4635), .IN2(n9443), .QN(n5278) );
  AOI222X1 U5152 ( .IN1(n9217), .IN2(divider_out[6]), .IN3(n9216), .IN4(
        degrees[6]), .IN5(degrees_tmp1[6]), .IN6(n9215), .QN(n5277) );
  AO21X1 U5153 ( .IN1(divider_out[5]), .IN2(n5295), .IN3(n4631), .Q(n5304) );
  NAND2X0 U5154 ( .IN1(divider_out[5]), .IN2(n9217), .QN(n4623) );
  NAND2X0 U5155 ( .IN1(degrees_tmp1[5]), .IN2(n9215), .QN(n4622) );
  NAND2X0 U5156 ( .IN1(degrees[5]), .IN2(n9216), .QN(n4621) );
  AND4X1 U5157 ( .IN1(n4627), .IN2(n4623), .IN3(n4622), .IN4(n4621), .Q(n5303)
         );
  AO21X1 U5158 ( .IN1(divider_out[4]), .IN2(n5295), .IN3(n4631), .Q(n5316) );
  NAND2X0 U5159 ( .IN1(divider_out[4]), .IN2(n9217), .QN(n4626) );
  NAND2X0 U5160 ( .IN1(n9215), .IN2(degrees_tmp1[4]), .QN(n4625) );
  NAND2X0 U5161 ( .IN1(degrees[4]), .IN2(n9216), .QN(n4624) );
  AND4X1 U5162 ( .IN1(n4627), .IN2(n4626), .IN3(n4625), .IN4(n4624), .Q(n5315)
         );
  AND2X1 U5163 ( .IN1(divider_out[3]), .IN2(n5295), .Q(n5288) );
  NAND2X0 U5164 ( .IN1(divider_out[3]), .IN2(n9217), .QN(n4630) );
  NAND2X0 U5165 ( .IN1(n9215), .IN2(degrees_tmp1[3]), .QN(n4629) );
  NAND2X0 U5166 ( .IN1(degrees[3]), .IN2(n9216), .QN(n4628) );
  AND4X1 U5167 ( .IN1(n5274), .IN2(n4630), .IN3(n4629), .IN4(n4628), .Q(n5287)
         );
  AO21X1 U5168 ( .IN1(divider_out[2]), .IN2(n5295), .IN3(n4631), .Q(n5326) );
  NAND2X0 U5169 ( .IN1(n9215), .IN2(degrees_tmp1[2]), .QN(n4634) );
  NAND2X0 U5170 ( .IN1(divider_out[2]), .IN2(n9217), .QN(n4633) );
  NAND2X0 U5171 ( .IN1(\a7/N2 ), .IN2(n9216), .QN(n4632) );
  AND4X1 U5172 ( .IN1(n4635), .IN2(n4634), .IN3(n4633), .IN4(n4632), .Q(n5325)
         );
  AND2X1 U5173 ( .IN1(divider_out[1]), .IN2(n5295), .Q(n4670) );
  NAND2X0 U5174 ( .IN1(divider_out[1]), .IN2(n9217), .QN(n4638) );
  NAND2X0 U5175 ( .IN1(n9215), .IN2(degrees_tmp1[1]), .QN(n4637) );
  NAND2X0 U5176 ( .IN1(\a7/N1 ), .IN2(n9216), .QN(n4636) );
  AND4X1 U5177 ( .IN1(n5274), .IN2(n4638), .IN3(n4637), .IN4(n4636), .Q(n4669)
         );
  AOI222X1 U5178 ( .IN1(n9217), .IN2(divider_out[0]), .IN3(n9216), .IN4(
        \a7/N0 ), .IN5(n9215), .IN6(degrees_tmp1[0]), .QN(n5296) );
  OR4X1 U5179 ( .IN1(degrees_tmp2[25]), .IN2(degrees_tmp2[18]), .IN3(
        degrees_tmp2[20]), .IN4(degrees_tmp2[22]), .Q(n4645) );
  OR4X1 U5180 ( .IN1(degrees_tmp2[17]), .IN2(degrees_tmp2[19]), .IN3(
        degrees_tmp2[27]), .IN4(degrees_tmp2[26]), .Q(n4644) );
  NOR4X0 U5181 ( .IN1(degrees_tmp2[7]), .IN2(degrees_tmp2[14]), .IN3(
        degrees_tmp2[29]), .IN4(degrees_tmp2[15]), .QN(n4642) );
  NOR4X0 U5182 ( .IN1(degrees_tmp2[28]), .IN2(degrees_tmp2[24]), .IN3(
        degrees_tmp2[30]), .IN4(degrees_tmp2[8]), .QN(n4641) );
  NOR4X0 U5183 ( .IN1(degrees_tmp2[13]), .IN2(degrees_tmp2[10]), .IN3(
        degrees_tmp2[21]), .IN4(degrees_tmp2[23]), .QN(n4640) );
  NOR4X0 U5184 ( .IN1(degrees_tmp2[11]), .IN2(degrees_tmp2[16]), .IN3(
        degrees_tmp2[12]), .IN4(degrees_tmp2[9]), .QN(n4639) );
  NAND4X0 U5185 ( .IN1(n4642), .IN2(n4641), .IN3(n4640), .IN4(n4639), .QN(
        n4643) );
  NOR4X0 U5186 ( .IN1(degrees_tmp2[31]), .IN2(n4645), .IN3(n4644), .IN4(n4643), 
        .QN(n5986) );
  NAND2X0 U5187 ( .IN1(n5986), .IN2(n9441), .QN(n6651) );
  INVX0 U5188 ( .INP(n6651), .ZN(n8220) );
  NAND2X0 U5189 ( .IN1(degrees_tmp2[3]), .IN2(degrees_tmp2[5]), .QN(n6921) );
  INVX0 U5190 ( .INP(n6921), .ZN(n5657) );
  NAND2X0 U5191 ( .IN1(n9436), .IN2(n9442), .QN(n9181) );
  INVX0 U5192 ( .INP(n9181), .ZN(n9080) );
  NOR2X0 U5193 ( .IN1(n9080), .IN2(n9440), .QN(n7956) );
  NAND4X0 U5194 ( .IN1(degrees_tmp2[2]), .IN2(n8220), .IN3(n5657), .IN4(n7956), 
        .QN(n8214) );
  NOR2X0 U5195 ( .IN1(degrees_tmp2[5]), .IN2(n9441), .QN(n8119) );
  NAND2X0 U5196 ( .IN1(n5986), .IN2(n8119), .QN(n8386) );
  INVX0 U5197 ( .INP(n8386), .ZN(n9047) );
  NAND2X0 U5198 ( .IN1(degrees_tmp2[3]), .IN2(n9434), .QN(n9060) );
  INVX0 U5199 ( .INP(n9060), .ZN(n8754) );
  NOR2X0 U5200 ( .IN1(n9436), .IN2(n9442), .QN(n8816) );
  NOR2X0 U5201 ( .IN1(degrees_tmp2[2]), .IN2(n8816), .QN(n6342) );
  INVX0 U5202 ( .INP(n6342), .ZN(n6797) );
  NAND2X0 U5203 ( .IN1(n8754), .IN2(n6797), .QN(n5786) );
  NAND2X0 U5204 ( .IN1(n9047), .IN2(n5786), .QN(n6234) );
  NAND2X0 U5205 ( .IN1(n8214), .IN2(n6234), .QN(\a5/N492 ) );
  NAND2X0 U5206 ( .IN1(n8119), .IN2(n9440), .QN(n5538) );
  INVX0 U5207 ( .INP(n5538), .ZN(n5937) );
  NAND2X0 U5208 ( .IN1(n5986), .IN2(n5937), .QN(n8268) );
  NAND2X0 U5209 ( .IN1(n9047), .IN2(n9060), .QN(n8422) );
  AO21X1 U5210 ( .IN1(n8268), .IN2(n6797), .IN3(n8422), .Q(n5783) );
  NAND2X0 U5211 ( .IN1(n6651), .IN2(n5783), .QN(\a2/N489 ) );
  NOR2X0 U5212 ( .IN1(degrees_tmp2[3]), .IN2(n9435), .QN(n8188) );
  NAND2X0 U5213 ( .IN1(n8188), .IN2(n9440), .QN(n6013) );
  INVX0 U5214 ( .INP(n6013), .ZN(n8242) );
  NAND2X0 U5215 ( .IN1(n9438), .IN2(n9436), .QN(n5588) );
  INVX0 U5216 ( .INP(n5588), .ZN(n5965) );
  NAND2X0 U5217 ( .IN1(n5965), .IN2(n9445), .QN(n7466) );
  INVX0 U5218 ( .INP(n7466), .ZN(n5863) );
  NAND2X0 U5219 ( .IN1(n8242), .IN2(n5863), .QN(n8212) );
  NAND2X0 U5220 ( .IN1(n8220), .IN2(n8212), .QN(n4646) );
  NAND2X0 U5221 ( .IN1(degrees_tmp2[3]), .IN2(n9435), .QN(n8595) );
  INVX0 U5222 ( .INP(n8595), .ZN(n7656) );
  NAND2X0 U5223 ( .IN1(n9445), .IN2(n9436), .QN(n8073) );
  INVX0 U5224 ( .INP(n5986), .ZN(n8213) );
  NOR2X0 U5225 ( .IN1(degrees_tmp2[5]), .IN2(n9440), .QN(n6710) );
  INVX0 U5226 ( .INP(n6710), .ZN(n7252) );
  NOR2X0 U5227 ( .IN1(n8213), .IN2(n7252), .QN(n5750) );
  INVX0 U5228 ( .INP(n5750), .ZN(n6893) );
  NOR2X0 U5229 ( .IN1(n8073), .IN2(n6893), .QN(n7582) );
  NAND2X0 U5230 ( .IN1(n7656), .IN2(n7582), .QN(n4675) );
  NAND2X0 U5231 ( .IN1(n4646), .IN2(n4675), .QN(\a3/N491 ) );
  NOR2X0 U5232 ( .IN1(n9437), .IN2(n9438), .QN(n4717) );
  INVX0 U5233 ( .INP(n4717), .ZN(n5355) );
  NOR2X0 U5234 ( .IN1(n8213), .IN2(n5355), .QN(n9105) );
  INVX0 U5235 ( .INP(n9105), .ZN(n9213) );
  NAND2X0 U5236 ( .IN1(n5986), .IN2(n9438), .QN(n8190) );
  NOR2X0 U5237 ( .IN1(degrees_tmp2[2]), .IN2(n9440), .QN(n8511) );
  INVX0 U5238 ( .INP(n8511), .ZN(n8909) );
  NOR2X0 U5239 ( .IN1(n8190), .IN2(n8909), .QN(n6173) );
  NAND2X0 U5240 ( .IN1(degrees_tmp2[3]), .IN2(n6173), .QN(n4763) );
  NOR2X0 U5241 ( .IN1(degrees_tmp2[0]), .IN2(n9442), .QN(n8760) );
  NAND2X0 U5242 ( .IN1(degrees_tmp2[0]), .IN2(n9442), .QN(n8282) );
  NOR2X0 U5243 ( .IN1(n8760), .IN2(n8728), .QN(n8727) );
  NOR2X0 U5244 ( .IN1(degrees_tmp2[3]), .IN2(n9434), .QN(n8572) );
  INVX0 U5245 ( .INP(n8572), .ZN(n8568) );
  NAND2X0 U5246 ( .IN1(n8220), .IN2(n8568), .QN(n6634) );
  OA21X1 U5247 ( .IN1(n4763), .IN2(n8727), .IN3(n6634), .Q(n4647) );
  NAND2X0 U5248 ( .IN1(n9213), .IN2(n4647), .QN(\a3/N490 ) );
  NAND2X0 U5249 ( .IN1(n8220), .IN2(n5965), .QN(n8937) );
  NOR2X0 U5250 ( .IN1(degrees_tmp2[2]), .IN2(n8937), .QN(n8074) );
  INVX0 U5251 ( .INP(n8268), .ZN(n8534) );
  NAND2X0 U5252 ( .IN1(n8534), .IN2(n9436), .QN(n8574) );
  NOR2X0 U5253 ( .IN1(n9445), .IN2(n8574), .QN(n6487) );
  NOR2X0 U5254 ( .IN1(n8074), .IN2(n6487), .QN(n4649) );
  NAND2X0 U5255 ( .IN1(n8595), .IN2(n8588), .QN(n4648) );
  NOR2X0 U5256 ( .IN1(n4649), .IN2(n4648), .QN(n4653) );
  NOR2X0 U5257 ( .IN1(n9437), .IN2(n9433), .QN(n6619) );
  NAND2X0 U5258 ( .IN1(n5986), .IN2(n6619), .QN(n7600) );
  NOR2X0 U5259 ( .IN1(n9445), .IN2(n9436), .QN(n6661) );
  NAND2X0 U5260 ( .IN1(n6661), .IN2(n9438), .QN(n5911) );
  NOR2X0 U5261 ( .IN1(n7600), .IN2(n5911), .QN(n8795) );
  INVX0 U5262 ( .INP(n8795), .ZN(n7480) );
  NAND2X0 U5263 ( .IN1(degrees_tmp2[2]), .IN2(n9438), .QN(n9132) );
  INVX0 U5264 ( .INP(n9132), .ZN(n8249) );
  NOR2X0 U5265 ( .IN1(n9435), .IN2(n8213), .QN(n5643) );
  NAND2X0 U5266 ( .IN1(n8249), .IN2(n5643), .QN(n7083) );
  INVX0 U5267 ( .INP(n7083), .ZN(n7214) );
  NAND2X0 U5268 ( .IN1(n8572), .IN2(n7214), .QN(n8840) );
  NAND2X0 U5269 ( .IN1(n9434), .IN2(n9441), .QN(n6401) );
  NOR2X0 U5270 ( .IN1(n8213), .IN2(n6401), .QN(n9190) );
  NAND2X0 U5271 ( .IN1(degrees_tmp2[2]), .IN2(n9190), .QN(n8124) );
  NAND2X0 U5272 ( .IN1(n9435), .IN2(n9438), .QN(n7402) );
  NOR2X0 U5273 ( .IN1(n8124), .IN2(n7402), .QN(n7653) );
  INVX0 U5274 ( .INP(n7653), .ZN(n8800) );
  NAND2X0 U5275 ( .IN1(n9080), .IN2(n9433), .QN(n8333) );
  INVX0 U5276 ( .INP(n8333), .ZN(n6207) );
  NAND2X0 U5277 ( .IN1(n9105), .IN2(n6207), .QN(n8592) );
  AND4X1 U5278 ( .IN1(n7480), .IN2(n8840), .IN3(n8800), .IN4(n8592), .Q(n4651)
         );
  NOR2X0 U5279 ( .IN1(degrees_tmp2[2]), .IN2(n8213), .QN(n8223) );
  INVX0 U5280 ( .INP(n8223), .ZN(n4700) );
  NOR2X0 U5281 ( .IN1(n4700), .IN2(n5538), .QN(n9074) );
  INVX0 U5282 ( .INP(n8816), .ZN(n9166) );
  NAND3X0 U5283 ( .IN1(n9074), .IN2(n9181), .IN3(n9166), .QN(n7331) );
  NAND2X0 U5284 ( .IN1(n9437), .IN2(n6173), .QN(n6308) );
  NAND2X0 U5285 ( .IN1(n8727), .IN2(n9433), .QN(n8123) );
  OA22X1 U5286 ( .IN1(n9433), .IN2(n7331), .IN3(n6308), .IN4(n8123), .Q(n4650)
         );
  NAND2X0 U5287 ( .IN1(n4717), .IN2(n9445), .QN(n5912) );
  NAND2X0 U5288 ( .IN1(n9434), .IN2(n5986), .QN(n4770) );
  NOR2X0 U5289 ( .IN1(n5912), .IN2(n4770), .QN(n6668) );
  NAND2X0 U5290 ( .IN1(n9433), .IN2(n9436), .QN(n8724) );
  NAND2X0 U5291 ( .IN1(n6668), .IN2(n8724), .QN(n7637) );
  NOR2X0 U5292 ( .IN1(n9438), .IN2(n9442), .QN(n8764) );
  INVX0 U5293 ( .INP(n8764), .ZN(n7717) );
  NAND2X0 U5294 ( .IN1(n9441), .IN2(n9436), .QN(n6049) );
  INVX0 U5295 ( .INP(n6049), .ZN(n6119) );
  NOR2X0 U5296 ( .IN1(n9434), .IN2(n8213), .QN(n5913) );
  NAND2X0 U5297 ( .IN1(n6119), .IN2(n5913), .QN(n6832) );
  NOR2X0 U5298 ( .IN1(n7717), .IN2(n6832), .QN(n7632) );
  NAND2X0 U5299 ( .IN1(degrees_tmp2[2]), .IN2(n7632), .QN(n6706) );
  NAND4X0 U5300 ( .IN1(n4651), .IN2(n4650), .IN3(n7637), .IN4(n6706), .QN(
        n4652) );
  NOR2X0 U5301 ( .IN1(n4653), .IN2(n4652), .QN(n4656) );
  NOR2X0 U5302 ( .IN1(n9434), .IN2(n9436), .QN(n7169) );
  NAND2X0 U5303 ( .IN1(n9435), .IN2(n9445), .QN(n9122) );
  NOR2X0 U5304 ( .IN1(n6651), .IN2(n9122), .QN(n8875) );
  INVX0 U5305 ( .INP(n8875), .ZN(n6337) );
  NOR2X0 U5306 ( .IN1(n9433), .IN2(n9445), .QN(n8699) );
  NAND2X0 U5307 ( .IN1(n5986), .IN2(n9435), .QN(n5758) );
  INVX0 U5308 ( .INP(n5758), .ZN(n5936) );
  NAND2X0 U5309 ( .IN1(n5936), .IN2(n9438), .QN(n8350) );
  INVX0 U5310 ( .INP(n8350), .ZN(n5553) );
  NAND2X0 U5311 ( .IN1(n8699), .IN2(n5553), .QN(n5651) );
  NOR2X0 U5312 ( .IN1(n9435), .IN2(n9213), .QN(n7093) );
  NAND2X0 U5313 ( .IN1(degrees_tmp2[3]), .IN2(n7093), .QN(n8761) );
  NAND2X0 U5314 ( .IN1(n8223), .IN2(n9441), .QN(n6510) );
  NOR2X0 U5315 ( .IN1(degrees_tmp2[3]), .IN2(n6510), .QN(n5423) );
  NAND2X0 U5316 ( .IN1(n5423), .IN2(n9438), .QN(n5975) );
  NAND4X0 U5317 ( .IN1(n6337), .IN2(n5651), .IN3(n8761), .IN4(n5975), .QN(
        n4654) );
  NAND2X0 U5318 ( .IN1(n7169), .IN2(n4654), .QN(n4655) );
  NAND2X0 U5319 ( .IN1(n4656), .IN2(n4655), .QN(\a2/N480 ) );
  NOR2X0 U5320 ( .IN1(n9434), .IN2(n9445), .QN(n7517) );
  NOR2X0 U5321 ( .IN1(degrees_tmp2[5]), .IN2(n7600), .QN(n6859) );
  NAND2X0 U5322 ( .IN1(n6859), .IN2(n9436), .QN(n8921) );
  NOR2X0 U5323 ( .IN1(n9433), .IN2(n8213), .QN(n5832) );
  INVX0 U5324 ( .INP(n5832), .ZN(n4755) );
  NOR2X0 U5325 ( .IN1(n4755), .IN2(n5538), .QN(n8408) );
  NAND2X0 U5326 ( .IN1(degrees_tmp2[2]), .IN2(n8408), .QN(n9127) );
  OA22X1 U5327 ( .IN1(n7517), .IN2(n8921), .IN3(n8727), .IN4(n9127), .Q(n4658)
         );
  NOR2X0 U5328 ( .IN1(n6049), .IN2(n5758), .QN(n8753) );
  NAND2X0 U5329 ( .IN1(n9433), .IN2(n8753), .QN(n9119) );
  INVX0 U5330 ( .INP(n9119), .ZN(n5352) );
  NOR2X0 U5331 ( .IN1(n9434), .IN2(n9438), .QN(n7437) );
  INVX0 U5332 ( .INP(n7437), .ZN(n7913) );
  NAND3X0 U5333 ( .IN1(degrees_tmp2[2]), .IN2(n5352), .IN3(n7913), .QN(n4657)
         );
  INVX0 U5334 ( .INP(n7600), .ZN(n9203) );
  NAND2X0 U5335 ( .IN1(n9445), .IN2(n9442), .QN(n7760) );
  NOR2X0 U5336 ( .IN1(n9440), .IN2(n7760), .QN(n7700) );
  NAND2X0 U5337 ( .IN1(n9203), .IN2(n7700), .QN(n8380) );
  NOR2X0 U5338 ( .IN1(n9437), .IN2(n5758), .QN(n5739) );
  NOR2X0 U5339 ( .IN1(n9433), .IN2(n8073), .QN(n5780) );
  NAND2X0 U5340 ( .IN1(n5739), .IN2(n5780), .QN(n7940) );
  NAND4X0 U5341 ( .IN1(n4658), .IN2(n4657), .IN3(n8380), .IN4(n7940), .QN(
        n4662) );
  NAND2X0 U5342 ( .IN1(n4717), .IN2(degrees_tmp2[0]), .QN(n4693) );
  INVX0 U5343 ( .INP(n4693), .ZN(n5545) );
  NAND2X0 U5344 ( .IN1(n5832), .IN2(n5545), .QN(n9098) );
  NAND2X0 U5345 ( .IN1(degrees_tmp2[2]), .IN2(n9434), .QN(n9032) );
  NOR2X0 U5346 ( .IN1(n9098), .IN2(n9032), .QN(n7333) );
  NAND2X0 U5347 ( .IN1(n9437), .IN2(n9433), .QN(n7552) );
  NOR2X0 U5348 ( .IN1(degrees_tmp2[5]), .IN2(n7552), .QN(n7050) );
  INVX0 U5349 ( .INP(n4770), .ZN(n8101) );
  NAND2X0 U5350 ( .IN1(n7050), .IN2(n8101), .QN(n8071) );
  INVX0 U5351 ( .INP(n8071), .ZN(n6100) );
  NOR2X0 U5352 ( .IN1(n7333), .IN2(n6100), .QN(n6819) );
  NOR2X0 U5353 ( .IN1(n9440), .IN2(n9436), .QN(n8995) );
  INVX0 U5354 ( .INP(n8995), .ZN(n8787) );
  INVX0 U5355 ( .INP(n8190), .ZN(n9210) );
  NOR2X0 U5356 ( .IN1(n8220), .IN2(n9210), .QN(n4728) );
  NOR2X0 U5357 ( .IN1(n9437), .IN2(n9445), .QN(n5472) );
  NOR2X0 U5358 ( .IN1(degrees_tmp2[2]), .IN2(n9441), .QN(n8022) );
  NOR2X0 U5359 ( .IN1(n5472), .IN2(n8022), .QN(n8510) );
  NOR2X0 U5360 ( .IN1(n4728), .IN2(n8510), .QN(n8354) );
  NAND2X0 U5361 ( .IN1(n8354), .IN2(n9442), .QN(n5615) );
  OA22X1 U5362 ( .IN1(n9080), .IN2(n6819), .IN3(n8787), .IN4(n5615), .Q(n4660)
         );
  NAND2X0 U5363 ( .IN1(n8223), .IN2(n9438), .QN(n5938) );
  NOR2X0 U5364 ( .IN1(n9437), .IN2(n5938), .QN(n7032) );
  NAND2X0 U5365 ( .IN1(degrees_tmp2[0]), .IN2(n9433), .QN(n9149) );
  INVX0 U5366 ( .INP(n9149), .ZN(n8883) );
  NOR2X0 U5367 ( .IN1(n8883), .IN2(n9440), .QN(n7012) );
  NAND2X0 U5368 ( .IN1(n7032), .IN2(n7012), .QN(n7944) );
  NOR2X0 U5369 ( .IN1(n9435), .IN2(n9433), .QN(n9073) );
  NOR2X0 U5370 ( .IN1(n4700), .IN2(n4693), .QN(n6449) );
  NAND2X0 U5371 ( .IN1(n9073), .IN2(n6449), .QN(n8043) );
  OR2X1 U5372 ( .IN1(n9434), .IN2(n9433), .Q(n6919) );
  INVX0 U5373 ( .INP(n6919), .ZN(n8675) );
  NAND2X0 U5374 ( .IN1(degrees_tmp2[0]), .IN2(n9438), .QN(n7920) );
  NOR2X0 U5375 ( .IN1(n5758), .IN2(n7920), .QN(n6016) );
  NAND2X0 U5376 ( .IN1(n8675), .IN2(n6016), .QN(n7981) );
  INVX0 U5377 ( .INP(n6619), .ZN(n7808) );
  NOR2X0 U5378 ( .IN1(n5758), .IN2(n7808), .QN(n5709) );
  NAND2X0 U5379 ( .IN1(n7517), .IN2(n5709), .QN(n6112) );
  NAND2X0 U5380 ( .IN1(n7981), .IN2(n6112), .QN(n8770) );
  NAND2X0 U5381 ( .IN1(n9132), .IN2(n8770), .QN(n4659) );
  NAND4X0 U5382 ( .IN1(n4660), .IN2(n7944), .IN3(n8043), .IN4(n4659), .QN(
        n4661) );
  NOR2X0 U5383 ( .IN1(n4662), .IN2(n4661), .QN(n4665) );
  NAND2X0 U5384 ( .IN1(n9047), .IN2(n6342), .QN(n9204) );
  NOR2X0 U5385 ( .IN1(n9435), .IN2(n9445), .QN(n8575) );
  INVX0 U5386 ( .INP(n8575), .ZN(n7745) );
  NOR2X0 U5387 ( .IN1(n9213), .IN2(n7745), .QN(n7654) );
  NAND2X0 U5388 ( .IN1(n7654), .IN2(n9436), .QN(n7326) );
  INVX0 U5389 ( .INP(n7920), .ZN(n8000) );
  NAND2X0 U5390 ( .IN1(n5986), .IN2(n8000), .QN(n6306) );
  NOR2X0 U5391 ( .IN1(degrees_tmp2[2]), .IN2(n6306), .QN(n6697) );
  NAND2X0 U5392 ( .IN1(n6697), .IN2(n9441), .QN(n8384) );
  NAND2X0 U5393 ( .IN1(n5643), .IN2(n9438), .QN(n6322) );
  NOR2X0 U5394 ( .IN1(n9437), .IN2(n6322), .QN(n8302) );
  NAND2X0 U5395 ( .IN1(degrees_tmp2[0]), .IN2(n8302), .QN(n8587) );
  NAND4X0 U5396 ( .IN1(n9204), .IN2(n7326), .IN3(n8384), .IN4(n8587), .QN(
        n4663) );
  NAND2X0 U5397 ( .IN1(n8572), .IN2(n4663), .QN(n4664) );
  NAND2X0 U5398 ( .IN1(n4665), .IN2(n4664), .QN(\a6/N478 ) );
  NAND3X0 U5399 ( .IN1(n5281), .IN2(n5280), .IN3(degrees_tmp1[1]), .QN(n4673)
         );
  NAND2X0 U5400 ( .IN1(n4743), .IN2(n4745), .QN(n5329) );
  NOR2X0 U5401 ( .IN1(n9216), .IN2(n5329), .QN(n5294) );
  NOR2X0 U5402 ( .IN1(n4667), .IN2(n4666), .QN(n4742) );
  NAND2X0 U5403 ( .IN1(n4742), .IN2(n4668), .QN(n5333) );
  NOR2X0 U5404 ( .IN1(n4743), .IN2(n5333), .QN(n5319) );
  FADDX1 U5405 ( .A(n4670), .B(n4669), .CI(n5296), .CO(n5324), .S(n4671) );
  AOI221X1 U5406 ( .IN1(\a7/N1 ), .IN2(n5294), .IN3(divider_out[1]), .IN4(
        n5319), .IN5(n4671), .QN(n4672) );
  NAND2X0 U5407 ( .IN1(n4673), .IN2(n4672), .QN(N325) );
  NAND4X0 U5408 ( .IN1(n9434), .IN2(degrees_tmp2[2]), .IN3(n5657), .IN4(n9181), 
        .QN(n4674) );
  NAND2X0 U5409 ( .IN1(n8220), .IN2(n4674), .QN(n8217) );
  NAND2X0 U5410 ( .IN1(n8217), .IN2(n4675), .QN(\a5/N491 ) );
  INVX0 U5411 ( .INP(n5938), .ZN(n6826) );
  NOR2X0 U5412 ( .IN1(n9434), .IN2(n8282), .QN(n7179) );
  NAND2X0 U5413 ( .IN1(n6826), .IN2(n7179), .QN(n7107) );
  INVX0 U5414 ( .INP(n7760), .ZN(n9082) );
  NAND3X0 U5415 ( .IN1(degrees_tmp2[3]), .IN2(n9047), .IN3(n9082), .QN(n8244)
         );
  NOR2X0 U5416 ( .IN1(degrees_tmp2[0]), .IN2(n9445), .QN(n8752) );
  OR2X1 U5417 ( .IN1(degrees_tmp2[3]), .IN2(n9442), .Q(n7736) );
  NOR2X0 U5418 ( .IN1(n9440), .IN2(n7736), .QN(n6017) );
  INVX0 U5419 ( .INP(n6017), .ZN(n7209) );
  NOR2X0 U5420 ( .IN1(n6651), .IN2(n7209), .QN(n7486) );
  NAND2X0 U5421 ( .IN1(n8752), .IN2(n7486), .QN(n6404) );
  NOR2X0 U5422 ( .IN1(n9434), .IN2(n9213), .QN(n5949) );
  NOR2X0 U5423 ( .IN1(n9435), .IN2(n8883), .QN(n5688) );
  NAND2X0 U5424 ( .IN1(n5949), .IN2(n5688), .QN(n7379) );
  NAND4X0 U5425 ( .IN1(n7107), .IN2(n8244), .IN3(n6404), .IN4(n7379), .QN(
        n4679) );
  NAND2X0 U5426 ( .IN1(degrees_tmp2[2]), .IN2(n9433), .QN(n9048) );
  INVX0 U5427 ( .INP(n9048), .ZN(n8825) );
  NAND2X0 U5428 ( .IN1(n8220), .IN2(n9440), .QN(n6069) );
  NOR2X0 U5429 ( .IN1(degrees_tmp2[5]), .IN2(n6069), .QN(n8181) );
  NAND2X0 U5430 ( .IN1(n8760), .IN2(n8181), .QN(n7060) );
  INVX0 U5431 ( .INP(n8022), .ZN(n8886) );
  NOR2X0 U5432 ( .IN1(n8190), .IN2(n8886), .QN(n6637) );
  INVX0 U5433 ( .INP(n6637), .ZN(n7534) );
  NOR2X0 U5434 ( .IN1(n9433), .IN2(n7534), .QN(n7421) );
  INVX0 U5435 ( .INP(n9073), .ZN(n7686) );
  NOR2X0 U5436 ( .IN1(n8386), .IN2(n7686), .QN(n7121) );
  NOR2X0 U5437 ( .IN1(n7421), .IN2(n7121), .QN(n6488) );
  INVX0 U5438 ( .INP(n7169), .ZN(n9061) );
  OA22X1 U5439 ( .IN1(n8825), .IN2(n7060), .IN3(n6488), .IN4(n9061), .Q(n4677)
         );
  NAND2X0 U5440 ( .IN1(n5986), .IN2(n7050), .QN(n6371) );
  INVX0 U5441 ( .INP(n6371), .ZN(n7936) );
  NAND2X0 U5442 ( .IN1(n7936), .IN2(n9436), .QN(n7011) );
  INVX0 U5443 ( .INP(n7517), .ZN(n8489) );
  NAND2X0 U5444 ( .IN1(n8489), .IN2(n8909), .QN(n9099) );
  NAND2X0 U5445 ( .IN1(n9435), .IN2(n8909), .QN(n6509) );
  NAND2X0 U5446 ( .IN1(n9099), .IN2(n6509), .QN(n7571) );
  NAND2X0 U5447 ( .IN1(degrees_tmp2[5]), .IN2(n5739), .QN(n8842) );
  INVX0 U5448 ( .INP(n8842), .ZN(n6261) );
  NOR2X0 U5449 ( .IN1(n9436), .IN2(n8568), .QN(n7389) );
  NAND2X0 U5450 ( .IN1(n6261), .IN2(n7389), .QN(n7662) );
  OA21X1 U5451 ( .IN1(n7011), .IN2(n7571), .IN3(n7662), .Q(n4676) );
  NOR2X0 U5452 ( .IN1(n9440), .IN2(n9442), .QN(n8424) );
  NOR2X0 U5453 ( .IN1(n8213), .IN2(n9436), .QN(n8301) );
  NAND2X0 U5454 ( .IN1(n6619), .IN2(n8301), .QN(n7746) );
  NOR2X0 U5455 ( .IN1(degrees_tmp2[2]), .IN2(n7746), .QN(n6584) );
  NAND2X0 U5456 ( .IN1(n8424), .IN2(n6584), .QN(n8584) );
  NAND2X0 U5457 ( .IN1(n9437), .IN2(degrees_tmp2[0]), .QN(n7298) );
  INVX0 U5458 ( .INP(n7298), .ZN(n6650) );
  NOR2X0 U5459 ( .IN1(degrees_tmp2[3]), .IN2(degrees_tmp2[5]), .QN(n8198) );
  INVX0 U5460 ( .INP(n8198), .ZN(n5757) );
  NOR2X0 U5461 ( .IN1(n5757), .IN2(n4770), .QN(n9202) );
  NAND2X0 U5462 ( .IN1(n6650), .IN2(n9202), .QN(n7025) );
  INVX0 U5463 ( .INP(n7025), .ZN(n8656) );
  NAND2X0 U5464 ( .IN1(n9435), .IN2(n8656), .QN(n8504) );
  NAND4X0 U5465 ( .IN1(n4677), .IN2(n4676), .IN3(n8584), .IN4(n8504), .QN(
        n4678) );
  NOR2X0 U5466 ( .IN1(n4679), .IN2(n4678), .QN(n4683) );
  INVX0 U5467 ( .INP(n8424), .ZN(n8822) );
  INVX0 U5468 ( .INP(n9190), .ZN(n7416) );
  NOR2X0 U5469 ( .IN1(n9438), .IN2(n7416), .QN(n9182) );
  NAND2X0 U5470 ( .IN1(n9182), .IN2(n8825), .QN(n9165) );
  NAND2X0 U5471 ( .IN1(n9105), .IN2(n5780), .QN(n8964) );
  INVX0 U5472 ( .INP(n6401), .ZN(n8940) );
  NAND2X0 U5473 ( .IN1(n8301), .IN2(n8940), .QN(n5803) );
  INVX0 U5474 ( .INP(n5803), .ZN(n5494) );
  NAND2X0 U5475 ( .IN1(degrees_tmp2[2]), .IN2(n5494), .QN(n6038) );
  INVX0 U5476 ( .INP(n8724), .ZN(n7784) );
  NOR2X0 U5477 ( .IN1(n9437), .IN2(n8190), .QN(n7699) );
  INVX0 U5478 ( .INP(n7699), .ZN(n6747) );
  NOR2X0 U5479 ( .IN1(n7784), .IN2(n6747), .QN(n8206) );
  NAND2X0 U5480 ( .IN1(n9434), .IN2(n8206), .QN(n4680) );
  NAND4X0 U5481 ( .IN1(n9165), .IN2(n8964), .IN3(n6038), .IN4(n4680), .QN(
        n4681) );
  NAND2X0 U5482 ( .IN1(n8822), .IN2(n4681), .QN(n4682) );
  NAND2X0 U5483 ( .IN1(n4683), .IN2(n4682), .QN(\a2/N451 ) );
  NAND2X0 U5484 ( .IN1(n8675), .IN2(n9438), .QN(n6369) );
  NOR2X0 U5485 ( .IN1(n4700), .IN2(n6369), .QN(n9076) );
  NAND2X0 U5486 ( .IN1(degrees_tmp2[0]), .IN2(n9076), .QN(n8651) );
  NAND2X0 U5487 ( .IN1(n5472), .IN2(n8301), .QN(n7291) );
  NOR2X0 U5488 ( .IN1(n7291), .IN2(n9060), .QN(n8179) );
  INVX0 U5489 ( .INP(n8179), .ZN(n7767) );
  NAND2X0 U5490 ( .IN1(n6710), .IN2(n9442), .QN(n6968) );
  NOR2X0 U5491 ( .IN1(n8213), .IN2(n6968), .QN(n6620) );
  INVX0 U5492 ( .INP(n6620), .ZN(n4779) );
  NOR2X0 U5493 ( .IN1(n4779), .IN2(n8886), .QN(n7984) );
  INVX0 U5494 ( .INP(n7984), .ZN(n9169) );
  INVX0 U5495 ( .INP(n8124), .ZN(n8485) );
  NAND2X0 U5496 ( .IN1(degrees_tmp2[5]), .IN2(n9442), .QN(n7706) );
  INVX0 U5497 ( .INP(n7706), .ZN(n7841) );
  NAND2X0 U5498 ( .IN1(n8485), .IN2(n7841), .QN(n9140) );
  NAND4X0 U5499 ( .IN1(n8651), .IN2(n7767), .IN3(n9169), .IN4(n9140), .QN(
        n4687) );
  INVX0 U5500 ( .INP(n8699), .ZN(n6198) );
  NAND2X0 U5501 ( .IN1(n9440), .IN2(n9436), .QN(n6836) );
  NOR2X0 U5502 ( .IN1(n6198), .IN2(n6836), .QN(n5872) );
  NAND2X0 U5503 ( .IN1(n9105), .IN2(n5872), .QN(n6814) );
  NAND2X0 U5504 ( .IN1(n9445), .IN2(n9440), .QN(n8474) );
  NOR2X0 U5505 ( .IN1(n7600), .IN2(n8474), .QN(n7921) );
  NAND2X0 U5506 ( .IN1(n9442), .IN2(n7921), .QN(n7096) );
  AND2X1 U5507 ( .IN1(n6814), .IN2(n7096), .Q(n7503) );
  NAND2X0 U5508 ( .IN1(n8760), .IN2(n9445), .QN(n8083) );
  INVX0 U5509 ( .INP(n8083), .ZN(n9209) );
  NAND3X0 U5510 ( .IN1(n8940), .IN2(n9210), .IN3(n9209), .QN(n7099) );
  NAND2X0 U5511 ( .IN1(n7517), .IN2(n9210), .QN(n8684) );
  NOR2X0 U5512 ( .IN1(n9442), .IN2(n8684), .QN(n7915) );
  NAND2X0 U5513 ( .IN1(n7915), .IN2(n9441), .QN(n7820) );
  NAND3X0 U5514 ( .IN1(degrees_tmp2[2]), .IN2(n5986), .IN3(n8119), .QN(n5624)
         );
  NAND2X0 U5515 ( .IN1(n9213), .IN2(n5624), .QN(n8954) );
  NAND2X0 U5516 ( .IN1(n9442), .IN2(n8954), .QN(n8400) );
  AO221X1 U5517 ( .IN1(n7820), .IN2(n6919), .IN3(n7820), .IN4(n8400), .IN5(
        n8883), .Q(n4685) );
  NOR2X0 U5518 ( .IN1(n9438), .IN2(n7600), .QN(n8529) );
  NAND2X0 U5519 ( .IN1(n9435), .IN2(n8529), .QN(n6311) );
  NOR2X0 U5520 ( .IN1(n9445), .IN2(n7736), .QN(n8240) );
  NAND2X0 U5521 ( .IN1(n9210), .IN2(n8240), .QN(n7293) );
  NAND2X0 U5522 ( .IN1(n6311), .IN2(n7293), .QN(n6686) );
  NAND2X0 U5523 ( .IN1(n8995), .IN2(n6686), .QN(n4684) );
  NAND4X0 U5524 ( .IN1(n7503), .IN2(n7099), .IN3(n4685), .IN4(n4684), .QN(
        n4686) );
  NOR2X0 U5525 ( .IN1(n4687), .IN2(n4686), .QN(n4691) );
  INVX0 U5526 ( .INP(n8474), .ZN(n8978) );
  NAND2X0 U5527 ( .IN1(n5986), .IN2(n6119), .QN(n6120) );
  NOR2X0 U5528 ( .IN1(n7717), .IN2(n6120), .QN(n8475) );
  NAND2X0 U5529 ( .IN1(n8978), .IN2(n8475), .QN(n6535) );
  INVX0 U5530 ( .INP(n6510), .ZN(n5766) );
  NAND2X0 U5531 ( .IN1(n9434), .IN2(n9080), .QN(n9046) );
  INVX0 U5532 ( .INP(n9046), .ZN(n6154) );
  NAND2X0 U5533 ( .IN1(n5766), .IN2(n6154), .QN(n8042) );
  NOR2X0 U5534 ( .IN1(n9435), .IN2(n8386), .QN(n5626) );
  INVX0 U5535 ( .INP(n5626), .ZN(n6887) );
  NOR2X0 U5536 ( .IN1(n7517), .IN2(n6887), .QN(n6438) );
  INVX0 U5537 ( .INP(n6438), .ZN(n4688) );
  NAND2X0 U5538 ( .IN1(n9434), .IN2(n4717), .QN(n5433) );
  NAND2X0 U5539 ( .IN1(n5538), .IN2(n5433), .QN(n8300) );
  NAND2X0 U5540 ( .IN1(n5986), .IN2(n8300), .QN(n8331) );
  INVX0 U5541 ( .INP(n8331), .ZN(n6698) );
  NAND2X0 U5542 ( .IN1(n8752), .IN2(n6698), .QN(n7444) );
  NAND4X0 U5543 ( .IN1(n6535), .IN2(n8042), .IN3(n4688), .IN4(n7444), .QN(
        n4689) );
  NAND2X0 U5544 ( .IN1(n9433), .IN2(n4689), .QN(n4690) );
  NAND2X0 U5545 ( .IN1(n4691), .IN2(n4690), .QN(\a4/N470 ) );
  NAND2X0 U5546 ( .IN1(degrees_tmp2[2]), .IN2(n5986), .QN(n5653) );
  INVX0 U5547 ( .INP(n5653), .ZN(n6493) );
  NAND2X0 U5548 ( .IN1(n5937), .IN2(n6493), .QN(n7510) );
  NOR2X0 U5549 ( .IN1(n8728), .IN2(n7510), .QN(n6929) );
  NAND2X0 U5550 ( .IN1(degrees_tmp2[2]), .IN2(n9435), .QN(n7233) );
  NOR2X0 U5551 ( .IN1(n5803), .IN2(n7233), .QN(n6914) );
  NOR2X0 U5552 ( .IN1(n6929), .IN2(n6914), .QN(n8915) );
  NAND2X0 U5553 ( .IN1(n9435), .IN2(n9440), .QN(n7945) );
  INVX0 U5554 ( .INP(n7945), .ZN(n9125) );
  NOR2X0 U5555 ( .IN1(n9435), .IN2(n9440), .QN(n8796) );
  NOR2X0 U5556 ( .IN1(n9125), .IN2(n8796), .QN(n9071) );
  INVX0 U5557 ( .INP(n9071), .ZN(n8171) );
  NAND2X0 U5558 ( .IN1(degrees_tmp2[2]), .IN2(n7945), .QN(n8938) );
  NAND2X0 U5559 ( .IN1(n8171), .IN2(n8938), .QN(n8227) );
  NOR2X0 U5560 ( .IN1(n6651), .IN2(n8227), .QN(n8395) );
  NOR2X0 U5561 ( .IN1(n8534), .IN2(n8395), .QN(n4692) );
  INVX0 U5562 ( .INP(n8760), .ZN(n8041) );
  OA22X1 U5563 ( .IN1(n4692), .IN2(n8724), .IN3(n8041), .IN4(n8422), .Q(n4694)
         );
  NAND2X0 U5564 ( .IN1(n6493), .IN2(n7050), .QN(n7394) );
  NOR2X0 U5565 ( .IN1(n8213), .IN2(n4693), .QN(n8567) );
  NAND2X0 U5566 ( .IN1(n8567), .IN2(n9071), .QN(n7988) );
  NAND4X0 U5567 ( .IN1(n8915), .IN2(n4694), .IN3(n7394), .IN4(n7988), .QN(
        n4696) );
  NAND2X0 U5568 ( .IN1(n9105), .IN2(n9436), .QN(n7679) );
  INVX0 U5569 ( .INP(n7679), .ZN(n8898) );
  NAND2X0 U5570 ( .IN1(n8898), .IN2(n8825), .QN(n8821) );
  NOR2X0 U5571 ( .IN1(degrees_tmp2[3]), .IN2(n8842), .QN(n8788) );
  NAND2X0 U5572 ( .IN1(n8788), .IN2(n9445), .QN(n5646) );
  INVX0 U5573 ( .INP(n5646), .ZN(n7832) );
  NAND2X0 U5574 ( .IN1(degrees_tmp2[0]), .IN2(n7832), .QN(n7459) );
  NAND2X0 U5575 ( .IN1(n7093), .IN2(n9445), .QN(n8564) );
  INVX0 U5576 ( .INP(n8564), .ZN(n8723) );
  NAND2X0 U5577 ( .IN1(n8675), .IN2(n8723), .QN(n5460) );
  NOR2X0 U5578 ( .IN1(n7600), .IN2(n7402), .QN(n5880) );
  NAND2X0 U5579 ( .IN1(n9434), .IN2(n9436), .QN(n8692) );
  NAND2X0 U5580 ( .IN1(n9061), .IN2(n8692), .QN(n8431) );
  NAND2X0 U5581 ( .IN1(n5880), .IN2(n8431), .QN(n8790) );
  NAND4X0 U5582 ( .IN1(n8821), .IN2(n7459), .IN3(n5460), .IN4(n8790), .QN(
        n4695) );
  NOR2X0 U5583 ( .IN1(n4696), .IN2(n4695), .QN(n4699) );
  INVX0 U5584 ( .INP(n6836), .ZN(n8467) );
  NOR2X0 U5585 ( .IN1(n8467), .IN2(n7686), .QN(n9104) );
  INVX0 U5586 ( .INP(n5472), .ZN(n6554) );
  NOR2X0 U5587 ( .IN1(n8213), .IN2(n6554), .QN(n6155) );
  INVX0 U5588 ( .INP(n6306), .ZN(n6613) );
  OA21X1 U5589 ( .IN1(n6155), .IN2(n6613), .IN3(n9132), .Q(n8241) );
  NAND2X0 U5590 ( .IN1(n9434), .IN2(n8241), .QN(n6361) );
  NAND2X0 U5591 ( .IN1(n7534), .IN2(n6361), .QN(n4697) );
  NAND2X0 U5592 ( .IN1(n9104), .IN2(n4697), .QN(n4698) );
  NAND2X0 U5593 ( .IN1(n4699), .IN2(n4698), .QN(\a1/N455 ) );
  INVX0 U5594 ( .INP(n6069), .ZN(n5419) );
  NAND2X0 U5595 ( .IN1(n5419), .IN2(n9433), .QN(n6606) );
  INVX0 U5596 ( .INP(n6606), .ZN(n6756) );
  INVX0 U5597 ( .INP(n8282), .ZN(n8728) );
  NAND2X0 U5598 ( .IN1(n8728), .IN2(n9445), .QN(n6635) );
  NAND2X0 U5599 ( .IN1(n6756), .IN2(n6635), .QN(n5781) );
  NOR2X0 U5600 ( .IN1(n9445), .IN2(n9166), .QN(n6243) );
  INVX0 U5601 ( .INP(n6243), .ZN(n8332) );
  OA21X1 U5602 ( .IN1(n9060), .IN2(n8332), .IN3(n9438), .Q(n6762) );
  OA21X1 U5603 ( .IN1(n6762), .IN2(n6651), .IN3(n6234), .Q(n6759) );
  NAND2X0 U5604 ( .IN1(n5781), .IN2(n6759), .QN(\a4/N489 ) );
  NAND2X0 U5605 ( .IN1(n9440), .IN2(n9442), .QN(n8531) );
  INVX0 U5606 ( .INP(n8531), .ZN(n8710) );
  NAND2X0 U5607 ( .IN1(n8710), .IN2(n5423), .QN(n5782) );
  NAND2X0 U5608 ( .IN1(n6759), .IN2(n5782), .QN(\a4/N490 ) );
  NOR2X0 U5609 ( .IN1(n6049), .IN2(n4700), .QN(n7198) );
  NAND2X0 U5610 ( .IN1(n8242), .IN2(n7198), .QN(n5785) );
  NAND2X0 U5611 ( .IN1(n5785), .IN2(n6759), .QN(\a4/N491 ) );
  NAND2X0 U5612 ( .IN1(n6756), .IN2(n7760), .QN(n8209) );
  NAND2X0 U5613 ( .IN1(n8209), .IN2(n6759), .QN(\a1/N488 ) );
  NAND2X0 U5614 ( .IN1(n9436), .IN2(n9082), .QN(n9128) );
  NOR2X0 U5615 ( .IN1(n7600), .IN2(n9128), .QN(n7296) );
  NAND2X0 U5616 ( .IN1(degrees_tmp2[5]), .IN2(n7296), .QN(n8029) );
  NOR2X0 U5617 ( .IN1(n9434), .IN2(n8029), .QN(n6896) );
  INVX0 U5618 ( .INP(n8692), .ZN(n8598) );
  NAND2X0 U5619 ( .IN1(n8598), .IN2(n9433), .QN(n5623) );
  INVX0 U5620 ( .INP(n5623), .ZN(n6678) );
  NAND2X0 U5621 ( .IN1(n9105), .IN2(n6678), .QN(n7738) );
  NOR2X0 U5622 ( .IN1(n5758), .IN2(n6369), .QN(n5353) );
  INVX0 U5623 ( .INP(n5353), .ZN(n7987) );
  INVX0 U5624 ( .INP(n8510), .ZN(n8780) );
  OA22X1 U5625 ( .IN1(n8575), .IN2(n7738), .IN3(n7987), .IN4(n8780), .Q(n4704)
         );
  INVX0 U5626 ( .INP(n5423), .ZN(n7566) );
  NOR2X0 U5627 ( .IN1(n7920), .IN2(n7566), .QN(n6347) );
  NAND2X0 U5628 ( .IN1(n6347), .IN2(n9442), .QN(n7764) );
  INVX0 U5629 ( .INP(n7764), .ZN(n9024) );
  NOR2X0 U5630 ( .IN1(n9434), .IN2(n7679), .QN(n6320) );
  NAND2X0 U5631 ( .IN1(degrees_tmp2[2]), .IN2(n6320), .QN(n9030) );
  NOR2X0 U5632 ( .IN1(n9442), .IN2(n9030), .QN(n6359) );
  NAND2X0 U5633 ( .IN1(n9433), .IN2(n9445), .QN(n7035) );
  INVX0 U5634 ( .INP(n7035), .ZN(n6649) );
  NAND3X0 U5635 ( .IN1(n9435), .IN2(n6649), .IN3(n5750), .QN(n7223) );
  NOR2X0 U5636 ( .IN1(n9441), .IN2(n7223), .QN(n6865) );
  NOR2X0 U5637 ( .IN1(n7600), .IN2(n9046), .QN(n6882) );
  NAND2X0 U5638 ( .IN1(degrees_tmp2[2]), .IN2(n6882), .QN(n8279) );
  INVX0 U5639 ( .INP(n8301), .ZN(n5482) );
  NOR2X0 U5640 ( .IN1(n5433), .IN2(n5482), .QN(n7761) );
  NAND2X0 U5641 ( .IN1(n8575), .IN2(n7761), .QN(n7446) );
  NOR2X0 U5642 ( .IN1(n6322), .IN2(n5623), .QN(n7269) );
  NAND2X0 U5643 ( .IN1(degrees_tmp2[2]), .IN2(n7269), .QN(n8208) );
  NAND2X0 U5644 ( .IN1(n9437), .IN2(n9442), .QN(n6979) );
  INVX0 U5645 ( .INP(n6979), .ZN(n6614) );
  NOR2X0 U5646 ( .IN1(n6614), .IN2(n8684), .QN(n6780) );
  NAND2X0 U5647 ( .IN1(degrees_tmp2[0]), .IN2(n6780), .QN(n4701) );
  NAND4X0 U5648 ( .IN1(n8279), .IN2(n7446), .IN3(n8208), .IN4(n4701), .QN(
        n4702) );
  NOR4X0 U5649 ( .IN1(n9024), .IN2(n6359), .IN3(n6865), .IN4(n4702), .QN(n4703) );
  NAND2X0 U5650 ( .IN1(n6613), .IN2(n9440), .QN(n7649) );
  INVX0 U5651 ( .INP(n7649), .ZN(n7484) );
  NAND2X0 U5652 ( .IN1(n7808), .IN2(n7552), .QN(n5442) );
  INVX0 U5653 ( .INP(n5442), .ZN(n7650) );
  NAND2X0 U5654 ( .IN1(n7484), .IN2(n7650), .QN(n7155) );
  INVX0 U5655 ( .INP(n8431), .ZN(n9023) );
  NOR2X0 U5656 ( .IN1(n9023), .IN2(n9433), .QN(n7451) );
  NAND2X0 U5657 ( .IN1(n8875), .IN2(n7451), .QN(n6701) );
  NAND4X0 U5658 ( .IN1(n4704), .IN2(n4703), .IN3(n7155), .IN4(n6701), .QN(
        n4705) );
  NOR2X0 U5659 ( .IN1(n6896), .IN2(n4705), .QN(n4707) );
  NAND2X0 U5660 ( .IN1(n9434), .IN2(n9433), .QN(n8229) );
  NAND2X0 U5661 ( .IN1(n6613), .IN2(n8022), .QN(n6908) );
  INVX0 U5662 ( .INP(n6908), .ZN(n6665) );
  NAND2X0 U5663 ( .IN1(n6665), .IN2(n9442), .QN(n8563) );
  INVX0 U5664 ( .INP(n8563), .ZN(n8674) );
  NAND2X0 U5665 ( .IN1(n8229), .IN2(n8674), .QN(n4706) );
  NAND2X0 U5666 ( .IN1(n4707), .IN2(n4706), .QN(\a6/N470 ) );
  NAND2X0 U5667 ( .IN1(degrees_tmp2[0]), .IN2(n9445), .QN(n7473) );
  NAND2X0 U5668 ( .IN1(n9434), .IN2(degrees_tmp2[5]), .QN(n8288) );
  NOR2X0 U5669 ( .IN1(n7808), .IN2(n8288), .QN(n7589) );
  NAND2X0 U5670 ( .IN1(n5986), .IN2(n7589), .QN(n8685) );
  NOR2X0 U5671 ( .IN1(n7473), .IN2(n8685), .QN(n7804) );
  INVX0 U5672 ( .INP(n9074), .ZN(n9029) );
  NOR2X0 U5673 ( .IN1(n9080), .IN2(n9029), .QN(n4712) );
  NOR2X0 U5674 ( .IN1(n9181), .IN2(n7510), .QN(n8483) );
  NOR2X0 U5675 ( .IN1(n9435), .IN2(n7784), .QN(n9026) );
  NAND2X0 U5676 ( .IN1(n6119), .IN2(n5832), .QN(n6464) );
  INVX0 U5677 ( .INP(n6464), .ZN(n4708) );
  NOR2X0 U5678 ( .IN1(n8575), .IN2(n9099), .QN(n7935) );
  AO22X1 U5679 ( .IN1(n5949), .IN2(n9026), .IN3(n4708), .IN4(n7935), .Q(n4711)
         );
  NAND2X0 U5680 ( .IN1(n9073), .IN2(n6665), .QN(n5727) );
  NOR2X0 U5681 ( .IN1(n7600), .IN2(n9166), .QN(n6941) );
  INVX0 U5682 ( .INP(n6941), .ZN(n8910) );
  NOR2X0 U5683 ( .IN1(degrees_tmp2[5]), .IN2(n8910), .QN(n6790) );
  INVX0 U5684 ( .INP(n6790), .ZN(n6578) );
  NOR2X0 U5685 ( .IN1(n9213), .IN2(n9048), .QN(n7678) );
  NAND2X0 U5686 ( .IN1(n7678), .IN2(n8041), .QN(n4709) );
  NAND4X0 U5687 ( .IN1(n5727), .IN2(n8042), .IN3(n6578), .IN4(n4709), .QN(
        n4710) );
  NOR4X0 U5688 ( .IN1(n4712), .IN2(n8483), .IN3(n4711), .IN4(n4710), .QN(n4713) );
  INVX0 U5689 ( .INP(n6369), .ZN(n4746) );
  NAND2X0 U5690 ( .IN1(n8301), .IN2(n4746), .QN(n6567) );
  NAND2X0 U5691 ( .IN1(n5986), .IN2(n8198), .QN(n6427) );
  INVX0 U5692 ( .INP(n6427), .ZN(n6417) );
  NAND2X0 U5693 ( .IN1(n6417), .IN2(n8598), .QN(n8267) );
  NOR2X0 U5694 ( .IN1(n9445), .IN2(n8267), .QN(n6672) );
  INVX0 U5695 ( .INP(n6672), .ZN(n8866) );
  NOR2X0 U5696 ( .IN1(n9047), .IN2(n9105), .QN(n6624) );
  NOR2X0 U5697 ( .IN1(n6624), .IN2(n9440), .QN(n6920) );
  NAND3X0 U5698 ( .IN1(n9435), .IN2(n8883), .IN3(n6920), .QN(n8235) );
  NAND4X0 U5699 ( .IN1(n4713), .IN2(n6567), .IN3(n8866), .IN4(n8235), .QN(
        n4714) );
  NOR2X0 U5700 ( .IN1(n7804), .IN2(n4714), .QN(n4716) );
  NAND2X0 U5701 ( .IN1(n6155), .IN2(n9433), .QN(n8597) );
  NOR2X0 U5702 ( .IN1(degrees_tmp2[5]), .IN2(n8597), .QN(n7414) );
  NAND2X0 U5703 ( .IN1(n8531), .IN2(n7414), .QN(n4715) );
  NAND2X0 U5704 ( .IN1(n4716), .IN2(n4715), .QN(\a1/N444 ) );
  NOR2X0 U5705 ( .IN1(n6651), .IN2(n7473), .QN(n8163) );
  INVX0 U5706 ( .INP(n7736), .ZN(n9031) );
  NOR2X0 U5707 ( .IN1(n9031), .IN2(n9073), .QN(n9054) );
  INVX0 U5708 ( .INP(n9054), .ZN(n8947) );
  NAND2X0 U5709 ( .IN1(n8163), .IN2(n8947), .QN(n4718) );
  NOR2X0 U5710 ( .IN1(n9048), .IN2(n6893), .QN(n6983) );
  NAND2X0 U5711 ( .IN1(n6650), .IN2(n6983), .QN(n8747) );
  NAND2X0 U5712 ( .IN1(n7517), .IN2(degrees_tmp2[0]), .QN(n8138) );
  NOR2X0 U5713 ( .IN1(n9213), .IN2(n8138), .QN(n8358) );
  NAND2X0 U5714 ( .IN1(n8358), .IN2(n9433), .QN(n8106) );
  NOR2X0 U5715 ( .IN1(n8213), .IN2(degrees_tmp2[3]), .QN(n7902) );
  NAND2X0 U5716 ( .IN1(n4717), .IN2(n7902), .QN(n8977) );
  INVX0 U5717 ( .INP(n8977), .ZN(n8186) );
  NAND2X0 U5718 ( .IN1(n9125), .IN2(n8186), .QN(n7786) );
  NAND4X0 U5719 ( .IN1(n4718), .IN2(n8747), .IN3(n8106), .IN4(n7786), .QN(
        n4724) );
  NOR2X0 U5720 ( .IN1(n7656), .IN2(n9436), .QN(n6343) );
  NOR2X0 U5721 ( .IN1(n9438), .IN2(n8124), .QN(n9188) );
  INVX0 U5722 ( .INP(n9188), .ZN(n7393) );
  NAND2X0 U5723 ( .IN1(n7517), .IN2(n8220), .QN(n8169) );
  INVX0 U5724 ( .INP(n8169), .ZN(n8697) );
  INVX0 U5725 ( .INP(n5913), .ZN(n4719) );
  NOR2X0 U5726 ( .IN1(n4719), .IN2(n7466), .QN(n6978) );
  NOR2X0 U5727 ( .IN1(n8697), .IN2(n6978), .QN(n4720) );
  OA22X1 U5728 ( .IN1(n6343), .IN2(n7393), .IN3(n4720), .IN4(n7686), .Q(n4722)
         );
  NAND2X0 U5729 ( .IN1(n7936), .IN2(n8467), .QN(n8885) );
  NOR2X0 U5730 ( .IN1(n8675), .IN2(n6017), .QN(n7655) );
  NOR2X0 U5731 ( .IN1(n6651), .IN2(n7920), .QN(n8447) );
  INVX0 U5732 ( .INP(n8447), .ZN(n8495) );
  OA22X1 U5733 ( .IN1(n9082), .IN2(n8885), .IN3(n7655), .IN4(n8495), .Q(n4721)
         );
  OR2X1 U5734 ( .IN1(n9445), .IN2(n7981), .Q(n6249) );
  NAND4X0 U5735 ( .IN1(n4722), .IN2(n4721), .IN3(n6535), .IN4(n6249), .QN(
        n4723) );
  NOR2X0 U5736 ( .IN1(n4724), .IN2(n4723), .QN(n4726) );
  INVX0 U5737 ( .INP(n4728), .ZN(n5761) );
  NAND2X0 U5738 ( .IN1(n5761), .IN2(n5442), .QN(n7596) );
  NOR2X0 U5739 ( .IN1(degrees_tmp2[0]), .IN2(n7596), .QN(n7971) );
  NAND2X0 U5740 ( .IN1(n8511), .IN2(n7971), .QN(n4725) );
  NAND2X0 U5741 ( .IN1(n4726), .IN2(n4725), .QN(\a5/N443 ) );
  NAND2X0 U5742 ( .IN1(n9190), .IN2(n9445), .QN(n7989) );
  NOR2X0 U5743 ( .IN1(n7402), .IN2(n7989), .QN(n7520) );
  NAND2X0 U5744 ( .IN1(degrees_tmp2[0]), .IN2(n7520), .QN(n9178) );
  NOR2X0 U5745 ( .IN1(degrees_tmp2[3]), .IN2(n8169), .QN(n8646) );
  NAND2X0 U5746 ( .IN1(n8646), .IN2(n9442), .QN(n9088) );
  NAND2X0 U5747 ( .IN1(n6649), .IN2(n5626), .QN(n7256) );
  NOR2X0 U5748 ( .IN1(n8883), .IN2(n9213), .QN(n9124) );
  NAND2X0 U5749 ( .IN1(n7700), .IN2(n9124), .QN(n4727) );
  NAND4X0 U5750 ( .IN1(n9178), .IN2(n9088), .IN3(n7256), .IN4(n4727), .QN(
        n4733) );
  NOR2X0 U5751 ( .IN1(degrees_tmp2[3]), .IN2(n8041), .QN(n6067) );
  NOR2X0 U5752 ( .IN1(n8249), .IN2(n4728), .QN(n7208) );
  NAND2X0 U5753 ( .IN1(n6067), .IN2(n7208), .QN(n8933) );
  NAND2X0 U5754 ( .IN1(n8825), .IN2(n6698), .QN(n6916) );
  OA22X1 U5755 ( .IN1(n9434), .IN2(n8933), .IN3(n6916), .IN4(n9442), .Q(n4731)
         );
  NOR2X0 U5756 ( .IN1(n9435), .IN2(n5938), .QN(n7735) );
  NAND2X0 U5757 ( .IN1(n9437), .IN2(n7735), .QN(n9212) );
  INVX0 U5758 ( .INP(n9212), .ZN(n6461) );
  NOR2X0 U5759 ( .IN1(n5938), .IN2(n7808), .QN(n6296) );
  NOR2X0 U5760 ( .IN1(n6461), .IN2(n6296), .QN(n6597) );
  NOR2X0 U5761 ( .IN1(degrees_tmp2[0]), .IN2(n6597), .QN(n6492) );
  NAND2X0 U5762 ( .IN1(n6492), .IN2(n9440), .QN(n6190) );
  NOR2X0 U5763 ( .IN1(n9437), .IN2(n9132), .QN(n5378) );
  NAND2X0 U5764 ( .IN1(n5378), .IN2(n8101), .QN(n8968) );
  NAND3X0 U5765 ( .IN1(n7025), .IN2(n8968), .IN3(n9127), .QN(n4729) );
  NAND2X0 U5766 ( .IN1(n4729), .IN2(n7233), .QN(n4730) );
  NAND2X0 U5767 ( .IN1(degrees_tmp2[3]), .IN2(n9445), .QN(n8645) );
  NAND2X0 U5768 ( .IN1(n8645), .IN2(n9048), .QN(n7597) );
  NOR2X0 U5769 ( .IN1(n9213), .IN2(n7597), .QN(n7698) );
  NAND2X0 U5770 ( .IN1(n9125), .IN2(n7698), .QN(n5466) );
  NAND4X0 U5771 ( .IN1(n4731), .IN2(n6190), .IN3(n4730), .IN4(n5466), .QN(
        n4732) );
  NOR2X0 U5772 ( .IN1(n4733), .IN2(n4732), .QN(n4735) );
  NOR2X0 U5773 ( .IN1(n8947), .IN2(n7649), .QN(n7090) );
  NAND2X0 U5774 ( .IN1(n7090), .IN2(n9441), .QN(n4734) );
  NAND2X0 U5775 ( .IN1(n4735), .IN2(n4734), .QN(\a6/N486 ) );
  NOR2X0 U5776 ( .IN1(n9433), .IN2(n8282), .QN(n6136) );
  NAND2X0 U5777 ( .IN1(n7699), .IN2(n6136), .QN(n6840) );
  NAND2X0 U5778 ( .IN1(n6710), .IN2(n9082), .QN(n5340) );
  OAI21X1 U5779 ( .IN1(n5912), .IN2(n6836), .IN3(n5340), .QN(n7901) );
  NAND2X0 U5780 ( .IN1(n5832), .IN2(n7901), .QN(n6201) );
  NAND2X0 U5781 ( .IN1(n6840), .IN2(n6201), .QN(n6146) );
  NOR2X0 U5782 ( .IN1(degrees_tmp2[0]), .IN2(n7393), .QN(n6213) );
  NAND2X0 U5783 ( .IN1(n9047), .IN2(n6017), .QN(n8737) );
  INVX0 U5784 ( .INP(n8737), .ZN(n8622) );
  INVX0 U5785 ( .INP(n5911), .ZN(n5985) );
  NAND2X0 U5786 ( .IN1(n5936), .IN2(n5985), .QN(n6959) );
  NOR2X0 U5787 ( .IN1(n8754), .IN2(n6959), .QN(n8676) );
  INVX0 U5788 ( .INP(n8073), .ZN(n9208) );
  NOR2X0 U5789 ( .IN1(n9208), .IN2(n6661), .QN(n9183) );
  NAND2X0 U5790 ( .IN1(n9190), .IN2(n9183), .QN(n5894) );
  NAND2X0 U5791 ( .IN1(n9105), .IN2(n8188), .QN(n6205) );
  INVX0 U5792 ( .INP(n6205), .ZN(n5895) );
  NOR2X0 U5793 ( .IN1(n5442), .IN2(n8684), .QN(n7457) );
  NOR2X0 U5794 ( .IN1(n5895), .IN2(n7457), .QN(n4736) );
  OA22X1 U5795 ( .IN1(n9435), .IN2(n5894), .IN3(degrees_tmp2[0]), .IN4(n4736), 
        .Q(n4737) );
  INVX0 U5796 ( .INP(n7402), .ZN(n8890) );
  NOR2X0 U5797 ( .IN1(degrees_tmp2[0]), .IN2(n8213), .QN(n8118) );
  NAND2X0 U5798 ( .IN1(n8890), .IN2(n8118), .QN(n8729) );
  NOR2X0 U5799 ( .IN1(n9434), .IN2(n8729), .QN(n5767) );
  INVX0 U5800 ( .INP(n5767), .ZN(n6588) );
  NOR2X0 U5801 ( .IN1(degrees_tmp2[2]), .IN2(n6588), .QN(n8888) );
  NAND2X0 U5802 ( .IN1(n8888), .IN2(n9441), .QN(n7781) );
  NAND2X0 U5803 ( .IN1(n6461), .IN2(n8787), .QN(n8797) );
  NAND4X0 U5804 ( .IN1(n4737), .IN2(n7662), .IN3(n7781), .IN4(n8797), .QN(
        n4738) );
  OR4X1 U5805 ( .IN1(n6213), .IN2(n8622), .IN3(n8676), .IN4(n4738), .Q(n4739)
         );
  NOR2X0 U5806 ( .IN1(n6146), .IN2(n4739), .QN(n4741) );
  INVX0 U5807 ( .INP(n8529), .ZN(n7876) );
  NOR2X0 U5808 ( .IN1(n7876), .IN2(n8938), .QN(n6090) );
  INVX0 U5809 ( .INP(n8796), .ZN(n8026) );
  NAND2X0 U5810 ( .IN1(n6090), .IN2(n8026), .QN(n4740) );
  NAND2X0 U5811 ( .IN1(n4741), .IN2(n4740), .QN(\a4/N438 ) );
  OR2X1 U5812 ( .IN1(n4743), .IN2(n4742), .Q(n4744) );
  NAND2X0 U5813 ( .IN1(n4745), .IN2(n4744), .QN(N357) );
  NOR2X0 U5814 ( .IN1(n6401), .IN2(n8350), .QN(n5696) );
  INVX0 U5815 ( .INP(n5696), .ZN(n7485) );
  NOR2X0 U5816 ( .IN1(n7485), .IN2(n7473), .QN(n8832) );
  NOR2X0 U5817 ( .IN1(n9149), .IN2(n6651), .QN(n6275) );
  INVX0 U5818 ( .INP(n6275), .ZN(n7234) );
  NOR2X0 U5819 ( .IN1(n8489), .IN2(n7234), .QN(n7827) );
  NAND2X0 U5820 ( .IN1(n8710), .IN2(n6155), .QN(n8578) );
  NOR2X0 U5821 ( .IN1(degrees_tmp2[0]), .IN2(n8578), .QN(n9009) );
  NOR2X0 U5822 ( .IN1(n8213), .IN2(n7209), .QN(n7109) );
  INVX0 U5823 ( .INP(n7109), .ZN(n6612) );
  NOR2X0 U5824 ( .IN1(n5911), .IN2(n6612), .QN(n6231) );
  NOR2X0 U5825 ( .IN1(degrees_tmp2[0]), .IN2(n9060), .QN(n5408) );
  NAND2X0 U5826 ( .IN1(n8220), .IN2(n5408), .QN(n9192) );
  NOR2X0 U5827 ( .IN1(n7717), .IN2(n9192), .QN(n6283) );
  NOR4X0 U5828 ( .IN1(n7827), .IN2(n9009), .IN3(n6231), .IN4(n6283), .QN(n4751) );
  NOR2X0 U5829 ( .IN1(n6205), .IN2(n6836), .QN(n5441) );
  NAND2X0 U5830 ( .IN1(n4746), .IN2(n8118), .QN(n7183) );
  NOR2X0 U5831 ( .IN1(n9442), .IN2(n7183), .QN(n6156) );
  NAND2X0 U5832 ( .IN1(n8119), .IN2(n8118), .QN(n8707) );
  INVX0 U5833 ( .INP(n8707), .ZN(n9033) );
  OA221X1 U5834 ( .IN1(n8898), .IN2(n9033), .IN3(n8898), .IN4(n8947), .IN5(
        n8511), .Q(n4748) );
  NOR2X0 U5835 ( .IN1(n7808), .IN2(n7083), .QN(n9187) );
  NAND2X0 U5836 ( .IN1(n9187), .IN2(n9436), .QN(n8135) );
  NAND3X0 U5837 ( .IN1(degrees_tmp2[2]), .IN2(n8567), .IN3(n8531), .QN(n7838)
         );
  OR2X1 U5838 ( .IN1(n8424), .IN2(n7838), .Q(n4764) );
  NAND4X0 U5839 ( .IN1(n7060), .IN2(n8135), .IN3(n4764), .IN4(n7940), .QN(
        n4747) );
  NOR4X0 U5840 ( .IN1(n5441), .IN2(n6156), .IN3(n4748), .IN4(n4747), .QN(n4750) );
  NOR2X0 U5841 ( .IN1(n8692), .IN2(n6371), .QN(n7483) );
  NAND2X0 U5842 ( .IN1(n7483), .IN2(n9442), .QN(n6696) );
  INVX0 U5843 ( .INP(n6696), .ZN(n6599) );
  NAND2X0 U5844 ( .IN1(degrees_tmp2[2]), .IN2(n6599), .QN(n6799) );
  INVX0 U5845 ( .INP(n8229), .ZN(n8730) );
  NOR2X0 U5846 ( .IN1(n8730), .IN2(n8675), .QN(n8461) );
  NOR2X0 U5847 ( .IN1(n9435), .IN2(n8461), .QN(n6403) );
  NAND2X0 U5848 ( .IN1(n7032), .IN2(n6403), .QN(n4749) );
  NAND4X0 U5849 ( .IN1(n4751), .IN2(n4750), .IN3(n6799), .IN4(n4749), .QN(
        n4752) );
  NOR2X0 U5850 ( .IN1(n8832), .IN2(n4752), .QN(n4754) );
  NOR2X0 U5851 ( .IN1(n9436), .IN2(n8474), .QN(n5516) );
  INVX0 U5852 ( .INP(n5516), .ZN(n7969) );
  NOR2X0 U5853 ( .IN1(n8386), .IN2(n7969), .QN(n6108) );
  NAND2X0 U5854 ( .IN1(n8588), .IN2(n6108), .QN(n4753) );
  NAND2X0 U5855 ( .IN1(n4754), .IN2(n4753), .QN(\a6/N453 ) );
  NAND2X0 U5856 ( .IN1(n6710), .IN2(n9203), .QN(n8515) );
  INVX0 U5857 ( .INP(n8515), .ZN(n9005) );
  NOR2X0 U5858 ( .IN1(n6100), .IN2(n9005), .QN(n7548) );
  NOR4X0 U5859 ( .IN1(n9435), .IN2(n8022), .IN3(n7548), .IN4(n6306), .QN(n5477) );
  NAND2X0 U5860 ( .IN1(n5986), .IN2(n5378), .QN(n9108) );
  NOR2X0 U5861 ( .IN1(n9433), .IN2(n9108), .QN(n5529) );
  INVX0 U5862 ( .INP(n5529), .ZN(n8882) );
  NAND2X0 U5863 ( .IN1(n9435), .IN2(n9441), .QN(n6946) );
  INVX0 U5864 ( .INP(n6946), .ZN(n7184) );
  NAND2X0 U5865 ( .IN1(n7902), .IN2(n7184), .QN(n7467) );
  INVX0 U5866 ( .INP(n7467), .ZN(n5843) );
  NAND2X0 U5867 ( .IN1(n5843), .IN2(n9440), .QN(n6398) );
  INVX0 U5868 ( .INP(n6661), .ZN(n8001) );
  NOR2X0 U5869 ( .IN1(n6398), .IN2(n8001), .QN(n5606) );
  INVX0 U5870 ( .INP(n5606), .ZN(n7225) );
  OA21X1 U5871 ( .IN1(n6836), .IN2(n8882), .IN3(n7225), .Q(n8023) );
  INVX0 U5872 ( .INP(n6487), .ZN(n6952) );
  NOR2X0 U5873 ( .IN1(n9442), .IN2(n6952), .QN(n8855) );
  NOR2X0 U5874 ( .IN1(n7298), .IN2(n7293), .QN(n7964) );
  NOR2X0 U5875 ( .IN1(n4755), .IN2(n5340), .QN(n8097) );
  INVX0 U5876 ( .INP(n8097), .ZN(n8183) );
  NAND3X0 U5877 ( .IN1(n8188), .IN2(n8101), .IN3(n5985), .QN(n7748) );
  NAND2X0 U5878 ( .IN1(n9076), .IN2(n9181), .QN(n9103) );
  NAND2X0 U5879 ( .IN1(n5545), .IN2(n7902), .QN(n8262) );
  INVX0 U5880 ( .INP(n8262), .ZN(n6325) );
  NAND2X0 U5881 ( .IN1(n6325), .IN2(n8171), .QN(n7322) );
  NAND4X0 U5882 ( .IN1(n8183), .IN2(n7748), .IN3(n9103), .IN4(n7322), .QN(
        n4757) );
  INVX0 U5883 ( .INP(n9099), .ZN(n8185) );
  NOR2X0 U5884 ( .IN1(n6651), .IN2(n8185), .QN(n8197) );
  NOR2X0 U5885 ( .IN1(n9438), .IN2(n9436), .QN(n7271) );
  NAND3X0 U5886 ( .IN1(n9082), .IN2(n8220), .IN3(n6836), .QN(n5361) );
  NOR2X0 U5887 ( .IN1(n8995), .IN2(n5361), .QN(n7918) );
  AO22X1 U5888 ( .IN1(n8197), .IN2(n7271), .IN3(n7918), .IN4(n9438), .Q(n4756)
         );
  NOR4X0 U5889 ( .IN1(n8855), .IN2(n7964), .IN3(n4757), .IN4(n4756), .QN(n4759) );
  NOR2X0 U5890 ( .IN1(n8489), .IN2(n9213), .QN(n9150) );
  NAND2X0 U5891 ( .IN1(n9150), .IN2(n9433), .QN(n6985) );
  NAND2X0 U5892 ( .IN1(n9080), .IN2(n7698), .QN(n4758) );
  NAND4X0 U5893 ( .IN1(n8023), .IN2(n4759), .IN3(n6985), .IN4(n4758), .QN(
        n4760) );
  NOR2X0 U5894 ( .IN1(n5477), .IN2(n4760), .QN(n4762) );
  NOR2X0 U5895 ( .IN1(n9440), .IN2(n7596), .QN(n6512) );
  NAND2X0 U5896 ( .IN1(n9209), .IN2(n6512), .QN(n4761) );
  NAND2X0 U5897 ( .IN1(n4762), .IN2(n4761), .QN(\a5/N447 ) );
  INVX0 U5898 ( .INP(n5460), .ZN(n6031) );
  INVX0 U5899 ( .INP(n6120), .ZN(n6623) );
  NAND2X0 U5900 ( .IN1(n8978), .IN2(n6623), .QN(n6060) );
  NAND2X0 U5901 ( .IN1(degrees_tmp2[3]), .IN2(n8760), .QN(n9197) );
  OA22X1 U5902 ( .IN1(n9054), .IN2(n6060), .IN3(n9197), .IN4(n8331), .Q(n4768)
         );
  NAND2X0 U5903 ( .IN1(n5843), .IN2(n7271), .QN(n7335) );
  INVX0 U5904 ( .INP(n7335), .ZN(n5745) );
  NAND2X0 U5905 ( .IN1(n9434), .IN2(n5745), .QN(n6786) );
  NAND2X0 U5906 ( .IN1(n9435), .IN2(n7198), .QN(n6373) );
  NOR2X0 U5907 ( .IN1(n5757), .IN2(n6373), .QN(n6147) );
  INVX0 U5908 ( .INP(n6147), .ZN(n5365) );
  AND2X1 U5909 ( .IN1(n6786), .IN2(n5365), .Q(n8620) );
  NAND2X0 U5910 ( .IN1(n5936), .IN2(n7050), .QN(n8550) );
  OA22X1 U5911 ( .IN1(n8727), .IN2(n7510), .IN3(n7969), .IN4(n8550), .Q(n4766)
         );
  NOR2X0 U5912 ( .IN1(n9108), .IN2(n8595), .QN(n9062) );
  NOR2X0 U5913 ( .IN1(n9032), .IN2(n6371), .QN(n9092) );
  NOR2X0 U5914 ( .IN1(n9062), .IN2(n9092), .QN(n8804) );
  NOR2X0 U5915 ( .IN1(degrees_tmp2[0]), .IN2(n8804), .QN(n7435) );
  NOR2X0 U5916 ( .IN1(n6979), .IN2(n4763), .QN(n9066) );
  INVX0 U5917 ( .INP(n9066), .ZN(n8720) );
  NAND2X0 U5918 ( .IN1(n6619), .IN2(n6613), .QN(n8104) );
  NOR2X0 U5919 ( .IN1(n8909), .IN2(n8104), .QN(n6000) );
  INVX0 U5920 ( .INP(n6000), .ZN(n8399) );
  NAND2X0 U5921 ( .IN1(n8720), .IN2(n8399), .QN(n6162) );
  NOR2X0 U5922 ( .IN1(n7435), .IN2(n6162), .QN(n4765) );
  AND4X1 U5923 ( .IN1(n8620), .IN2(n4766), .IN3(n4765), .IN4(n4764), .Q(n4767)
         );
  NAND2X0 U5924 ( .IN1(n7654), .IN2(n8467), .QN(n7495) );
  NAND2X0 U5925 ( .IN1(n6155), .IN2(n8188), .QN(n7657) );
  NAND2X0 U5926 ( .IN1(n7252), .IN2(n7913), .QN(n7405) );
  OR2X1 U5927 ( .IN1(n7657), .IN2(n7405), .Q(n7938) );
  NAND4X0 U5928 ( .IN1(n4768), .IN2(n4767), .IN3(n7495), .IN4(n7938), .QN(
        n4769) );
  NOR2X0 U5929 ( .IN1(n6031), .IN2(n4769), .QN(n4772) );
  NOR2X0 U5930 ( .IN1(n8240), .IN2(n9082), .QN(n8446) );
  INVX0 U5931 ( .INP(n8446), .ZN(n8145) );
  NOR2X0 U5932 ( .IN1(n7920), .IN2(n4770), .QN(n6934) );
  NAND2X0 U5933 ( .IN1(n8145), .IN2(n6934), .QN(n4771) );
  NAND2X0 U5934 ( .IN1(n4772), .IN2(n4771), .QN(\a2/N440 ) );
  NOR2X0 U5935 ( .IN1(n8041), .IN2(n7600), .QN(n8289) );
  INVX0 U5936 ( .INP(n8289), .ZN(n4773) );
  NAND2X0 U5937 ( .IN1(n7517), .IN2(n8753), .QN(n8926) );
  INVX0 U5938 ( .INP(n7597), .ZN(n8667) );
  NAND2X0 U5939 ( .IN1(n8667), .IN2(n5949), .QN(n6217) );
  NAND4X0 U5940 ( .IN1(n7107), .IN2(n4773), .IN3(n8926), .IN4(n6217), .QN(
        n4778) );
  NAND2X0 U5941 ( .IN1(n9210), .IN2(n8171), .QN(n5488) );
  OR2X1 U5942 ( .IN1(n8645), .IN2(n5488), .Q(n7583) );
  OA22X1 U5943 ( .IN1(n9441), .IN2(n7583), .IN3(n7597), .IN4(n7485), .Q(n4776)
         );
  NOR2X0 U5944 ( .IN1(n9105), .IN2(n8534), .QN(n9205) );
  INVX0 U5945 ( .INP(n6136), .ZN(n4774) );
  NAND2X0 U5946 ( .IN1(n9437), .IN2(n9440), .QN(n5363) );
  NAND2X0 U5947 ( .IN1(n8760), .IN2(n6417), .QN(n8591) );
  OA22X1 U5948 ( .IN1(n9205), .IN2(n4774), .IN3(n5363), .IN4(n8591), .Q(n4775)
         );
  INVX0 U5949 ( .INP(n6347), .ZN(n9110) );
  NAND2X0 U5950 ( .IN1(n9031), .IN2(n5494), .QN(n7377) );
  NAND4X0 U5951 ( .IN1(n4776), .IN2(n4775), .IN3(n9110), .IN4(n7377), .QN(
        n4777) );
  NOR2X0 U5952 ( .IN1(n4778), .IN2(n4777), .QN(n4782) );
  INVX0 U5953 ( .INP(n8302), .ZN(n8317) );
  NAND2X0 U5954 ( .IN1(n9190), .IN2(n9080), .QN(n7392) );
  NAND4X0 U5955 ( .IN1(n4779), .IN2(n8317), .IN3(n8707), .IN4(n7392), .QN(
        n4780) );
  NAND2X0 U5956 ( .IN1(n8825), .IN2(n4780), .QN(n4781) );
  NAND2X0 U5957 ( .IN1(n4782), .IN2(n4781), .QN(\a1/N443 ) );
  NOR2X0 U5958 ( .IN1(rst), .IN2(n5330), .QN(\a7/N37 ) );
  NAND2X0 U5959 ( .IN1(n4787), .IN2(n4789), .QN(n4785) );
  NAND3X0 U5960 ( .IN1(degrees[28]), .IN2(degrees[29]), .IN3(n4785), .QN(n4783) );
  NAND2X0 U5961 ( .IN1(degrees[31]), .IN2(n4783), .QN(n4795) );
  NOR2X0 U5962 ( .IN1(degrees[30]), .IN2(n4795), .QN(n4813) );
  NAND4X0 U5963 ( .IN1(degrees[28]), .IN2(degrees[31]), .IN3(degrees[29]), 
        .IN4(n4785), .QN(n4793) );
  NAND2X0 U5964 ( .IN1(degrees[31]), .IN2(degrees[30]), .QN(n4784) );
  NAND2X0 U5965 ( .IN1(n4793), .IN2(n4784), .QN(n4788) );
  NAND2X0 U5966 ( .IN1(n4785), .IN2(n4788), .QN(n4791) );
  MUX21X1 U5967 ( .IN1(n4792), .IN2(degrees[28]), .S(n4791), .Q(n4811) );
  AND2X1 U5968 ( .IN1(n4789), .IN2(n4788), .Q(n4786) );
  OAI22X1 U5969 ( .IN1(n4787), .IN2(n4786), .IN3(n4785), .IN4(n4784), .QN(
        n4808) );
  MUX21X1 U5970 ( .IN1(degrees[26]), .IN2(n4789), .S(n4788), .Q(n4803) );
  NOR2X0 U5971 ( .IN1(n4803), .IN2(degrees[25]), .QN(n4806) );
  INVX0 U5972 ( .INP(n4806), .ZN(n4790) );
  NAND3X0 U5973 ( .IN1(n4811), .IN2(n4808), .IN3(n4790), .QN(n4797) );
  NOR2X0 U5974 ( .IN1(n4792), .IN2(n4791), .QN(n4794) );
  OA21X1 U5975 ( .IN1(degrees[29]), .IN2(n4794), .IN3(n4793), .Q(n4798) );
  AO21X1 U5976 ( .IN1(n4813), .IN2(n4797), .IN3(n4798), .Q(n4800) );
  AND2X1 U5977 ( .IN1(degrees[30]), .IN2(n4795), .Q(n4814) );
  INVX0 U5978 ( .INP(n4798), .ZN(n4796) );
  NAND2X0 U5979 ( .IN1(n4797), .IN2(n4796), .QN(n4812) );
  AO21X1 U5980 ( .IN1(n4814), .IN2(n4812), .IN3(n4813), .Q(n4801) );
  NAND3X0 U5981 ( .IN1(n4798), .IN2(n4801), .IN3(n4797), .QN(n4799) );
  NAND2X0 U5982 ( .IN1(n4800), .IN2(n4799), .QN(n4831) );
  INVX0 U5983 ( .INP(n4801), .ZN(n4805) );
  MUX21X1 U5984 ( .IN1(n4802), .IN2(degrees[25]), .S(n4805), .Q(n4818) );
  NOR2X0 U5985 ( .IN1(degrees[24]), .IN2(n4818), .QN(n4819) );
  INVX0 U5986 ( .INP(n4819), .ZN(n4807) );
  NOR2X0 U5987 ( .IN1(degrees[25]), .IN2(n4805), .QN(n4804) );
  XOR2X1 U5988 ( .IN1(n4804), .IN2(n4803), .Q(n4820) );
  NOR2X0 U5989 ( .IN1(n4806), .IN2(n4805), .QN(n4809) );
  XOR2X1 U5990 ( .IN1(n4808), .IN2(n4809), .Q(n4823) );
  NAND3X0 U5991 ( .IN1(n4807), .IN2(n4820), .IN3(n4823), .QN(n4826) );
  NAND2X0 U5992 ( .IN1(n4809), .IN2(n4808), .QN(n4810) );
  XOR2X1 U5993 ( .IN1(n4811), .IN2(n4810), .Q(n4828) );
  AND2X1 U5994 ( .IN1(n4826), .IN2(n4828), .Q(n4833) );
  NOR2X0 U5995 ( .IN1(n4831), .IN2(n4833), .QN(n4815) );
  MUX21X1 U5996 ( .IN1(n4814), .IN2(n4813), .S(n4812), .Q(n4829) );
  NOR2X0 U5997 ( .IN1(n4815), .IN2(n4829), .QN(n4824) );
  MUX21X1 U5998 ( .IN1(n4816), .IN2(degrees[24]), .S(n4824), .Q(n4836) );
  NOR2X0 U5999 ( .IN1(n4836), .IN2(degrees[23]), .QN(n4838) );
  NOR2X0 U6000 ( .IN1(degrees[24]), .IN2(n4824), .QN(n4817) );
  XNOR2X1 U6001 ( .IN1(n4818), .IN2(n4817), .Q(n4840) );
  NOR2X0 U6002 ( .IN1(n4838), .IN2(n4840), .QN(n4842) );
  NOR2X0 U6003 ( .IN1(n4819), .IN2(n4824), .QN(n4821) );
  XOR2X1 U6004 ( .IN1(n4821), .IN2(n4820), .Q(n4844) );
  NAND2X0 U6005 ( .IN1(n4842), .IN2(n4844), .QN(n4852) );
  NAND2X0 U6006 ( .IN1(n4821), .IN2(n4820), .QN(n4822) );
  XOR2X1 U6007 ( .IN1(n4823), .IN2(n4822), .Q(n4850) );
  NAND2X0 U6008 ( .IN1(n4852), .IN2(n4850), .QN(n4845) );
  NAND2X0 U6009 ( .IN1(n4829), .IN2(n4826), .QN(n4827) );
  NOR2X0 U6010 ( .IN1(n4828), .IN2(n4824), .QN(n4825) );
  AOI22X1 U6011 ( .IN1(n4828), .IN2(n4827), .IN3(n4826), .IN4(n4825), .QN(
        n4846) );
  AND2X1 U6012 ( .IN1(n4845), .IN2(n4846), .Q(n4834) );
  INVX0 U6013 ( .INP(n4829), .ZN(n4830) );
  NOR2X0 U6014 ( .IN1(n4833), .IN2(n4830), .QN(n4832) );
  MUX21X1 U6015 ( .IN1(n4833), .IN2(n4832), .S(n4831), .Q(n4848) );
  NOR2X0 U6016 ( .IN1(n4834), .IN2(n4848), .QN(n4847) );
  MUX21X1 U6017 ( .IN1(n4835), .IN2(degrees[23]), .S(n4847), .Q(n4855) );
  NOR2X0 U6018 ( .IN1(degrees[22]), .IN2(n4855), .QN(n4857) );
  NOR2X0 U6019 ( .IN1(degrees[23]), .IN2(n4847), .QN(n4837) );
  XNOR2X1 U6020 ( .IN1(n4837), .IN2(n4836), .Q(n4858) );
  NOR2X0 U6021 ( .IN1(n4838), .IN2(n4847), .QN(n4839) );
  XOR2X1 U6022 ( .IN1(n4840), .IN2(n4839), .Q(n4864) );
  NOR3X0 U6023 ( .IN1(n4857), .IN2(n4858), .IN3(n4864), .QN(n4866) );
  INVX0 U6024 ( .INP(n4847), .ZN(n4841) );
  NAND2X0 U6025 ( .IN1(n4842), .IN2(n4841), .QN(n4843) );
  XNOR2X1 U6026 ( .IN1(n4844), .IN2(n4843), .Q(n4870) );
  NOR2X0 U6027 ( .IN1(n4866), .IN2(n4870), .QN(n4875) );
  MUX21X1 U6028 ( .IN1(n4846), .IN2(n4848), .S(n4845), .Q(n4853) );
  INVX0 U6029 ( .INP(n4853), .ZN(n4874) );
  INVX0 U6030 ( .INP(n4875), .ZN(n4873) );
  NOR2X0 U6031 ( .IN1(n4850), .IN2(n4847), .QN(n4851) );
  NAND2X0 U6032 ( .IN1(n4852), .IN2(n4848), .QN(n4849) );
  AO22X1 U6033 ( .IN1(n4852), .IN2(n4851), .IN3(n4850), .IN4(n4849), .Q(n4872)
         );
  NOR2X0 U6034 ( .IN1(n4875), .IN2(n4872), .QN(n4854) );
  NOR2X0 U6035 ( .IN1(n4854), .IN2(n4853), .QN(n4865) );
  NOR2X0 U6036 ( .IN1(degrees[22]), .IN2(n4865), .QN(n4856) );
  XNOR2X1 U6037 ( .IN1(n4856), .IN2(n4855), .Q(n4883) );
  NOR2X0 U6038 ( .IN1(n4857), .IN2(n4865), .QN(n4862) );
  INVX0 U6039 ( .INP(n4858), .ZN(n4861) );
  XNOR2X1 U6040 ( .IN1(n4862), .IN2(n4861), .Q(n4887) );
  OR2X1 U6041 ( .IN1(n4883), .IN2(n4887), .Q(n4860) );
  MUX21X1 U6042 ( .IN1(n4859), .IN2(degrees[22]), .S(n4865), .Q(n4881) );
  NOR2X0 U6043 ( .IN1(degrees[21]), .IN2(n4881), .QN(n4880) );
  NOR2X0 U6044 ( .IN1(n4860), .IN2(n4880), .QN(n4877) );
  NAND2X0 U6045 ( .IN1(n4862), .IN2(n4861), .QN(n4863) );
  XOR2X1 U6046 ( .IN1(n4864), .IN2(n4863), .Q(n4879) );
  NOR2X0 U6047 ( .IN1(n4877), .IN2(n4879), .QN(n4890) );
  OR2X1 U6048 ( .IN1(n4865), .IN2(n4866), .Q(n4869) );
  INVX0 U6049 ( .INP(n4866), .ZN(n4868) );
  NOR2X0 U6050 ( .IN1(n4870), .IN2(n4874), .QN(n4867) );
  AOI22X1 U6051 ( .IN1(n4870), .IN2(n4869), .IN3(n4868), .IN4(n4867), .QN(
        n4891) );
  OR2X1 U6052 ( .IN1(n4890), .IN2(n4891), .Q(n4871) );
  OA221X1 U6053 ( .IN1(n4875), .IN2(n4874), .IN3(n4873), .IN4(n4872), .IN5(
        n4871), .Q(n4888) );
  MUX21X1 U6054 ( .IN1(degrees[21]), .IN2(n4876), .S(n4888), .Q(n4895) );
  NOR2X0 U6055 ( .IN1(n4877), .IN2(n4888), .QN(n4878) );
  XOR2X1 U6056 ( .IN1(n4879), .IN2(n4878), .Q(n4899) );
  NOR2X0 U6057 ( .IN1(n4880), .IN2(n4888), .QN(n4884) );
  XNOR2X1 U6058 ( .IN1(n4883), .IN2(n4884), .Q(n4906) );
  NAND2X0 U6059 ( .IN1(n4895), .IN2(n4896), .QN(n4900) );
  NOR2X0 U6060 ( .IN1(degrees[21]), .IN2(n4888), .QN(n4882) );
  XNOR2X1 U6061 ( .IN1(n4882), .IN2(n4881), .Q(n4903) );
  INVX0 U6062 ( .INP(n4903), .ZN(n4901) );
  NAND3X0 U6063 ( .IN1(n4906), .IN2(n4900), .IN3(n4901), .QN(n4912) );
  INVX0 U6064 ( .INP(n4883), .ZN(n4885) );
  NAND2X0 U6065 ( .IN1(n4885), .IN2(n4884), .QN(n4886) );
  XNOR2X1 U6066 ( .IN1(n4887), .IN2(n4886), .Q(n4908) );
  NAND2X0 U6067 ( .IN1(n4912), .IN2(n4908), .QN(n4897) );
  NAND2X0 U6068 ( .IN1(n4899), .IN2(n4897), .QN(n4893) );
  INVX0 U6069 ( .INP(n4888), .ZN(n4889) );
  NAND2X0 U6070 ( .IN1(n4891), .IN2(n4889), .QN(n4892) );
  MUX21X1 U6071 ( .IN1(n4892), .IN2(n4891), .S(n4890), .Q(n4910) );
  NAND2X0 U6072 ( .IN1(n4893), .IN2(n4910), .QN(n4909) );
  INVX0 U6073 ( .INP(n4909), .ZN(n4904) );
  NOR2X0 U6074 ( .IN1(degrees[20]), .IN2(n4904), .QN(n4894) );
  XNOR2X1 U6075 ( .IN1(n4895), .IN2(n4894), .Q(n4928) );
  MUX21X1 U6076 ( .IN1(n4896), .IN2(degrees[20]), .S(n4909), .Q(n4919) );
  NAND2X0 U6077 ( .IN1(n4919), .IN2(n4921), .QN(n4917) );
  NOR2X0 U6078 ( .IN1(n4899), .IN2(n4904), .QN(n4898) );
  MUX21X1 U6079 ( .IN1(n4899), .IN2(n4898), .S(n4897), .Q(n4922) );
  NAND2X0 U6080 ( .IN1(n4900), .IN2(n4909), .QN(n4902) );
  XNOR2X1 U6081 ( .IN1(n4901), .IN2(n4902), .Q(n4931) );
  NAND3X0 U6082 ( .IN1(n4931), .IN2(n4917), .IN3(n4928), .QN(n4923) );
  INVX0 U6083 ( .INP(n4923), .ZN(n4907) );
  NOR2X0 U6084 ( .IN1(n4903), .IN2(n4902), .QN(n4905) );
  OA22X1 U6085 ( .IN1(n4906), .IN2(n4905), .IN3(n4904), .IN4(n4912), .Q(n4924)
         );
  NOR2X0 U6086 ( .IN1(n4907), .IN2(n4924), .QN(n4936) );
  INVX0 U6087 ( .INP(n4908), .ZN(n4914) );
  NAND2X0 U6088 ( .IN1(n4909), .IN2(n4912), .QN(n4913) );
  NOR2X0 U6089 ( .IN1(n4914), .IN2(n4910), .QN(n4911) );
  AO22X1 U6090 ( .IN1(n4914), .IN2(n4913), .IN3(n4912), .IN4(n4911), .Q(n4935)
         );
  INVX0 U6091 ( .INP(n4935), .ZN(n4915) );
  NOR2X0 U6092 ( .IN1(n4936), .IN2(n4915), .QN(n4916) );
  NOR2X0 U6093 ( .IN1(n4922), .IN2(n4916), .QN(n4920) );
  INVX0 U6094 ( .INP(n4920), .ZN(n4933) );
  AND2X1 U6095 ( .IN1(n4917), .IN2(n4933), .Q(n4929) );
  XOR2X1 U6096 ( .IN1(n4928), .IN2(n4929), .Q(n4939) );
  NOR2X0 U6097 ( .IN1(degrees[19]), .IN2(n4920), .QN(n4918) );
  XNOR2X1 U6098 ( .IN1(n4919), .IN2(n4918), .Q(n4949) );
  MUX21X1 U6099 ( .IN1(n4921), .IN2(degrees[19]), .S(n4920), .Q(n4947) );
  NOR2X0 U6100 ( .IN1(degrees[18]), .IN2(n4947), .QN(n4937) );
  NOR2X0 U6101 ( .IN1(n4935), .IN2(n4936), .QN(n4934) );
  AO21X1 U6102 ( .IN1(n4922), .IN2(n4923), .IN3(n4924), .Q(n4926) );
  NAND3X0 U6103 ( .IN1(n4924), .IN2(n4933), .IN3(n4923), .QN(n4925) );
  NAND2X0 U6104 ( .IN1(n4926), .IN2(n4925), .QN(n4941) );
  NAND2X0 U6105 ( .IN1(n4939), .IN2(n4949), .QN(n4927) );
  NOR2X0 U6106 ( .IN1(n4937), .IN2(n4927), .QN(n4943) );
  NAND2X0 U6107 ( .IN1(n4929), .IN2(n4928), .QN(n4930) );
  XNOR2X1 U6108 ( .IN1(n4931), .IN2(n4930), .Q(n4945) );
  NOR2X0 U6109 ( .IN1(n4943), .IN2(n4945), .QN(n4940) );
  NOR2X0 U6110 ( .IN1(n4941), .IN2(n4940), .QN(n4932) );
  AO221X1 U6111 ( .IN1(n4936), .IN2(n4935), .IN3(n4934), .IN4(n4933), .IN5(
        n4932), .Q(n4951) );
  INVX0 U6112 ( .INP(n4951), .ZN(n4946) );
  NOR2X0 U6113 ( .IN1(n4937), .IN2(n4946), .QN(n4950) );
  NAND2X0 U6114 ( .IN1(n4949), .IN2(n4950), .QN(n4938) );
  XNOR2X1 U6115 ( .IN1(n4939), .IN2(n4938), .Q(n4961) );
  NAND2X0 U6116 ( .IN1(n4941), .IN2(n4951), .QN(n4942) );
  MUX21X1 U6117 ( .IN1(n4942), .IN2(n4941), .S(n4940), .Q(n4957) );
  NOR2X0 U6118 ( .IN1(n4943), .IN2(n4946), .QN(n4944) );
  XNOR2X1 U6119 ( .IN1(n4945), .IN2(n4944), .Q(n4975) );
  INVX0 U6120 ( .INP(n4975), .ZN(n4955) );
  INVX0 U6121 ( .INP(n4961), .ZN(n4954) );
  NOR2X0 U6122 ( .IN1(degrees[18]), .IN2(n4946), .QN(n4948) );
  XNOR2X1 U6123 ( .IN1(n4948), .IN2(n4947), .Q(n4966) );
  XNOR2X1 U6124 ( .IN1(n4950), .IN2(n4949), .Q(n4970) );
  NOR2X0 U6125 ( .IN1(n4966), .IN2(n4970), .QN(n4953) );
  MUX21X1 U6126 ( .IN1(n4952), .IN2(degrees[18]), .S(n4951), .Q(n4965) );
  NAND2X0 U6127 ( .IN1(n4965), .IN2(n4963), .QN(n4962) );
  NAND2X0 U6128 ( .IN1(n4953), .IN2(n4962), .QN(n4959) );
  NAND2X0 U6129 ( .IN1(n4954), .IN2(n4959), .QN(n4973) );
  NAND2X0 U6130 ( .IN1(n4955), .IN2(n4973), .QN(n4956) );
  NAND2X0 U6131 ( .IN1(n4957), .IN2(n4956), .QN(n4972) );
  NAND2X0 U6132 ( .IN1(n4972), .IN2(n4959), .QN(n4960) );
  NOR2X0 U6133 ( .IN1(n4961), .IN2(n4957), .QN(n4958) );
  AO22X1 U6134 ( .IN1(n4961), .IN2(n4960), .IN3(n4959), .IN4(n4958), .Q(n4978)
         );
  AND2X1 U6135 ( .IN1(n4962), .IN2(n4972), .Q(n4967) );
  XNOR2X1 U6136 ( .IN1(n4966), .IN2(n4967), .Q(n4989) );
  MUX21X1 U6137 ( .IN1(n4963), .IN2(degrees[17]), .S(n4972), .Q(n4982) );
  NAND2X0 U6138 ( .IN1(n4982), .IN2(n4977), .QN(n4984) );
  AND2X1 U6139 ( .IN1(n4963), .IN2(n4972), .Q(n4964) );
  XNOR2X1 U6140 ( .IN1(n4965), .IN2(n4964), .Q(n4986) );
  NAND3X0 U6141 ( .IN1(n4989), .IN2(n4984), .IN3(n4986), .QN(n4995) );
  INVX0 U6142 ( .INP(n4966), .ZN(n4968) );
  NAND2X0 U6143 ( .IN1(n4968), .IN2(n4967), .QN(n4969) );
  XOR2X1 U6144 ( .IN1(n4970), .IN2(n4969), .Q(n4997) );
  INVX0 U6145 ( .INP(n4997), .ZN(n4971) );
  NAND2X0 U6146 ( .IN1(n4995), .IN2(n4971), .QN(n4979) );
  NAND2X0 U6147 ( .IN1(n4978), .IN2(n4979), .QN(n4976) );
  NAND2X0 U6148 ( .IN1(n4975), .IN2(n4972), .QN(n4974) );
  MUX21X1 U6149 ( .IN1(n4975), .IN2(n4974), .S(n4973), .Q(n4993) );
  NAND2X0 U6150 ( .IN1(n4976), .IN2(n4993), .QN(n4992) );
  MUX21X1 U6151 ( .IN1(n4977), .IN2(degrees[16]), .S(n4992), .Q(n5002) );
  NAND2X0 U6152 ( .IN1(n5002), .IN2(n5000), .QN(n4999) );
  INVX0 U6153 ( .INP(n4978), .ZN(n4981) );
  NAND2X0 U6154 ( .IN1(n4992), .IN2(n4981), .QN(n4980) );
  MUX21X1 U6155 ( .IN1(n4981), .IN2(n4980), .S(n4979), .Q(n5003) );
  INVX0 U6156 ( .INP(n4992), .ZN(n4990) );
  NOR2X0 U6157 ( .IN1(degrees[16]), .IN2(n4990), .QN(n4983) );
  XNOR2X1 U6158 ( .IN1(n4983), .IN2(n4982), .Q(n5009) );
  AND2X1 U6159 ( .IN1(n4984), .IN2(n4992), .Q(n4987) );
  XOR2X1 U6160 ( .IN1(n4987), .IN2(n4986), .Q(n5011) );
  AND2X1 U6161 ( .IN1(n5009), .IN2(n5011), .Q(n4985) );
  NAND2X0 U6162 ( .IN1(n4985), .IN2(n4999), .QN(n5005) );
  INVX0 U6163 ( .INP(n5005), .ZN(n4991) );
  AND2X1 U6164 ( .IN1(n4987), .IN2(n4986), .Q(n4988) );
  OA22X1 U6165 ( .IN1(n4995), .IN2(n4990), .IN3(n4989), .IN4(n4988), .Q(n5007)
         );
  NOR2X0 U6166 ( .IN1(n4991), .IN2(n5007), .QN(n5013) );
  NAND2X0 U6167 ( .IN1(n4992), .IN2(n4995), .QN(n4996) );
  NOR2X0 U6168 ( .IN1(n4997), .IN2(n4993), .QN(n4994) );
  AOI22X1 U6169 ( .IN1(n4997), .IN2(n4996), .IN3(n4995), .IN4(n4994), .QN(
        n5014) );
  OR2X1 U6170 ( .IN1(n5013), .IN2(n5014), .Q(n4998) );
  NAND2X0 U6171 ( .IN1(n5003), .IN2(n4998), .QN(n5012) );
  AND2X1 U6172 ( .IN1(n4999), .IN2(n5012), .Q(n5008) );
  XOR2X1 U6173 ( .IN1(n5008), .IN2(n5009), .Q(n5019) );
  MUX21X1 U6174 ( .IN1(degrees[15]), .IN2(n5000), .S(n5012), .Q(n5027) );
  NOR2X0 U6175 ( .IN1(n5027), .IN2(degrees[14]), .QN(n5031) );
  AND2X1 U6176 ( .IN1(n5000), .IN2(n5012), .Q(n5001) );
  XOR2X1 U6177 ( .IN1(n5002), .IN2(n5001), .Q(n5033) );
  NOR2X0 U6178 ( .IN1(n5031), .IN2(n5033), .QN(n5017) );
  NAND2X0 U6179 ( .IN1(n5012), .IN2(n5005), .QN(n5006) );
  NOR2X0 U6180 ( .IN1(n5007), .IN2(n5003), .QN(n5004) );
  AO22X1 U6181 ( .IN1(n5007), .IN2(n5006), .IN3(n5005), .IN4(n5004), .Q(n5037)
         );
  NAND2X0 U6182 ( .IN1(n5017), .IN2(n5019), .QN(n5026) );
  NAND2X0 U6183 ( .IN1(n5009), .IN2(n5008), .QN(n5010) );
  XOR2X1 U6184 ( .IN1(n5011), .IN2(n5010), .Q(n5024) );
  NAND2X0 U6185 ( .IN1(n5026), .IN2(n5024), .QN(n5020) );
  NAND2X0 U6186 ( .IN1(n5037), .IN2(n5020), .QN(n5016) );
  NAND2X0 U6187 ( .IN1(n5014), .IN2(n5012), .QN(n5015) );
  MUX21X1 U6188 ( .IN1(n5015), .IN2(n5014), .S(n5013), .Q(n5021) );
  NAND2X0 U6189 ( .IN1(n5016), .IN2(n5021), .QN(n5035) );
  NAND2X0 U6190 ( .IN1(n5017), .IN2(n5035), .QN(n5018) );
  XOR2X1 U6191 ( .IN1(n5019), .IN2(n5018), .Q(n5041) );
  INVX0 U6192 ( .INP(n5020), .ZN(n5038) );
  NOR2X0 U6193 ( .IN1(n5037), .IN2(n5038), .QN(n5036) );
  INVX0 U6194 ( .INP(n5035), .ZN(n5030) );
  NOR2X0 U6195 ( .IN1(n5024), .IN2(n5030), .QN(n5025) );
  INVX0 U6196 ( .INP(n5021), .ZN(n5022) );
  NAND2X0 U6197 ( .IN1(n5026), .IN2(n5022), .QN(n5023) );
  AO22X1 U6198 ( .IN1(n5026), .IN2(n5025), .IN3(n5024), .IN4(n5023), .Q(n5055)
         );
  NOR2X0 U6199 ( .IN1(degrees[14]), .IN2(n5030), .QN(n5028) );
  XOR2X1 U6200 ( .IN1(n5028), .IN2(n5027), .Q(n5048) );
  INVX0 U6201 ( .INP(degrees[14]), .ZN(n5029) );
  MUX21X1 U6202 ( .IN1(n5029), .IN2(degrees[14]), .S(n5030), .Q(n5045) );
  NOR2X0 U6203 ( .IN1(degrees[13]), .IN2(n5045), .QN(n5047) );
  INVX0 U6204 ( .INP(n5047), .ZN(n5042) );
  NOR2X0 U6205 ( .IN1(n5031), .IN2(n5030), .QN(n5032) );
  XNOR2X1 U6206 ( .IN1(n5033), .IN2(n5032), .Q(n5044) );
  NAND3X0 U6207 ( .IN1(n5048), .IN2(n5042), .IN3(n5044), .QN(n5039) );
  AND2X1 U6208 ( .IN1(n5039), .IN2(n5041), .Q(n5054) );
  NOR2X0 U6209 ( .IN1(n5055), .IN2(n5054), .QN(n5034) );
  AO221X1 U6210 ( .IN1(n5038), .IN2(n5037), .IN3(n5036), .IN4(n5035), .IN5(
        n5034), .Q(n5053) );
  NAND2X0 U6211 ( .IN1(n5053), .IN2(n5039), .QN(n5040) );
  XNOR2X1 U6212 ( .IN1(n5041), .IN2(n5040), .Q(n5077) );
  NAND3X0 U6213 ( .IN1(n5042), .IN2(n5053), .IN3(n5048), .QN(n5043) );
  XNOR2X1 U6214 ( .IN1(n5044), .IN2(n5043), .Q(n5073) );
  INVX0 U6215 ( .INP(n5053), .ZN(n5050) );
  NOR2X0 U6216 ( .IN1(degrees[13]), .IN2(n5050), .QN(n5046) );
  XOR2X1 U6217 ( .IN1(n5046), .IN2(n5045), .Q(n5065) );
  NOR2X0 U6218 ( .IN1(n5047), .IN2(n5050), .QN(n5049) );
  XOR2X1 U6219 ( .IN1(n5049), .IN2(n5048), .Q(n5067) );
  NAND2X0 U6220 ( .IN1(n5065), .IN2(n5067), .QN(n5052) );
  MUX21X1 U6221 ( .IN1(degrees[13]), .IN2(n5051), .S(n5050), .Q(n5059) );
  AND2X1 U6222 ( .IN1(n5059), .IN2(n5058), .Q(n5062) );
  NOR2X0 U6223 ( .IN1(n5052), .IN2(n5062), .QN(n5068) );
  NOR2X0 U6224 ( .IN1(n5073), .IN2(n5068), .QN(n5076) );
  OR2X1 U6225 ( .IN1(n5077), .IN2(n5076), .Q(n5057) );
  NAND2X0 U6226 ( .IN1(n5053), .IN2(n5055), .QN(n5056) );
  MUX21X1 U6227 ( .IN1(n5056), .IN2(n5055), .S(n5054), .Q(n5069) );
  NAND2X0 U6228 ( .IN1(n5057), .IN2(n5069), .QN(n5075) );
  INVX0 U6229 ( .INP(n5075), .ZN(n5061) );
  MUX21X1 U6230 ( .IN1(n5058), .IN2(degrees[12]), .S(n5061), .Q(n5090) );
  NOR2X0 U6231 ( .IN1(degrees[11]), .IN2(n5090), .QN(n5087) );
  INVX0 U6232 ( .INP(n5087), .ZN(n5063) );
  NOR2X0 U6233 ( .IN1(degrees[12]), .IN2(n5061), .QN(n5060) );
  XNOR2X1 U6234 ( .IN1(n5060), .IN2(n5059), .Q(n5092) );
  NOR2X0 U6235 ( .IN1(n5062), .IN2(n5061), .QN(n5064) );
  XOR2X1 U6236 ( .IN1(n5064), .IN2(n5065), .Q(n5095) );
  NAND3X0 U6237 ( .IN1(n5063), .IN2(n5092), .IN3(n5095), .QN(n5085) );
  NAND2X0 U6238 ( .IN1(n5065), .IN2(n5064), .QN(n5066) );
  XOR2X1 U6239 ( .IN1(n5067), .IN2(n5066), .Q(n5083) );
  NAND2X0 U6240 ( .IN1(n5085), .IN2(n5083), .QN(n5074) );
  INVX0 U6241 ( .INP(n5074), .ZN(n5100) );
  INVX0 U6242 ( .INP(n5068), .ZN(n5071) );
  NAND2X0 U6243 ( .IN1(n5075), .IN2(n5071), .QN(n5072) );
  NOR2X0 U6244 ( .IN1(n5073), .IN2(n5069), .QN(n5070) );
  AO22X1 U6245 ( .IN1(n5073), .IN2(n5072), .IN3(n5071), .IN4(n5070), .Q(n5099)
         );
  NOR2X0 U6246 ( .IN1(n5099), .IN2(n5100), .QN(n5098) );
  NAND2X0 U6247 ( .IN1(n5099), .IN2(n5074), .QN(n5079) );
  NAND2X0 U6248 ( .IN1(n5077), .IN2(n5075), .QN(n5078) );
  MUX21X1 U6249 ( .IN1(n5078), .IN2(n5077), .S(n5076), .Q(n5080) );
  NAND2X0 U6250 ( .IN1(n5079), .IN2(n5080), .QN(n5097) );
  INVX0 U6251 ( .INP(n5097), .ZN(n5088) );
  NOR2X0 U6252 ( .IN1(n5083), .IN2(n5088), .QN(n5084) );
  INVX0 U6253 ( .INP(n5080), .ZN(n5081) );
  NAND2X0 U6254 ( .IN1(n5085), .IN2(n5081), .QN(n5082) );
  AO22X1 U6255 ( .IN1(n5085), .IN2(n5084), .IN3(n5083), .IN4(n5082), .Q(n5114)
         );
  MUX21X1 U6256 ( .IN1(n5086), .IN2(degrees[11]), .S(n5088), .Q(n5102) );
  NOR2X0 U6257 ( .IN1(degrees[10]), .IN2(n5102), .QN(n5104) );
  NOR2X0 U6258 ( .IN1(n5087), .IN2(n5088), .QN(n5093) );
  XOR2X1 U6259 ( .IN1(n5092), .IN2(n5093), .Q(n5108) );
  NOR2X0 U6260 ( .IN1(degrees[11]), .IN2(n5088), .QN(n5089) );
  XOR2X1 U6261 ( .IN1(n5090), .IN2(n5089), .Q(n5106) );
  NAND2X0 U6262 ( .IN1(n5108), .IN2(n5106), .QN(n5091) );
  NOR2X0 U6263 ( .IN1(n5104), .IN2(n5091), .QN(n5109) );
  NAND2X0 U6264 ( .IN1(n5093), .IN2(n5092), .QN(n5094) );
  XNOR2X1 U6265 ( .IN1(n5095), .IN2(n5094), .Q(n5111) );
  NOR2X0 U6266 ( .IN1(n5109), .IN2(n5111), .QN(n5116) );
  NOR2X0 U6267 ( .IN1(n5114), .IN2(n5116), .QN(n5096) );
  AOI221X1 U6268 ( .IN1(n5100), .IN2(n5099), .IN3(n5098), .IN4(n5097), .IN5(
        n5096), .QN(n5113) );
  MUX21X1 U6269 ( .IN1(n5101), .IN2(degrees[10]), .S(n5113), .Q(n5128) );
  NOR2X0 U6270 ( .IN1(degrees[9]), .IN2(n5128), .QN(n5125) );
  NOR2X0 U6271 ( .IN1(degrees[10]), .IN2(n5113), .QN(n5103) );
  XNOR2X1 U6272 ( .IN1(n5103), .IN2(n5102), .Q(n5129) );
  NOR2X0 U6273 ( .IN1(n5104), .IN2(n5113), .QN(n5105) );
  XNOR2X1 U6274 ( .IN1(n5105), .IN2(n5106), .Q(n5133) );
  NOR3X0 U6275 ( .IN1(n5125), .IN2(n5129), .IN3(n5133), .QN(n5118) );
  NAND2X0 U6276 ( .IN1(n5106), .IN2(n5105), .QN(n5107) );
  XNOR2X1 U6277 ( .IN1(n5108), .IN2(n5107), .Q(n5124) );
  NOR2X0 U6278 ( .IN1(n5118), .IN2(n5124), .QN(n5112) );
  INVX0 U6279 ( .INP(n5112), .ZN(n5136) );
  NOR2X0 U6280 ( .IN1(n5109), .IN2(n5113), .QN(n5110) );
  XNOR2X1 U6281 ( .IN1(n5111), .IN2(n5110), .Q(n5135) );
  NAND2X0 U6282 ( .IN1(n5136), .IN2(n5135), .QN(n5138) );
  NOR2X0 U6283 ( .IN1(n5112), .IN2(n5135), .QN(n5117) );
  NOR2X0 U6284 ( .IN1(n5116), .IN2(n5113), .QN(n5115) );
  MUX21X1 U6285 ( .IN1(n5116), .IN2(n5115), .S(n5114), .Q(n5119) );
  NOR2X0 U6286 ( .IN1(n5117), .IN2(n5119), .QN(n5137) );
  OR2X1 U6287 ( .IN1(n5137), .IN2(n5118), .Q(n5123) );
  INVX0 U6288 ( .INP(n5118), .ZN(n5122) );
  INVX0 U6289 ( .INP(n5119), .ZN(n5120) );
  NOR2X0 U6290 ( .IN1(n5124), .IN2(n5120), .QN(n5121) );
  AO22X1 U6291 ( .IN1(n5124), .IN2(n5123), .IN3(n5122), .IN4(n5121), .Q(n5155)
         );
  NOR2X0 U6292 ( .IN1(n5125), .IN2(n5137), .QN(n5131) );
  XNOR2X1 U6293 ( .IN1(n5129), .IN2(n5131), .Q(n5147) );
  MUX21X1 U6294 ( .IN1(degrees[9]), .IN2(n5126), .S(n5137), .Q(n5142) );
  NAND2X0 U6295 ( .IN1(n5142), .IN2(n5139), .QN(n5140) );
  NOR2X0 U6296 ( .IN1(degrees[9]), .IN2(n5137), .QN(n5127) );
  XOR2X1 U6297 ( .IN1(n5128), .IN2(n5127), .Q(n5144) );
  NAND3X0 U6298 ( .IN1(n5147), .IN2(n5140), .IN3(n5144), .QN(n5148) );
  INVX0 U6299 ( .INP(n5129), .ZN(n5130) );
  NAND2X0 U6300 ( .IN1(n5131), .IN2(n5130), .QN(n5132) );
  XNOR2X1 U6301 ( .IN1(n5133), .IN2(n5132), .Q(n5151) );
  NAND2X0 U6302 ( .IN1(n5148), .IN2(n5151), .QN(n5153) );
  NAND2X0 U6303 ( .IN1(n5155), .IN2(n5153), .QN(n5134) );
  OA221X1 U6304 ( .IN1(n5138), .IN2(n5137), .IN3(n5136), .IN4(n5135), .IN5(
        n5134), .Q(n5152) );
  MUX21X1 U6305 ( .IN1(n5139), .IN2(degrees[8]), .S(n5152), .Q(n5159) );
  NOR2X0 U6306 ( .IN1(degrees[7]), .IN2(n5159), .QN(n5157) );
  INVX0 U6307 ( .INP(n5152), .ZN(n5149) );
  AND2X1 U6308 ( .IN1(n5140), .IN2(n5149), .Q(n5145) );
  XOR2X1 U6309 ( .IN1(n5144), .IN2(n5145), .Q(n5164) );
  NOR2X0 U6310 ( .IN1(degrees[8]), .IN2(n5152), .QN(n5141) );
  XNOR2X1 U6311 ( .IN1(n5142), .IN2(n5141), .Q(n5162) );
  NAND2X0 U6312 ( .IN1(n5164), .IN2(n5162), .QN(n5143) );
  OR2X1 U6313 ( .IN1(n5157), .IN2(n5143), .Q(n5173) );
  NAND2X0 U6314 ( .IN1(n5145), .IN2(n5144), .QN(n5146) );
  XOR2X1 U6315 ( .IN1(n5147), .IN2(n5146), .Q(n5171) );
  AND2X1 U6316 ( .IN1(n5173), .IN2(n5171), .Q(n5167) );
  NAND2X0 U6317 ( .IN1(n5149), .IN2(n5148), .QN(n5150) );
  XNOR2X1 U6318 ( .IN1(n5151), .IN2(n5150), .Q(n5165) );
  NOR2X0 U6319 ( .IN1(n5167), .IN2(n5165), .QN(n5156) );
  NOR2X0 U6320 ( .IN1(n5155), .IN2(n5152), .QN(n5154) );
  MUX21X1 U6321 ( .IN1(n5155), .IN2(n5154), .S(n5153), .Q(n5169) );
  NOR2X0 U6322 ( .IN1(n5156), .IN2(n5169), .QN(n5168) );
  MUX21X1 U6323 ( .IN1(degrees[7]), .IN2(n5244), .S(n5168), .Q(n5182) );
  AND2X1 U6324 ( .IN1(n5251), .IN2(n5182), .Q(n5180) );
  NOR2X0 U6325 ( .IN1(n5157), .IN2(n5168), .QN(n5161) );
  XOR2X1 U6326 ( .IN1(n5162), .IN2(n5161), .Q(n5187) );
  NOR2X0 U6327 ( .IN1(degrees[7]), .IN2(n5168), .QN(n5158) );
  XOR2X1 U6328 ( .IN1(n5159), .IN2(n5158), .Q(n5185) );
  NAND2X0 U6329 ( .IN1(n5187), .IN2(n5185), .QN(n5160) );
  OR2X1 U6330 ( .IN1(n5180), .IN2(n5160), .Q(n5179) );
  NAND2X0 U6331 ( .IN1(n5162), .IN2(n5161), .QN(n5163) );
  XOR2X1 U6332 ( .IN1(n5164), .IN2(n5163), .Q(n5177) );
  NOR2X0 U6333 ( .IN1(n5167), .IN2(n5168), .QN(n5166) );
  MUX21X1 U6334 ( .IN1(n5167), .IN2(n5166), .S(n5165), .Q(n5175) );
  AND2X1 U6335 ( .IN1(n5179), .IN2(n5177), .Q(n5191) );
  NOR2X0 U6336 ( .IN1(n5171), .IN2(n5168), .QN(n5172) );
  NAND2X0 U6337 ( .IN1(n5173), .IN2(n5169), .QN(n5170) );
  AO22X1 U6338 ( .IN1(n5173), .IN2(n5172), .IN3(n5171), .IN4(n5170), .Q(n5189)
         );
  NOR2X0 U6339 ( .IN1(n5191), .IN2(n5189), .QN(n5174) );
  NOR2X0 U6340 ( .IN1(n5175), .IN2(n5174), .QN(n5188) );
  NOR2X0 U6341 ( .IN1(n5177), .IN2(n5188), .QN(n5178) );
  NAND2X0 U6342 ( .IN1(n5179), .IN2(n5175), .QN(n5176) );
  AO22X1 U6343 ( .IN1(n5179), .IN2(n5178), .IN3(n5177), .IN4(n5176), .Q(n5201)
         );
  MUX21X1 U6344 ( .IN1(degrees[6]), .IN2(n5251), .S(n5188), .Q(n5195) );
  AND2X1 U6345 ( .IN1(n5256), .IN2(n5195), .Q(n5193) );
  NOR2X0 U6346 ( .IN1(n5180), .IN2(n5188), .QN(n5184) );
  XOR2X1 U6347 ( .IN1(n5185), .IN2(n5184), .Q(n5200) );
  NOR2X0 U6348 ( .IN1(degrees[6]), .IN2(n5188), .QN(n5181) );
  XNOR2X1 U6349 ( .IN1(n5182), .IN2(n5181), .Q(n5198) );
  NAND2X0 U6350 ( .IN1(n5200), .IN2(n5198), .QN(n5183) );
  OR2X1 U6351 ( .IN1(n5193), .IN2(n5183), .Q(n5209) );
  NAND2X0 U6352 ( .IN1(n5185), .IN2(n5184), .QN(n5186) );
  XOR2X1 U6353 ( .IN1(n5187), .IN2(n5186), .Q(n5207) );
  AND2X1 U6354 ( .IN1(n5209), .IN2(n5207), .Q(n5203) );
  NOR2X0 U6355 ( .IN1(n5201), .IN2(n5203), .QN(n5192) );
  NOR2X0 U6356 ( .IN1(n5191), .IN2(n5188), .QN(n5190) );
  MUX21X1 U6357 ( .IN1(n5191), .IN2(n5190), .S(n5189), .Q(n5205) );
  NOR2X0 U6358 ( .IN1(n5192), .IN2(n5205), .QN(n5204) );
  MUX21X1 U6359 ( .IN1(n5256), .IN2(degrees[5]), .S(n5204), .Q(n5216) );
  NOR2X0 U6360 ( .IN1(degrees[4]), .IN2(n5216), .QN(n5219) );
  NOR2X0 U6361 ( .IN1(n5193), .IN2(n5204), .QN(n5197) );
  XOR2X1 U6362 ( .IN1(n5198), .IN2(n5197), .Q(n5223) );
  NOR2X0 U6363 ( .IN1(degrees[5]), .IN2(n5204), .QN(n5194) );
  XNOR2X1 U6364 ( .IN1(n5195), .IN2(n5194), .Q(n5221) );
  NAND2X0 U6365 ( .IN1(n5223), .IN2(n5221), .QN(n5196) );
  OR2X1 U6366 ( .IN1(n5219), .IN2(n5196), .Q(n5215) );
  NAND2X0 U6367 ( .IN1(n5198), .IN2(n5197), .QN(n5199) );
  XOR2X1 U6368 ( .IN1(n5200), .IN2(n5199), .Q(n5213) );
  NOR2X0 U6369 ( .IN1(n5203), .IN2(n5204), .QN(n5202) );
  MUX21X1 U6370 ( .IN1(n5203), .IN2(n5202), .S(n5201), .Q(n5211) );
  AND2X1 U6371 ( .IN1(n5215), .IN2(n5213), .Q(n5226) );
  NOR2X0 U6372 ( .IN1(n5207), .IN2(n5204), .QN(n5208) );
  NAND2X0 U6373 ( .IN1(n5209), .IN2(n5205), .QN(n5206) );
  AO22X1 U6374 ( .IN1(n5209), .IN2(n5208), .IN3(n5207), .IN4(n5206), .Q(n5227)
         );
  NOR2X0 U6375 ( .IN1(n5226), .IN2(n5227), .QN(n5210) );
  NOR2X0 U6376 ( .IN1(n5211), .IN2(n5210), .QN(n5224) );
  NOR2X0 U6377 ( .IN1(n5213), .IN2(n5224), .QN(n5214) );
  NAND2X0 U6378 ( .IN1(n5215), .IN2(n5211), .QN(n5212) );
  AO22X1 U6379 ( .IN1(n5215), .IN2(n5214), .IN3(n5213), .IN4(n5212), .Q(n5264)
         );
  NOR2X0 U6380 ( .IN1(degrees[4]), .IN2(n5224), .QN(n5217) );
  XNOR2X1 U6381 ( .IN1(n5217), .IN2(n5216), .Q(n5235) );
  MUX21X1 U6382 ( .IN1(n5218), .IN2(degrees[4]), .S(n5224), .Q(n5231) );
  NOR2X0 U6383 ( .IN1(degrees[3]), .IN2(n5231), .QN(n5234) );
  NOR2X0 U6384 ( .IN1(n5219), .IN2(n5224), .QN(n5220) );
  XNOR2X1 U6385 ( .IN1(n5220), .IN2(n5221), .Q(n5236) );
  NOR3X0 U6386 ( .IN1(n5235), .IN2(n5234), .IN3(n5236), .QN(n5239) );
  NAND2X0 U6387 ( .IN1(n5221), .IN2(n5220), .QN(n5222) );
  XNOR2X1 U6388 ( .IN1(n5223), .IN2(n5222), .Q(n5238) );
  NOR2X0 U6389 ( .IN1(n5239), .IN2(n5238), .QN(n5266) );
  NOR2X0 U6390 ( .IN1(n5264), .IN2(n5266), .QN(n5268) );
  INVX0 U6391 ( .INP(n5224), .ZN(n5225) );
  NAND2X0 U6392 ( .IN1(n5227), .IN2(n5225), .QN(n5228) );
  MUX21X1 U6393 ( .IN1(n5228), .IN2(n5227), .S(n5226), .Q(n5229) );
  INVX0 U6394 ( .INP(n5229), .ZN(n5240) );
  NOR2X0 U6395 ( .IN1(n5268), .IN2(n5240), .QN(n5265) );
  NOR2X0 U6396 ( .IN1(degrees[3]), .IN2(n5265), .QN(n5232) );
  AND2X1 U6397 ( .IN1(degrees[3]), .IN2(n5265), .Q(n5230) );
  INVX0 U6398 ( .INP(rst), .ZN(n5269) );
  OA21X1 U6399 ( .IN1(n5232), .IN2(n5230), .IN3(n5269), .Q(\a7/N38 ) );
  XNOR2X1 U6400 ( .IN1(n5232), .IN2(n5231), .Q(n5233) );
  NOR2X0 U6401 ( .IN1(rst), .IN2(n5233), .QN(\a7/N39 ) );
  NOR2X0 U6402 ( .IN1(n5234), .IN2(n5265), .QN(n5261) );
  INVX0 U6403 ( .INP(n5235), .ZN(n5260) );
  NAND2X0 U6404 ( .IN1(n5261), .IN2(n5260), .QN(n5263) );
  XNOR2X1 U6405 ( .IN1(n5236), .IN2(n5263), .Q(n5237) );
  NOR2X0 U6406 ( .IN1(rst), .IN2(n5237), .QN(\a7/N41 ) );
  OA21X1 U6407 ( .IN1(n5239), .IN2(n5265), .IN3(n5238), .Q(n5242) );
  AND2X1 U6408 ( .IN1(n5266), .IN2(n5240), .Q(n5241) );
  OA21X1 U6409 ( .IN1(n5242), .IN2(n5241), .IN3(n5269), .Q(\a7/N42 ) );
  INVX0 U6410 ( .INP(n5243), .ZN(N334) );
  AND2X1 U6411 ( .IN1(n5245), .IN2(n5244), .Q(n5246) );
  MUX21X1 U6412 ( .IN1(degrees_tmp1[7]), .IN2(n5246), .S(n5281), .Q(n4528) );
  MUX21X1 U6413 ( .IN1(degrees_tmp1[1]), .IN2(\a7/N1 ), .S(n5281), .Q(n4522)
         );
  MUX21X1 U6414 ( .IN1(degrees_tmp1[0]), .IN2(\a7/N0 ), .S(n5281), .Q(n4520)
         );
  MUX21X1 U6415 ( .IN1(degrees_tmp1[2]), .IN2(n5330), .S(n5281), .Q(n4523) );
  NOR2X0 U6416 ( .IN1(n5247), .IN2(n5330), .QN(n5249) );
  INVX0 U6417 ( .INP(n5253), .ZN(n5248) );
  OR2X1 U6418 ( .IN1(n5249), .IN2(n5248), .Q(n5250) );
  MUX21X1 U6419 ( .IN1(degrees_tmp1[3]), .IN2(n5250), .S(n5281), .Q(n4524) );
  MUX21X1 U6420 ( .IN1(degrees[6]), .IN2(n5251), .S(n5257), .Q(n5252) );
  MUX21X1 U6421 ( .IN1(degrees_tmp1[6]), .IN2(n5252), .S(n5281), .Q(n4527) );
  NAND2X0 U6422 ( .IN1(degrees[4]), .IN2(n5253), .QN(n5255) );
  OA21X1 U6423 ( .IN1(degrees[4]), .IN2(n5253), .IN3(n5255), .Q(n5254) );
  MUX21X1 U6424 ( .IN1(degrees_tmp1[4]), .IN2(n5254), .S(n5281), .Q(n4525) );
  NAND2X0 U6425 ( .IN1(n5256), .IN2(n5255), .QN(n5258) );
  AND2X1 U6426 ( .IN1(n5258), .IN2(n5257), .Q(n5259) );
  MUX21X1 U6427 ( .IN1(degrees_tmp1[5]), .IN2(n5259), .S(n5281), .Q(n4526) );
  OR2X1 U6428 ( .IN1(n5261), .IN2(n5260), .Q(n5262) );
  AND3X1 U6429 ( .IN1(n5263), .IN2(n5269), .IN3(n5262), .Q(\a7/N40 ) );
  OA21X1 U6430 ( .IN1(n5266), .IN2(n5265), .IN3(n5264), .Q(n5267) );
  NOR3X0 U6431 ( .IN1(rst), .IN2(n5268), .IN3(n5267), .QN(\a7/N43 ) );
  AND2X1 U6432 ( .IN1(\a7/N1 ), .IN2(n5269), .Q(\a7/N36 ) );
  AND2X1 U6433 ( .IN1(\a7/N0 ), .IN2(n5269), .Q(\a7/N35 ) );
  FADDX1 U6434 ( .A(n5272), .B(n5271), .CI(n5270), .CO(n5273), .S(N331) );
  FADDX1 U6435 ( .A(n5275), .B(n5274), .CI(n5273), .CO(n5243), .S(N332) );
  FADDX1 U6436 ( .A(n5278), .B(n5277), .CI(n5276), .CO(n5270), .S(n5279) );
  INVX0 U6437 ( .INP(n5279), .ZN(n5285) );
  NAND2X0 U6438 ( .IN1(n5294), .IN2(degrees[6]), .QN(n5284) );
  NAND2X0 U6439 ( .IN1(divider_out[6]), .IN2(n5319), .QN(n5283) );
  AND2X1 U6440 ( .IN1(n5281), .IN2(n5280), .Q(n5328) );
  NAND2X0 U6441 ( .IN1(degrees_tmp1[6]), .IN2(n5328), .QN(n5282) );
  NAND4X0 U6442 ( .IN1(n5285), .IN2(n5284), .IN3(n5283), .IN4(n5282), .QN(N330) );
  NAND2X0 U6443 ( .IN1(n5294), .IN2(degrees[3]), .QN(n5293) );
  NAND2X0 U6444 ( .IN1(n5328), .IN2(degrees_tmp1[3]), .QN(n5292) );
  FADDX1 U6445 ( .A(n5288), .B(n5287), .CI(n5286), .CO(n5314), .S(n5289) );
  INVX0 U6446 ( .INP(n5289), .ZN(n5291) );
  NAND2X0 U6447 ( .IN1(n5319), .IN2(divider_out[3]), .QN(n5290) );
  NAND4X0 U6448 ( .IN1(n5293), .IN2(n5292), .IN3(n5291), .IN4(n5290), .QN(N327) );
  NAND2X0 U6449 ( .IN1(n5294), .IN2(\a7/N0 ), .QN(n5301) );
  NAND2X0 U6450 ( .IN1(n5328), .IN2(degrees_tmp1[0]), .QN(n5300) );
  AND2X1 U6451 ( .IN1(divider_out[0]), .IN2(n5295), .Q(n5297) );
  XOR2X1 U6452 ( .IN1(n5297), .IN2(n5296), .Q(n5299) );
  NAND2X0 U6453 ( .IN1(n5319), .IN2(divider_out[0]), .QN(n5298) );
  NAND4X0 U6454 ( .IN1(n5301), .IN2(n5300), .IN3(n5299), .IN4(n5298), .QN(N324) );
  FADDX1 U6455 ( .A(n5304), .B(n5303), .CI(n5302), .CO(n5276), .S(n5305) );
  INVX0 U6456 ( .INP(n5305), .ZN(n5313) );
  NOR2X0 U6457 ( .IN1(n5329), .IN2(n5306), .QN(n5318) );
  NAND2X0 U6458 ( .IN1(n5318), .IN2(degrees[5]), .QN(n5312) );
  NAND2X0 U6459 ( .IN1(degrees_tmp1[5]), .IN2(n5328), .QN(n5311) );
  INVX0 U6460 ( .INP(n5307), .ZN(n5309) );
  NAND3X0 U6461 ( .IN1(divider_out[5]), .IN2(n5309), .IN3(n5308), .QN(n5310)
         );
  NAND4X0 U6462 ( .IN1(n5313), .IN2(n5312), .IN3(n5311), .IN4(n5310), .QN(N329) );
  FADDX1 U6463 ( .A(n5316), .B(n5315), .CI(n5314), .CO(n5302), .S(n5317) );
  INVX0 U6464 ( .INP(n5317), .ZN(n5323) );
  NAND2X0 U6465 ( .IN1(n5318), .IN2(degrees[4]), .QN(n5322) );
  NAND2X0 U6466 ( .IN1(n5328), .IN2(degrees_tmp1[4]), .QN(n5321) );
  NAND3X0 U6467 ( .IN1(n5319), .IN2(divider_out[4]), .IN3(n9439), .QN(n5320)
         );
  NAND4X0 U6468 ( .IN1(n5323), .IN2(n5322), .IN3(n5321), .IN4(n5320), .QN(N328) );
  FADDX1 U6469 ( .A(n5326), .B(n5325), .CI(n5324), .CO(n5286), .S(n5327) );
  INVX0 U6470 ( .INP(n5327), .ZN(n5337) );
  NAND2X0 U6471 ( .IN1(n5328), .IN2(degrees_tmp1[2]), .QN(n5336) );
  NOR2X0 U6472 ( .IN1(n5330), .IN2(n5329), .QN(n9219) );
  NAND2X0 U6473 ( .IN1(n9219), .IN2(n5331), .QN(n5335) );
  OR3X1 U6474 ( .IN1(n5333), .IN2(divider_out[7]), .IN3(n5332), .Q(n5334) );
  NAND4X0 U6475 ( .IN1(n5337), .IN2(n5336), .IN3(n5335), .IN4(n5334), .QN(N326) );
  INVX0 U6476 ( .INP(n9108), .ZN(n8180) );
  NAND2X0 U6477 ( .IN1(n8180), .IN2(n5408), .QN(n8713) );
  INVX0 U6478 ( .INP(n8713), .ZN(n7064) );
  NAND2X0 U6479 ( .IN1(n6275), .IN2(n9442), .QN(n7257) );
  NOR2X0 U6480 ( .IN1(n7257), .IN2(n8909), .QN(n6930) );
  NAND2X0 U6481 ( .IN1(n5766), .IN2(n6067), .QN(n6726) );
  NOR2X0 U6482 ( .IN1(n8288), .IN2(n6726), .QN(n6561) );
  NOR4X0 U6483 ( .IN1(n7064), .IN2(n6100), .IN3(n6930), .IN4(n6561), .QN(n5345) );
  NAND2X0 U6484 ( .IN1(n9125), .IN2(n6613), .QN(n7554) );
  NOR2X0 U6485 ( .IN1(n7035), .IN2(n7554), .QN(n7640) );
  NOR2X0 U6486 ( .IN1(degrees_tmp2[3]), .IN2(n8598), .QN(n7213) );
  INVX0 U6487 ( .INP(n6155), .ZN(n7168) );
  NOR2X0 U6488 ( .IN1(n9442), .IN2(n7168), .QN(n6148) );
  OA21X1 U6489 ( .IN1(n7169), .IN2(n7213), .IN3(n6148), .Q(n5339) );
  NOR2X0 U6490 ( .IN1(n7876), .IN2(degrees_tmp2[2]), .QN(n7645) );
  NAND2X0 U6491 ( .IN1(degrees_tmp2[0]), .IN2(n7645), .QN(n6238) );
  NAND2X0 U6492 ( .IN1(n7827), .IN2(n9438), .QN(n7616) );
  NAND2X0 U6493 ( .IN1(n6238), .IN2(n7616), .QN(n8931) );
  NOR2X0 U6494 ( .IN1(degrees_tmp2[5]), .IN2(n5653), .QN(n7167) );
  NAND2X0 U6495 ( .IN1(n7167), .IN2(n6067), .QN(n8167) );
  NOR2X0 U6496 ( .IN1(n8268), .IN2(n8595), .QN(n7355) );
  INVX0 U6497 ( .INP(n8752), .ZN(n8004) );
  NAND2X0 U6498 ( .IN1(n7355), .IN2(n8004), .QN(n7722) );
  NAND4X0 U6499 ( .IN1(n8800), .IN2(n5727), .IN3(n8167), .IN4(n7722), .QN(
        n5338) );
  NOR4X0 U6500 ( .IN1(n7640), .IN2(n5339), .IN3(n8931), .IN4(n5338), .QN(n5344) );
  NAND2X0 U6501 ( .IN1(n8710), .IN2(n8954), .QN(n6878) );
  INVX0 U6502 ( .INP(n5340), .ZN(n5906) );
  NAND2X0 U6503 ( .IN1(n5986), .IN2(n5906), .QN(n6051) );
  NAND2X0 U6504 ( .IN1(n8875), .IN2(n9440), .QN(n8349) );
  NAND3X0 U6505 ( .IN1(n6878), .IN2(n6051), .IN3(n8349), .QN(n5341) );
  NAND2X0 U6506 ( .IN1(degrees_tmp2[3]), .IN2(n9436), .QN(n8649) );
  INVX0 U6507 ( .INP(n8649), .ZN(n6182) );
  NAND2X0 U6508 ( .IN1(n5341), .IN2(n6182), .QN(n5343) );
  NAND2X0 U6509 ( .IN1(n9188), .IN2(n5688), .QN(n5342) );
  NAND4X0 U6510 ( .IN1(n5345), .IN2(n5344), .IN3(n5343), .IN4(n5342), .QN(
        \a6/N437 ) );
  NOR2X0 U6511 ( .IN1(n7035), .IN2(n8190), .QN(n6412) );
  NAND2X0 U6512 ( .IN1(n9435), .IN2(n6412), .QN(n8246) );
  NOR2X0 U6513 ( .IN1(n9437), .IN2(n8246), .QN(n8459) );
  NAND2X0 U6514 ( .IN1(n9182), .IN2(n8240), .QN(n8820) );
  INVX0 U6515 ( .INP(n7746), .ZN(n8512) );
  NAND2X0 U6516 ( .IN1(n9434), .IN2(n8512), .QN(n8438) );
  NAND4X0 U6517 ( .IN1(n8820), .IN2(n8651), .IN3(n8438), .IN4(n7748), .QN(
        n5351) );
  NAND3X0 U6518 ( .IN1(n8188), .IN2(n8220), .IN3(n8431), .QN(n8421) );
  OA22X1 U6519 ( .IN1(n8752), .IN2(n6311), .IN3(n9445), .IN4(n8421), .Q(n5346)
         );
  INVX0 U6520 ( .INP(n7473), .ZN(n7880) );
  NAND2X0 U6521 ( .IN1(n7093), .IN2(n7880), .QN(n9058) );
  NAND3X0 U6522 ( .IN1(n5346), .IN2(n8380), .IN3(n9058), .QN(n5350) );
  NAND2X0 U6523 ( .IN1(n6613), .IN2(n8511), .QN(n6466) );
  NAND2X0 U6524 ( .IN1(n5657), .IN2(n6623), .QN(n8706) );
  OA22X1 U6525 ( .IN1(n7552), .IN2(n6466), .IN3(n7745), .IN4(n8706), .Q(n5348)
         );
  NOR2X0 U6526 ( .IN1(degrees_tmp2[0]), .IN2(n7534), .QN(n8823) );
  NAND3X0 U6527 ( .IN1(n8823), .IN2(n8531), .IN3(n8822), .QN(n5520) );
  INVX0 U6528 ( .INP(n7510), .ZN(n7033) );
  NAND4X0 U6529 ( .IN1(n7033), .IN2(n9433), .IN3(n8041), .IN4(n8282), .QN(
        n5347) );
  NAND2X0 U6530 ( .IN1(n6320), .IN2(n9433), .QN(n9111) );
  INVX0 U6531 ( .INP(n9111), .ZN(n6163) );
  NAND2X0 U6532 ( .IN1(n9435), .IN2(n6163), .QN(n8878) );
  NAND4X0 U6533 ( .IN1(n5348), .IN2(n5520), .IN3(n5347), .IN4(n8878), .QN(
        n5349) );
  OR4X1 U6534 ( .IN1(n8459), .IN2(n5351), .IN3(n5350), .IN4(n5349), .Q(
        \a6/N459 ) );
  NAND2X0 U6535 ( .IN1(n8816), .IN2(n8697), .QN(n7789) );
  NOR2X0 U6536 ( .IN1(degrees_tmp2[5]), .IN2(n7789), .QN(n8310) );
  INVX0 U6537 ( .INP(n9182), .ZN(n7404) );
  NOR2X0 U6538 ( .IN1(n7404), .IN2(n9122), .QN(n6220) );
  INVX0 U6539 ( .INP(n8567), .ZN(n7347) );
  NOR2X0 U6540 ( .IN1(n7347), .IN2(n9122), .QN(n6891) );
  NOR4X0 U6541 ( .IN1(n7486), .IN2(n8310), .IN3(n6220), .IN4(n6891), .QN(n5360) );
  NOR2X0 U6542 ( .IN1(n7291), .IN2(n6013), .QN(n8458) );
  NOR2X0 U6543 ( .IN1(n8213), .IN2(n5912), .QN(n8731) );
  NAND2X0 U6544 ( .IN1(n8731), .IN2(n7784), .QN(n7182) );
  NOR2X0 U6545 ( .IN1(n9434), .IN2(n7182), .QN(n7425) );
  NOR2X0 U6546 ( .IN1(n8458), .IN2(n7425), .QN(n6169) );
  NAND2X0 U6547 ( .IN1(n5832), .IN2(n8300), .QN(n5369) );
  NOR2X0 U6548 ( .IN1(degrees_tmp2[0]), .IN2(n6427), .QN(n7359) );
  INVX0 U6549 ( .INP(n7359), .ZN(n9130) );
  INVX0 U6550 ( .INP(n8550), .ZN(n6274) );
  NAND2X0 U6551 ( .IN1(n6274), .IN2(n9032), .QN(n8020) );
  OA221X1 U6552 ( .IN1(n7745), .IN2(n5369), .IN3(n7745), .IN4(n9130), .IN5(
        n8020), .Q(n5354) );
  NAND2X0 U6553 ( .IN1(degrees_tmp2[5]), .IN2(n5352), .QN(n6135) );
  NAND2X0 U6554 ( .IN1(n6119), .IN2(n5353), .QN(n8835) );
  AND4X1 U6555 ( .IN1(n6169), .IN2(n5354), .IN3(n6135), .IN4(n8835), .Q(n5359)
         );
  NOR2X0 U6556 ( .IN1(n8649), .IN2(n8268), .QN(n8638) );
  NAND2X0 U6557 ( .IN1(n8638), .IN2(n9445), .QN(n7857) );
  NAND3X0 U6558 ( .IN1(n9073), .IN2(n5761), .IN3(n8780), .QN(n5356) );
  NOR2X0 U6559 ( .IN1(n5355), .IN2(n5653), .QN(n6805) );
  INVX0 U6560 ( .INP(n6805), .ZN(n9053) );
  NAND3X0 U6561 ( .IN1(n5356), .IN2(n9053), .IN3(n5975), .QN(n5357) );
  NAND2X0 U6562 ( .IN1(n5357), .IN2(n8995), .QN(n5358) );
  NAND4X0 U6563 ( .IN1(n5360), .IN2(n5359), .IN3(n7857), .IN4(n5358), .QN(
        \a6/N479 ) );
  NAND2X0 U6564 ( .IN1(n7167), .IN2(n8188), .QN(n8996) );
  NOR2X0 U6565 ( .IN1(n8940), .IN2(n8996), .QN(n6333) );
  INVX0 U6566 ( .INP(n7233), .ZN(n9084) );
  AO21X1 U6567 ( .IN1(n8331), .IN2(n5361), .IN3(n9084), .Q(n5362) );
  OA22X1 U6568 ( .IN1(degrees_tmp2[3]), .IN2(n5362), .IN3(n7548), .IN4(n9166), 
        .Q(n5367) );
  NAND2X0 U6569 ( .IN1(n9082), .IN2(n8186), .QN(n7558) );
  NAND2X0 U6570 ( .IN1(n7656), .IN2(n9150), .QN(n6892) );
  NOR2X0 U6571 ( .IN1(n7168), .IN2(n6919), .QN(n5673) );
  NAND2X0 U6572 ( .IN1(n8816), .IN2(n5673), .QN(n8799) );
  INVX0 U6573 ( .INP(n5363), .ZN(n5473) );
  NOR2X0 U6574 ( .IN1(n8940), .IN2(n5473), .QN(n8824) );
  INVX0 U6575 ( .INP(n8824), .ZN(n8630) );
  NAND3X0 U6576 ( .IN1(n7167), .IN2(degrees_tmp2[3]), .IN3(n8630), .QN(n5364)
         );
  AND4X1 U6577 ( .IN1(n7558), .IN2(n6892), .IN3(n8799), .IN4(n5364), .Q(n5366)
         );
  NOR2X0 U6578 ( .IN1(n9433), .IN2(n8474), .QN(n6327) );
  NAND2X0 U6579 ( .IN1(n6327), .IN2(n8302), .QN(n6557) );
  NAND4X0 U6580 ( .IN1(n5367), .IN2(n5366), .IN3(n5365), .IN4(n6557), .QN(
        n5368) );
  AO21X1 U6581 ( .IN1(n6333), .IN2(n9436), .IN3(n5368), .Q(\a6/N487 ) );
  NOR2X0 U6582 ( .IN1(degrees_tmp2[2]), .IN2(n6311), .QN(n8058) );
  NAND2X0 U6583 ( .IN1(degrees_tmp2[0]), .IN2(n8058), .QN(n8454) );
  NAND2X0 U6584 ( .IN1(n9197), .IN2(n9149), .QN(n7528) );
  NAND2X0 U6585 ( .IN1(n7032), .IN2(n7528), .QN(n5933) );
  MUX21X1 U6586 ( .IN1(n8454), .IN2(n5933), .S(n9434), .Q(n5377) );
  NAND2X0 U6587 ( .IN1(degrees_tmp2[2]), .IN2(n8567), .QN(n8423) );
  NOR2X0 U6588 ( .IN1(n8531), .IN2(n8423), .QN(n7192) );
  NAND2X0 U6589 ( .IN1(n8447), .IN2(n9433), .QN(n7174) );
  NOR2X0 U6590 ( .IN1(n9435), .IN2(n7174), .QN(n7415) );
  NOR2X0 U6591 ( .IN1(n9212), .IN2(n8649), .QN(n8324) );
  NAND2X0 U6592 ( .IN1(n9105), .IN2(n8752), .QN(n7638) );
  NOR2X0 U6593 ( .IN1(n9442), .IN2(n7638), .QN(n7507) );
  NOR2X0 U6594 ( .IN1(n8324), .IN2(n7507), .QN(n5809) );
  NAND2X0 U6595 ( .IN1(n5529), .IN2(n8995), .QN(n7730) );
  NOR2X0 U6596 ( .IN1(n9436), .IN2(n7035), .QN(n7049) );
  NAND2X0 U6597 ( .IN1(n6620), .IN2(n7049), .QN(n7065) );
  NOR2X0 U6598 ( .IN1(n9435), .IN2(n5369), .QN(n6068) );
  NAND2X0 U6599 ( .IN1(n6068), .IN2(n9445), .QN(n5370) );
  NAND4X0 U6600 ( .IN1(n5809), .IN2(n7730), .IN3(n7065), .IN4(n5370), .QN(
        n5374) );
  NOR2X0 U6601 ( .IN1(n9434), .IN2(n9108), .QN(n7806) );
  NAND2X0 U6602 ( .IN1(n7806), .IN2(n9436), .QN(n7873) );
  NOR2X0 U6603 ( .IN1(n8190), .IN2(n7945), .QN(n9184) );
  NAND2X0 U6604 ( .IN1(n8649), .IN2(n9149), .QN(n9001) );
  NAND2X0 U6605 ( .IN1(n9184), .IN2(n9001), .QN(n7386) );
  OA22X1 U6606 ( .IN1(n9031), .IN2(n7873), .IN3(n9441), .IN4(n7386), .Q(n5372)
         );
  NOR2X0 U6607 ( .IN1(n8731), .IN2(n7167), .QN(n7391) );
  NOR2X0 U6608 ( .IN1(n7391), .IN2(n8229), .QN(n7970) );
  NAND2X0 U6609 ( .IN1(n7970), .IN2(n9436), .QN(n5371) );
  NOR2X0 U6610 ( .IN1(degrees_tmp2[3]), .IN2(n7291), .QN(n8848) );
  NAND2X0 U6611 ( .IN1(n8848), .IN2(n9442), .QN(n5951) );
  NAND2X0 U6612 ( .IN1(n6182), .IN2(n9188), .QN(n5897) );
  NAND4X0 U6613 ( .IN1(n5372), .IN2(n5371), .IN3(n5951), .IN4(n5897), .QN(
        n5373) );
  NOR4X0 U6614 ( .IN1(n7192), .IN2(n7415), .IN3(n5374), .IN4(n5373), .QN(n5376) );
  NOR2X0 U6615 ( .IN1(n8489), .IN2(n6624), .QN(n6638) );
  INVX0 U6616 ( .INP(n6638), .ZN(n8960) );
  NOR2X0 U6617 ( .IN1(n9434), .IN2(n5938), .QN(n7195) );
  NAND2X0 U6618 ( .IN1(n9435), .IN2(n7195), .QN(n9002) );
  AO221X1 U6619 ( .IN1(n8960), .IN2(n6049), .IN3(n8960), .IN4(n9002), .IN5(
        degrees_tmp2[3]), .Q(n5375) );
  NOR2X0 U6620 ( .IN1(n9440), .IN2(n8842), .QN(n8519) );
  NAND2X0 U6621 ( .IN1(n8699), .IN2(n8519), .QN(n8657) );
  NAND4X0 U6622 ( .IN1(n5377), .IN2(n5376), .IN3(n5375), .IN4(n8657), .QN(
        \a5/N454 ) );
  NOR2X0 U6623 ( .IN1(n9197), .IN2(n8684), .QN(n6352) );
  NAND2X0 U6624 ( .IN1(n6417), .IN2(n6614), .QN(n8880) );
  NOR2X0 U6625 ( .IN1(n8467), .IN2(n8880), .QN(n6221) );
  NOR2X0 U6626 ( .IN1(n6371), .IN2(n8083), .QN(n5958) );
  NOR4X0 U6627 ( .IN1(n8458), .IN2(n6352), .IN3(n6221), .IN4(n5958), .QN(n5384) );
  NOR2X0 U6628 ( .IN1(n9082), .IN2(n9433), .QN(n7417) );
  NAND2X0 U6629 ( .IN1(n6119), .IN2(n5750), .QN(n7875) );
  NAND2X0 U6630 ( .IN1(n8534), .IN2(n8727), .QN(n7939) );
  OA22X1 U6631 ( .IN1(n7417), .IN2(n7875), .IN3(n9433), .IN4(n7939), .Q(n5383)
         );
  NOR2X0 U6632 ( .IN1(n8890), .IN2(n7841), .QN(n6936) );
  NAND2X0 U6633 ( .IN1(n8220), .IN2(n6936), .QN(n5842) );
  NOR2X0 U6634 ( .IN1(n8213), .IN2(n7233), .QN(n6143) );
  NAND2X0 U6635 ( .IN1(n5937), .IN2(n6143), .QN(n8891) );
  INVX0 U6636 ( .INP(n6051), .ZN(n8496) );
  NAND2X0 U6637 ( .IN1(n8496), .IN2(n9433), .QN(n6915) );
  NAND2X0 U6638 ( .IN1(n5378), .IN2(n8301), .QN(n8705) );
  NAND3X0 U6639 ( .IN1(n6060), .IN2(n8705), .IN3(n7393), .QN(n5379) );
  NAND2X0 U6640 ( .IN1(n5379), .IN2(n9073), .QN(n5380) );
  AND4X1 U6641 ( .IN1(n8584), .IN2(n8891), .IN3(n6915), .IN4(n5380), .Q(n5381)
         );
  OA221X1 U6642 ( .IN1(n9061), .IN2(n5975), .IN3(n9061), .IN4(n5842), .IN5(
        n5381), .Q(n5382) );
  NAND2X0 U6643 ( .IN1(n8788), .IN2(n9032), .QN(n7910) );
  NAND4X0 U6644 ( .IN1(n5384), .IN2(n5383), .IN3(n5382), .IN4(n7910), .QN(
        \a4/N459 ) );
  NAND3X0 U6645 ( .IN1(n8249), .IN2(n5913), .IN3(n9442), .QN(n6835) );
  NOR2X0 U6646 ( .IN1(degrees_tmp2[0]), .IN2(n6835), .QN(n8319) );
  NOR2X0 U6647 ( .IN1(n7600), .IN2(n6635), .QN(n7869) );
  INVX0 U6648 ( .INP(n9197), .ZN(n5995) );
  NOR2X0 U6649 ( .IN1(n5995), .IN2(n8728), .QN(n8122) );
  NOR2X0 U6650 ( .IN1(n8122), .IN2(n8268), .QN(n6521) );
  NAND2X0 U6651 ( .IN1(n8754), .IN2(n6805), .QN(n7288) );
  INVX0 U6652 ( .INP(n7632), .ZN(n6925) );
  NAND2X0 U6653 ( .IN1(n9437), .IN2(n6934), .QN(n5385) );
  NAND2X0 U6654 ( .IN1(n7184), .IN2(n6613), .QN(n8470) );
  NAND4X0 U6655 ( .IN1(n6925), .IN2(n5385), .IN3(n8470), .IN4(n7392), .QN(
        n5386) );
  NAND2X0 U6656 ( .IN1(n8825), .IN2(n5386), .QN(n5388) );
  INVX0 U6657 ( .INP(n6412), .ZN(n8261) );
  NOR2X0 U6658 ( .IN1(n9125), .IN2(n6614), .QN(n8528) );
  OR2X1 U6659 ( .IN1(n8261), .IN2(n8528), .Q(n6341) );
  NAND2X0 U6660 ( .IN1(n9105), .IN2(n5516), .QN(n8846) );
  AO21X1 U6661 ( .IN1(n7558), .IN2(n8846), .IN3(n7179), .Q(n5387) );
  NAND4X0 U6662 ( .IN1(n7288), .IN2(n5388), .IN3(n6341), .IN4(n5387), .QN(
        n5389) );
  NOR4X0 U6663 ( .IN1(n8319), .IN2(n7869), .IN3(n6521), .IN4(n5389), .QN(n5390) );
  NAND2X0 U6664 ( .IN1(n8529), .IN2(n9209), .QN(n8336) );
  NAND2X0 U6665 ( .IN1(n8424), .IN2(n6417), .QN(n7839) );
  OR2X1 U6666 ( .IN1(n6049), .IN2(n7839), .Q(n8099) );
  NOR2X0 U6667 ( .IN1(n6651), .IN2(n8645), .QN(n8640) );
  NAND3X0 U6668 ( .IN1(n8640), .IN2(n9438), .IN3(n7945), .QN(n5474) );
  NAND4X0 U6669 ( .IN1(n5390), .IN2(n8336), .IN3(n8099), .IN4(n5474), .QN(
        \a4/N476 ) );
  INVX0 U6670 ( .INP(n9001), .ZN(n8876) );
  NOR2X0 U6671 ( .IN1(n8876), .IN2(n8578), .QN(n5394) );
  NAND2X0 U6672 ( .IN1(n5766), .IN2(n8816), .QN(n7533) );
  NAND2X0 U6673 ( .IN1(n7093), .IN2(n9436), .QN(n6485) );
  NOR2X0 U6674 ( .IN1(n6554), .IN2(n8729), .QN(n7297) );
  INVX0 U6675 ( .INP(n7297), .ZN(n8778) );
  NAND3X0 U6676 ( .IN1(n7533), .IN2(n6485), .IN3(n8778), .QN(n5391) );
  NAND2X0 U6677 ( .IN1(n5391), .IN2(n8572), .QN(n5392) );
  NOR2X0 U6678 ( .IN1(n9445), .IN2(n7876), .QN(n6353) );
  NAND2X0 U6679 ( .IN1(n6353), .IN2(n9166), .QN(n8245) );
  NAND4X0 U6680 ( .IN1(n8380), .IN2(n7940), .IN3(n5392), .IN4(n8245), .QN(
        n5393) );
  NOR3X0 U6681 ( .IN1(n5394), .IN2(n8058), .IN3(n5393), .QN(n5396) );
  NAND2X0 U6682 ( .IN1(n8249), .IN2(n6941), .QN(n7499) );
  NAND2X0 U6683 ( .IN1(n8188), .IN2(n5750), .QN(n7954) );
  NOR2X0 U6684 ( .IN1(n9437), .IN2(n7954), .QN(n5722) );
  NAND2X0 U6685 ( .IN1(n5722), .IN2(n8073), .QN(n5395) );
  NAND4X0 U6686 ( .IN1(n5396), .IN2(n8820), .IN3(n7499), .IN4(n5395), .QN(
        \a4/N485 ) );
  OA22X1 U6687 ( .IN1(n9084), .IN2(n6567), .IN3(n5615), .IN4(n5623), .Q(n5402)
         );
  NOR2X0 U6688 ( .IN1(n9434), .IN2(n6510), .QN(n8468) );
  INVX0 U6689 ( .INP(n8468), .ZN(n9003) );
  NOR2X0 U6690 ( .IN1(n9003), .IN2(n6921), .QN(n8407) );
  NAND2X0 U6691 ( .IN1(degrees_tmp2[2]), .IN2(n9005), .QN(n7445) );
  NOR2X0 U6692 ( .IN1(n7168), .IN2(n9060), .QN(n6360) );
  NAND2X0 U6693 ( .IN1(n9435), .IN2(n6360), .QN(n7378) );
  NAND2X0 U6694 ( .IN1(n7445), .IN2(n7378), .QN(n8559) );
  NAND2X0 U6695 ( .IN1(n7679), .IN2(n6306), .QN(n6709) );
  NAND2X0 U6696 ( .IN1(n6017), .IN2(n6709), .QN(n5397) );
  NAND2X0 U6697 ( .IN1(n6710), .IN2(n8163), .QN(n8304) );
  NOR2X0 U6698 ( .IN1(n6651), .IN2(n9061), .QN(n9172) );
  NAND2X0 U6699 ( .IN1(n9435), .IN2(n9172), .QN(n9050) );
  NAND3X0 U6700 ( .IN1(n5397), .IN2(n8304), .IN3(n9050), .QN(n5400) );
  NAND2X0 U6701 ( .IN1(n8572), .IN2(n6148), .QN(n8070) );
  INVX0 U6702 ( .INP(n7394), .ZN(n8432) );
  NAND2X0 U6703 ( .IN1(n8432), .IN2(n9023), .QN(n7782) );
  INVX0 U6704 ( .INP(n8731), .ZN(n7463) );
  NOR2X0 U6705 ( .IN1(degrees_tmp2[0]), .IN2(n7463), .QN(n8460) );
  NAND2X0 U6706 ( .IN1(n8710), .IN2(n8460), .QN(n7763) );
  INVX0 U6707 ( .INP(n5780), .ZN(n6366) );
  NAND2X0 U6708 ( .IN1(n6366), .IN2(n8001), .QN(n7438) );
  NAND2X0 U6709 ( .IN1(n7093), .IN2(n7438), .QN(n5398) );
  NAND4X0 U6710 ( .IN1(n8070), .IN2(n7782), .IN3(n7763), .IN4(n5398), .QN(
        n5399) );
  NOR4X0 U6711 ( .IN1(n8407), .IN2(n8559), .IN3(n5400), .IN4(n5399), .QN(n5401) );
  INVX0 U6712 ( .INP(n5880), .ZN(n8596) );
  NAND2X0 U6713 ( .IN1(n7050), .IN2(n6143), .QN(n7431) );
  NAND4X0 U6714 ( .IN1(n5402), .IN2(n5401), .IN3(n8596), .IN4(n7431), .QN(
        \a3/N440 ) );
  NOR2X0 U6715 ( .IN1(n7645), .IN2(n8723), .QN(n7821) );
  NAND2X0 U6716 ( .IN1(n9445), .IN2(n6709), .QN(n8530) );
  OA22X1 U6717 ( .IN1(n7821), .IN2(n6836), .IN3(n8530), .IN4(n7209), .Q(n5407)
         );
  NOR2X0 U6718 ( .IN1(n6119), .IN2(n6650), .QN(n8247) );
  AND3X1 U6719 ( .IN1(n6412), .IN2(n8247), .IN3(n9442), .Q(n5405) );
  NAND2X0 U6720 ( .IN1(n5832), .IN2(n5472), .QN(n6967) );
  NOR2X0 U6721 ( .IN1(n9061), .IN2(n6967), .QN(n6399) );
  NAND3X0 U6722 ( .IN1(n8825), .IN2(n7093), .IN3(n9436), .QN(n8347) );
  NAND2X0 U6723 ( .IN1(n7981), .IN2(n8347), .QN(n7795) );
  NAND2X0 U6724 ( .IN1(degrees_tmp2[2]), .IN2(n9172), .QN(n8889) );
  INVX0 U6725 ( .INP(n9032), .ZN(n6194) );
  NAND2X0 U6726 ( .IN1(n6194), .IN2(n6623), .QN(n8763) );
  INVX0 U6727 ( .INP(n8763), .ZN(n7282) );
  NAND2X0 U6728 ( .IN1(n9435), .IN2(n7282), .QN(n8669) );
  OA22X1 U6729 ( .IN1(n6936), .IN2(n8889), .IN3(n9433), .IN4(n8669), .Q(n5403)
         );
  NOR2X0 U6730 ( .IN1(n9434), .IN2(n7600), .QN(n6758) );
  NAND2X0 U6731 ( .IN1(n9080), .IN2(n6758), .QN(n9041) );
  OR2X1 U6732 ( .IN1(n8167), .IN2(n9434), .Q(n6763) );
  NAND2X0 U6733 ( .IN1(n9437), .IN2(n6613), .QN(n8445) );
  INVX0 U6734 ( .INP(n8445), .ZN(n5695) );
  NOR2X0 U6735 ( .IN1(n6649), .IN2(n8461), .QN(n6947) );
  NAND2X0 U6736 ( .IN1(n5695), .IN2(n6947), .QN(n6687) );
  NAND4X0 U6737 ( .IN1(n5403), .IN2(n9041), .IN3(n6763), .IN4(n6687), .QN(
        n5404) );
  NOR4X0 U6738 ( .IN1(n5405), .IN2(n6399), .IN3(n7795), .IN4(n5404), .QN(n5406) );
  NAND2X0 U6739 ( .IN1(degrees_tmp2[3]), .IN2(degrees_tmp2[0]), .QN(n7800) );
  INVX0 U6740 ( .INP(n7800), .ZN(n9037) );
  INVX0 U6741 ( .INP(n6968), .ZN(n7615) );
  NAND2X0 U6742 ( .IN1(n7615), .IN2(n8220), .QN(n5616) );
  NAND2X0 U6743 ( .IN1(n9212), .IN2(n5616), .QN(n7618) );
  NAND2X0 U6744 ( .IN1(n9037), .IN2(n7618), .QN(n5792) );
  NAND3X0 U6745 ( .IN1(n5407), .IN2(n5406), .IN3(n5792), .QN(\a3/N470 ) );
  INVX0 U6746 ( .INP(n5624), .ZN(n5931) );
  NOR2X0 U6747 ( .IN1(n5766), .IN2(n7033), .QN(n5430) );
  NOR2X0 U6748 ( .IN1(n5430), .IN2(n8649), .QN(n7621) );
  OA21X1 U6749 ( .IN1(n6710), .IN2(n5931), .IN3(n7621), .Q(n5412) );
  NOR2X0 U6750 ( .IN1(n9436), .IN2(n6606), .QN(n9156) );
  OA21X1 U6751 ( .IN1(n9156), .IN2(n6983), .IN3(n8041), .Q(n5411) );
  NOR2X0 U6752 ( .IN1(n7600), .IN2(n9181), .QN(n6271) );
  NAND2X0 U6753 ( .IN1(n6271), .IN2(n9032), .QN(n5536) );
  NOR2X0 U6754 ( .IN1(n5408), .IN2(n7169), .QN(n8573) );
  INVX0 U6755 ( .INP(n8573), .ZN(n7239) );
  NAND2X0 U6756 ( .IN1(n6148), .IN2(n7239), .QN(n5409) );
  NAND4X0 U6757 ( .IN1(n8800), .IN2(n6985), .IN3(n5536), .IN4(n5409), .QN(
        n5410) );
  NOR4X0 U6758 ( .IN1(n5412), .IN2(n5411), .IN3(n7795), .IN4(n5410), .QN(n5415) );
  NOR2X0 U6759 ( .IN1(n7416), .IN2(n9435), .QN(n6235) );
  NAND2X0 U6760 ( .IN1(n8000), .IN2(n6235), .QN(n9159) );
  INVX0 U6761 ( .INP(n9159), .ZN(n7354) );
  NAND2X0 U6762 ( .IN1(degrees_tmp2[3]), .IN2(n7354), .QN(n8868) );
  INVX0 U6763 ( .INP(n6322), .ZN(n8826) );
  INVX0 U6764 ( .INP(n8645), .ZN(n9189) );
  NAND3X0 U6765 ( .IN1(n8826), .IN2(n9189), .IN3(n9436), .QN(n8524) );
  NOR2X0 U6766 ( .IN1(n7169), .IN2(n8796), .QN(n8639) );
  NAND2X0 U6767 ( .IN1(n7936), .IN2(n8639), .QN(n6600) );
  NAND3X0 U6768 ( .IN1(n6600), .IN2(n6925), .IN3(n8262), .QN(n5413) );
  NAND2X0 U6769 ( .IN1(n5413), .IN2(n9445), .QN(n5414) );
  NAND4X0 U6770 ( .IN1(n5415), .IN2(n8868), .IN3(n8524), .IN4(n5414), .QN(
        \a2/N473 ) );
  INVX0 U6771 ( .INP(n8684), .ZN(n6392) );
  NAND2X0 U6772 ( .IN1(n6649), .IN2(n9190), .QN(n9100) );
  INVX0 U6773 ( .INP(n9100), .ZN(n7666) );
  NOR2X0 U6774 ( .IN1(n6392), .IN2(n7666), .QN(n5416) );
  NAND2X0 U6775 ( .IN1(n8301), .IN2(n8198), .QN(n8527) );
  NOR2X0 U6776 ( .IN1(n9440), .IN2(n8527), .QN(n6980) );
  INVX0 U6777 ( .INP(n6980), .ZN(n8779) );
  OA22X1 U6778 ( .IN1(n7656), .IN2(n5416), .IN3(n9084), .IN4(n8779), .Q(n5421)
         );
  NOR2X0 U6779 ( .IN1(n6946), .IN2(n6427), .QN(n8330) );
  NOR2X0 U6780 ( .IN1(n6296), .IN2(n8330), .QN(n7588) );
  INVX0 U6781 ( .INP(n7011), .ZN(n7858) );
  NAND2X0 U6782 ( .IN1(n9082), .IN2(n7858), .QN(n6937) );
  NAND2X0 U6783 ( .IN1(n6758), .IN2(n7760), .QN(n5418) );
  NAND2X0 U6784 ( .IN1(n6353), .IN2(n9181), .QN(n5417) );
  AND4X1 U6785 ( .IN1(n7588), .IN2(n6937), .IN3(n5418), .IN4(n5417), .Q(n5420)
         );
  NAND2X0 U6786 ( .IN1(n8000), .IN2(n5419), .QN(n7585) );
  NAND2X0 U6787 ( .IN1(n6119), .IN2(n6620), .QN(n7633) );
  NAND4X0 U6788 ( .IN1(n5421), .IN2(n5420), .IN3(n7585), .IN4(n7633), .QN(
        \a2/N485 ) );
  NOR2X0 U6789 ( .IN1(n7402), .IN2(n5803), .QN(n8379) );
  NOR2X0 U6790 ( .IN1(n5938), .IN2(n8282), .QN(n7809) );
  NAND2X0 U6791 ( .IN1(n7809), .IN2(n9060), .QN(n7834) );
  NOR2X0 U6792 ( .IN1(n8728), .IN2(n7394), .QN(n8162) );
  NAND2X0 U6793 ( .IN1(n9434), .IN2(n8162), .QN(n7743) );
  NOR2X0 U6794 ( .IN1(n6510), .IN2(n7402), .QN(n8566) );
  NAND2X0 U6795 ( .IN1(n8566), .IN2(n9060), .QN(n5422) );
  NAND4X0 U6796 ( .IN1(n7834), .IN2(n7743), .IN3(n6135), .IN4(n5422), .QN(
        n5428) );
  NAND2X0 U6797 ( .IN1(n6155), .IN2(n8728), .QN(n6888) );
  NOR2X0 U6798 ( .IN1(n9440), .IN2(n6888), .QN(n8272) );
  NAND2X0 U6799 ( .IN1(n8272), .IN2(n9433), .QN(n9112) );
  NAND2X0 U6800 ( .IN1(n5423), .IN2(n7437), .QN(n8869) );
  NAND2X0 U6801 ( .IN1(n8728), .IN2(n8468), .QN(n8817) );
  NAND4X0 U6802 ( .IN1(n9112), .IN2(n8869), .IN3(n8817), .IN4(n8584), .QN(
        n5427) );
  NAND2X0 U6803 ( .IN1(n7359), .IN2(n9440), .QN(n7471) );
  NAND2X0 U6804 ( .IN1(n6859), .IN2(n9440), .QN(n9129) );
  NAND3X0 U6805 ( .IN1(n7471), .IN2(n7679), .IN3(n9129), .QN(n5424) );
  NAND2X0 U6806 ( .IN1(n5424), .IN2(n8575), .QN(n5425) );
  NAND2X0 U6807 ( .IN1(n9125), .IN2(n6412), .QN(n8673) );
  NAND4X0 U6808 ( .IN1(n6398), .IN2(n5425), .IN3(n8713), .IN4(n8673), .QN(
        n5426) );
  NOR4X0 U6809 ( .IN1(n8379), .IN2(n5428), .IN3(n5427), .IN4(n5426), .QN(n5429) );
  NOR2X0 U6810 ( .IN1(n9445), .IN2(n8842), .QN(n7518) );
  NAND2X0 U6811 ( .IN1(n7518), .IN2(n9440), .QN(n8131) );
  NOR2X0 U6812 ( .IN1(n9433), .IN2(n9181), .QN(n5708) );
  NAND2X0 U6813 ( .IN1(n9182), .IN2(n5708), .QN(n6845) );
  NAND4X0 U6814 ( .IN1(n5429), .IN2(n8131), .IN3(n7857), .IN4(n6845), .QN(
        \a1/N449 ) );
  NAND3X0 U6815 ( .IN1(n8185), .IN2(n6274), .IN3(n8073), .QN(n5527) );
  OA21X1 U6816 ( .IN1(n5430), .IN2(n8282), .IN3(n5527), .Q(n5438) );
  NOR2X0 U6817 ( .IN1(n9435), .IN2(n8268), .QN(n7816) );
  NOR3X0 U6818 ( .IN1(n5696), .IN2(n7816), .IN3(n6392), .QN(n5431) );
  OA22X1 U6819 ( .IN1(n9084), .IN2(n5803), .IN3(n5431), .IN4(n8649), .Q(n5437)
         );
  NAND2X0 U6820 ( .IN1(n9182), .IN2(n9433), .QN(n8922) );
  NOR2X0 U6821 ( .IN1(n9436), .IN2(n8922), .QN(n7358) );
  INVX0 U6822 ( .INP(n5643), .ZN(n5432) );
  NOR2X0 U6823 ( .IN1(n5433), .IN2(n5432), .QN(n5751) );
  INVX0 U6824 ( .INP(n8188), .ZN(n8588) );
  NOR2X0 U6825 ( .IN1(n5965), .IN2(n7271), .QN(n6575) );
  INVX0 U6826 ( .INP(n6575), .ZN(n8987) );
  NOR2X0 U6827 ( .IN1(n8588), .IN2(n8987), .QN(n6508) );
  AND2X1 U6828 ( .IN1(n8220), .IN2(n6508), .Q(n5435) );
  NAND2X0 U6829 ( .IN1(degrees_tmp2[0]), .IN2(n8097), .QN(n6414) );
  NOR2X0 U6830 ( .IN1(n7252), .IN2(n6651), .QN(n9195) );
  NAND2X0 U6831 ( .IN1(n9195), .IN2(n9445), .QN(n6286) );
  NOR2X0 U6832 ( .IN1(n6306), .IN2(n8645), .QN(n7843) );
  NAND2X0 U6833 ( .IN1(n7843), .IN2(n9441), .QN(n8624) );
  NAND3X0 U6834 ( .IN1(n5739), .IN2(n8978), .IN3(n7784), .QN(n7362) );
  NAND4X0 U6835 ( .IN1(n6414), .IN2(n6286), .IN3(n8624), .IN4(n7362), .QN(
        n5434) );
  NOR4X0 U6836 ( .IN1(n7358), .IN2(n5751), .IN3(n5435), .IN4(n5434), .QN(n5436) );
  NAND4X0 U6837 ( .IN1(n5438), .IN2(n5437), .IN3(n5436), .IN4(n6892), .QN(
        \a1/N477 ) );
  NOR2X0 U6838 ( .IN1(n7746), .IN2(n7571), .QN(n5440) );
  AO22X1 U6839 ( .IN1(n8496), .IN2(n7784), .IN3(n7645), .IN4(n8171), .Q(n7630)
         );
  INVX0 U6840 ( .INP(n7761), .ZN(n9020) );
  NAND2X0 U6841 ( .IN1(n7654), .IN2(n9433), .QN(n7308) );
  INVX0 U6842 ( .INP(n5616), .ZN(n7311) );
  NAND2X0 U6843 ( .IN1(n8752), .IN2(n7311), .QN(n6517) );
  NAND4X0 U6844 ( .IN1(n9020), .IN2(n8563), .IN3(n7308), .IN4(n6517), .QN(
        n5439) );
  NOR4X0 U6845 ( .IN1(n5441), .IN2(n5440), .IN3(n7630), .IN4(n5439), .QN(n5445) );
  NAND2X0 U6846 ( .IN1(n8534), .IN2(n6136), .QN(n8492) );
  INVX0 U6847 ( .INP(n8247), .ZN(n7914) );
  AO221X1 U6848 ( .IN1(n8778), .IN2(n5938), .IN3(n8778), .IN4(n7914), .IN5(
        n8568), .Q(n5444) );
  NAND2X0 U6849 ( .IN1(n9436), .IN2(n5442), .QN(n7388) );
  NAND2X0 U6850 ( .IN1(n7808), .IN2(n7388), .QN(n6391) );
  NAND3X0 U6851 ( .IN1(n5750), .IN2(n9435), .IN3(n6391), .QN(n5734) );
  OR2X1 U6852 ( .IN1(n9445), .IN2(n5734), .Q(n5443) );
  NAND4X0 U6853 ( .IN1(n5445), .IN2(n8492), .IN3(n5444), .IN4(n5443), .QN(
        \a6/N436 ) );
  INVX0 U6854 ( .INP(n7763), .ZN(n5449) );
  NOR2X0 U6855 ( .IN1(n6651), .IN2(n7945), .QN(n8988) );
  AND2X1 U6856 ( .IN1(degrees_tmp2[2]), .IN2(n8988), .Q(n5448) );
  NAND2X0 U6857 ( .IN1(n9436), .IN2(n7945), .QN(n7897) );
  NOR2X0 U6858 ( .IN1(n6371), .IN2(n7897), .QN(n6545) );
  INVX0 U6859 ( .INP(n6545), .ZN(n8252) );
  NAND4X0 U6860 ( .IN1(n7394), .IN2(n7293), .IN3(n8685), .IN4(n8252), .QN(
        n5447) );
  NAND2X0 U6861 ( .IN1(n6859), .IN2(n7169), .QN(n8007) );
  NAND2X0 U6862 ( .IN1(n8988), .IN2(n9438), .QN(n8751) );
  NAND2X0 U6863 ( .IN1(n8978), .IN2(n6016), .QN(n8925) );
  NAND4X0 U6864 ( .IN1(n7873), .IN2(n8007), .IN3(n8751), .IN4(n8925), .QN(
        n5446) );
  NOR4X0 U6865 ( .IN1(n5449), .IN2(n5448), .IN3(n5447), .IN4(n5446), .QN(n5451) );
  NAND2X0 U6866 ( .IN1(n8220), .IN2(n5872), .QN(n5450) );
  NAND4X0 U6867 ( .IN1(n5451), .IN2(n6135), .IN3(n9159), .IN4(n5450), .QN(
        \a6/N438 ) );
  NOR2X0 U6868 ( .IN1(n6650), .IN2(n6915), .QN(n5459) );
  NAND2X0 U6869 ( .IN1(n8000), .IN2(n7921), .QN(n8053) );
  NAND4X0 U6870 ( .IN1(n9041), .IN2(n5727), .IN3(n7378), .IN4(n8053), .QN(
        n5458) );
  INVX0 U6871 ( .INP(n9127), .ZN(n9014) );
  NAND2X0 U6872 ( .IN1(n9014), .IN2(n9181), .QN(n6298) );
  NAND3X0 U6873 ( .IN1(n8754), .IN2(n8753), .IN3(n9438), .QN(n7172) );
  INVX0 U6874 ( .INP(n8288), .ZN(n6434) );
  NAND3X0 U6875 ( .IN1(n8875), .IN2(n6434), .IN3(n9433), .QN(n6904) );
  NAND3X0 U6876 ( .IN1(n6298), .IN2(n7172), .IN3(n6904), .QN(n5457) );
  NOR2X0 U6877 ( .IN1(n6554), .IN2(n6322), .QN(n7133) );
  INVX0 U6878 ( .INP(n7133), .ZN(n6150) );
  NOR2X0 U6879 ( .IN1(n6150), .IN2(n8724), .QN(n7908) );
  NOR2X0 U6880 ( .IN1(n6891), .IN2(n7908), .QN(n5831) );
  NAND2X0 U6881 ( .IN1(n8816), .IN2(n8354), .QN(n7034) );
  NAND2X0 U6882 ( .IN1(n7699), .IN2(n9209), .QN(n7965) );
  NAND3X0 U6883 ( .IN1(n7034), .IN2(n7965), .IN3(n9053), .QN(n5452) );
  NAND2X0 U6884 ( .IN1(n5452), .IN2(n8572), .QN(n5455) );
  NAND2X0 U6885 ( .IN1(n9433), .IN2(n9166), .QN(n6804) );
  NAND3X0 U6886 ( .IN1(n9182), .IN2(n8073), .IN3(n6804), .QN(n5454) );
  INVX0 U6887 ( .INP(n8727), .ZN(n9019) );
  NAND2X0 U6888 ( .IN1(n9092), .IN2(n9019), .QN(n5453) );
  NAND4X0 U6889 ( .IN1(n5831), .IN2(n5455), .IN3(n5454), .IN4(n5453), .QN(
        n5456) );
  OR4X1 U6890 ( .IN1(n5459), .IN2(n5458), .IN3(n5457), .IN4(n5456), .Q(
        \a6/N439 ) );
  NOR2X0 U6891 ( .IN1(n7945), .IN2(n6371), .QN(n8005) );
  NOR2X0 U6892 ( .IN1(n7358), .IN2(n8005), .QN(n7604) );
  NOR2X0 U6893 ( .IN1(n8649), .IN2(n6322), .QN(n6782) );
  NAND2X0 U6894 ( .IN1(n6782), .IN2(n9441), .QN(n8406) );
  OA22X1 U6895 ( .IN1(degrees_tmp2[0]), .IN2(n5460), .IN3(n9440), .IN4(n8406), 
        .Q(n5465) );
  INVX0 U6896 ( .INP(n7654), .ZN(n6811) );
  NOR2X0 U6897 ( .IN1(n8883), .IN2(n9442), .QN(n8484) );
  OA22X1 U6898 ( .IN1(n8675), .IN2(n6811), .IN3(n8484), .IN4(n7534), .Q(n5463)
         );
  NAND2X0 U6899 ( .IN1(n9190), .IN2(n7880), .QN(n9027) );
  NAND2X0 U6900 ( .IN1(n9105), .IN2(n6836), .QN(n5632) );
  NOR2X0 U6901 ( .IN1(n9434), .IN2(n8821), .QN(n6528) );
  NOR2X0 U6902 ( .IN1(n8727), .IN2(n7566), .QN(n8112) );
  NOR2X0 U6903 ( .IN1(n8350), .IN2(n8138), .QN(n8359) );
  NOR4X0 U6904 ( .IN1(n6528), .IN2(n8112), .IN3(n6672), .IN4(n8359), .QN(n5461) );
  OA221X1 U6905 ( .IN1(n8595), .IN2(n9027), .IN3(n8595), .IN4(n5632), .IN5(
        n5461), .Q(n5462) );
  NOR2X0 U6906 ( .IN1(n7600), .IN2(n8282), .QN(n7063) );
  NAND2X0 U6907 ( .IN1(n8249), .IN2(n7063), .QN(n7450) );
  NAND2X0 U6908 ( .IN1(n8408), .IN2(n8041), .QN(n6264) );
  AND4X1 U6909 ( .IN1(n5463), .IN2(n5462), .IN3(n7450), .IN4(n6264), .Q(n5464)
         );
  NAND4X0 U6910 ( .IN1(n7604), .IN2(n5465), .IN3(n5464), .IN4(n7781), .QN(
        \a6/N440 ) );
  NOR2X0 U6911 ( .IN1(n9436), .IN2(n7596), .QN(n7703) );
  NAND2X0 U6912 ( .IN1(n8575), .IN2(n7703), .QN(n8664) );
  NOR2X0 U6913 ( .IN1(n9440), .IN2(n8664), .QN(n5471) );
  NOR2X0 U6914 ( .IN1(n7035), .IN2(n6893), .QN(n5971) );
  NAND2X0 U6915 ( .IN1(n5971), .IN2(n8282), .QN(n8694) );
  NAND4X0 U6916 ( .IN1(n6414), .IN2(n8694), .IN3(n7335), .IN4(n8042), .QN(
        n5470) );
  NAND2X0 U6917 ( .IN1(n6649), .IN2(n7816), .QN(n7111) );
  NOR2X0 U6918 ( .IN1(n8568), .IN2(n6306), .QN(n6523) );
  NAND2X0 U6919 ( .IN1(n6523), .IN2(n9441), .QN(n8156) );
  NAND4X0 U6920 ( .IN1(n5466), .IN2(n7111), .IN3(n8156), .IN4(n7495), .QN(
        n5469) );
  NAND2X0 U6921 ( .IN1(n6296), .IN2(n9442), .QN(n8126) );
  NOR2X0 U6922 ( .IN1(n9445), .IN2(n7987), .QN(n7934) );
  NAND2X0 U6923 ( .IN1(n6650), .IN2(n7934), .QN(n5837) );
  NOR2X0 U6924 ( .IN1(n9433), .IN2(n6836), .QN(n8955) );
  NAND2X0 U6925 ( .IN1(n7208), .IN2(n8955), .QN(n5467) );
  NAND4X0 U6926 ( .IN1(n5734), .IN2(n8126), .IN3(n5837), .IN4(n5467), .QN(
        n5468) );
  OR4X1 U6927 ( .IN1(n5471), .IN2(n5470), .IN3(n5469), .IN4(n5468), .Q(
        \a6/N441 ) );
  NAND2X0 U6928 ( .IN1(n9080), .IN2(n5750), .QN(n7714) );
  NOR2X0 U6929 ( .IN1(n8645), .IN2(n7714), .QN(n7751) );
  INVX0 U6930 ( .INP(n8955), .ZN(n5901) );
  NOR2X0 U6931 ( .IN1(n7463), .IN2(n5901), .QN(n7677) );
  INVX0 U6932 ( .INP(n8240), .ZN(n6833) );
  NOR2X0 U6933 ( .IN1(n7347), .IN2(n6833), .QN(n7561) );
  NOR4X0 U6934 ( .IN1(n6487), .IN2(n7751), .IN3(n7677), .IN4(n7561), .QN(n5481) );
  AOI22X1 U6935 ( .IN1(n5472), .IN2(n7359), .IN3(n6207), .IN4(n8197), .QN(
        n5480) );
  INVX0 U6936 ( .INP(n6148), .ZN(n5823) );
  OA22X1 U6937 ( .IN1(n8171), .IN2(n7011), .IN3(n5823), .IN4(n7405), .Q(n5479)
         );
  NAND2X0 U6938 ( .IN1(n5473), .IN2(n7843), .QN(n7922) );
  INVX0 U6939 ( .INP(n7922), .ZN(n5984) );
  NOR2X0 U6940 ( .IN1(n7169), .IN2(n5474), .QN(n5476) );
  NAND2X0 U6941 ( .IN1(n8000), .IN2(n8875), .QN(n7729) );
  NAND2X0 U6942 ( .IN1(n9440), .IN2(n9181), .QN(n9045) );
  NOR2X0 U6943 ( .IN1(degrees_tmp2[3]), .IN2(n9045), .QN(n6507) );
  NAND2X0 U6944 ( .IN1(n7699), .IN2(n6507), .QN(n7376) );
  NOR2X0 U6945 ( .IN1(n7233), .IN2(n6120), .QN(n7254) );
  NAND2X0 U6946 ( .IN1(n8675), .IN2(n7254), .QN(n6442) );
  NAND3X0 U6947 ( .IN1(n7729), .IN2(n7376), .IN3(n6442), .QN(n5475) );
  NOR4X0 U6948 ( .IN1(n5984), .IN2(n5477), .IN3(n5476), .IN4(n5475), .QN(n5478) );
  NAND4X0 U6949 ( .IN1(n5481), .IN2(n5480), .IN3(n5479), .IN4(n5478), .QN(
        \a6/N442 ) );
  INVX0 U6950 ( .INP(n6967), .ZN(n5816) );
  NAND2X0 U6951 ( .IN1(n5816), .IN2(n9019), .QN(n8192) );
  INVX0 U6952 ( .INP(n9183), .ZN(n7164) );
  NAND2X0 U6953 ( .IN1(n8988), .IN2(n7164), .QN(n8164) );
  OA22X1 U6954 ( .IN1(n9440), .IN2(n8192), .IN3(n9438), .IN4(n8164), .Q(n5487)
         );
  NOR2X0 U6955 ( .IN1(n9435), .IN2(n8705), .QN(n9171) );
  NOR2X0 U6956 ( .IN1(degrees_tmp2[0]), .IN2(n8882), .QN(n9154) );
  NOR2X0 U6957 ( .IN1(n9171), .IN2(n9154), .QN(n6134) );
  OA22X1 U6958 ( .IN1(n8796), .IN2(n6238), .IN3(n6650), .IN4(n7293), .Q(n5486)
         );
  NAND2X0 U6959 ( .IN1(n9080), .IN2(n6637), .QN(n6312) );
  NAND2X0 U6960 ( .IN1(n6100), .IN2(n9166), .QN(n6975) );
  NAND3X0 U6961 ( .IN1(n6312), .IN2(n7485), .IN3(n6975), .QN(n5484) );
  NAND2X0 U6962 ( .IN1(n9434), .IN2(n9203), .QN(n6574) );
  INVX0 U6963 ( .INP(n6574), .ZN(n5547) );
  NAND2X0 U6964 ( .IN1(n8000), .IN2(n5547), .QN(n7862) );
  NAND3X0 U6965 ( .IN1(n5965), .IN2(n6758), .IN3(n9442), .QN(n7716) );
  NAND2X0 U6966 ( .IN1(n7862), .IN2(n7716), .QN(n6587) );
  NOR2X0 U6967 ( .IN1(n7416), .IN2(n8724), .QN(n9123) );
  NOR2X0 U6968 ( .IN1(n5538), .IN2(n5482), .QN(n7521) );
  AO22X1 U6969 ( .IN1(n8575), .IN2(n9123), .IN3(n8667), .IN4(n7521), .Q(n5483)
         );
  NOR4X0 U6970 ( .IN1(n6983), .IN2(n5484), .IN3(n6587), .IN4(n5483), .QN(n5485) );
  NAND4X0 U6971 ( .IN1(n5487), .IN2(n6134), .IN3(n5486), .IN4(n5485), .QN(
        \a6/N443 ) );
  NAND2X0 U6972 ( .IN1(n6182), .IN2(n9032), .QN(n6323) );
  NOR2X0 U6973 ( .IN1(n5488), .IN2(n6323), .QN(n6475) );
  NOR2X0 U6974 ( .IN1(n8461), .IN2(n8386), .QN(n9164) );
  AND2X1 U6975 ( .IN1(n9164), .IN2(n9445), .Q(n7898) );
  NAND2X0 U6976 ( .IN1(n8710), .IN2(n5931), .QN(n8452) );
  INVX0 U6977 ( .INP(n7291), .ZN(n7428) );
  NAND2X0 U6978 ( .IN1(n7428), .IN2(n6434), .QN(n8068) );
  NAND2X0 U6979 ( .IN1(n8475), .IN2(n9445), .QN(n8571) );
  NAND3X0 U6980 ( .IN1(n8452), .IN2(n8068), .IN3(n8571), .QN(n5491) );
  NAND2X0 U6981 ( .IN1(n7745), .IN2(n9122), .QN(n9155) );
  NAND2X0 U6982 ( .IN1(n5547), .IN2(n9155), .QN(n5489) );
  NOR2X0 U6983 ( .IN1(degrees_tmp2[3]), .IN2(n7416), .QN(n7501) );
  NAND2X0 U6984 ( .IN1(n7501), .IN2(n9019), .QN(n5500) );
  NAND3X0 U6985 ( .IN1(n5489), .IN2(n5500), .IN3(n6975), .QN(n5490) );
  NOR4X0 U6986 ( .IN1(n6475), .IN2(n7898), .IN3(n5491), .IN4(n5490), .QN(n5492) );
  INVX0 U6987 ( .INP(n8869), .ZN(n5640) );
  NAND2X0 U6988 ( .IN1(n5640), .IN2(n8282), .QN(n6534) );
  NAND4X0 U6989 ( .IN1(n5492), .IN2(n9088), .IN3(n6534), .IN4(n7616), .QN(
        \a6/N444 ) );
  NOR2X0 U6990 ( .IN1(degrees_tmp2[0]), .IN2(n7656), .QN(n6736) );
  NAND2X0 U6991 ( .IN1(n6173), .IN2(n6736), .QN(n5556) );
  INVX0 U6992 ( .INP(n6947), .ZN(n5493) );
  OA22X1 U6993 ( .IN1(n9441), .IN2(n5556), .IN3(n8317), .IN4(n5493), .Q(n5499)
         );
  NOR2X0 U6994 ( .IN1(degrees_tmp2[3]), .IN2(n6959), .QN(n8436) );
  NOR2X0 U6995 ( .IN1(n7876), .IN2(n7760), .QN(n6771) );
  NAND2X0 U6996 ( .IN1(n6623), .IN2(n8511), .QN(n8979) );
  NOR2X0 U6997 ( .IN1(n7736), .IN2(n8979), .QN(n6451) );
  NOR2X0 U6998 ( .IN1(n8041), .IN2(n8268), .QN(n8942) );
  OR2X1 U6999 ( .IN1(n8005), .IN2(n8942), .Q(n8773) );
  NOR4X0 U7000 ( .IN1(n8436), .IN2(n6771), .IN3(n6451), .IN4(n8773), .QN(n5497) );
  NOR2X0 U7001 ( .IN1(n5494), .IN2(n6320), .QN(n5495) );
  OA22X1 U7002 ( .IN1(n8796), .IN2(n8705), .IN3(n8667), .IN4(n5495), .Q(n5496)
         );
  NOR2X0 U7003 ( .IN1(n8213), .IN2(n6369), .QN(n5716) );
  NAND2X0 U7004 ( .IN1(n8752), .IN2(n5716), .QN(n8200) );
  AND4X1 U7005 ( .IN1(n5497), .IN2(n5496), .IN3(n8891), .IN4(n8200), .Q(n5498)
         );
  NAND4X0 U7006 ( .IN1(n5499), .IN2(n5498), .IN3(n5897), .IN4(n7834), .QN(
        \a6/N445 ) );
  NOR2X0 U7007 ( .IN1(n9445), .IN2(n8880), .QN(n7850) );
  OA21X1 U7008 ( .IN1(n6261), .IN2(n9184), .IN3(n9037), .Q(n5504) );
  NOR2X0 U7009 ( .IN1(n6651), .IN2(n7969), .QN(n6034) );
  NAND2X0 U7010 ( .IN1(n6034), .IN2(n9438), .QN(n7294) );
  OA22X1 U7011 ( .IN1(n9054), .IN2(n6308), .IN3(n8188), .IN4(n7294), .Q(n5502)
         );
  INVX0 U7012 ( .INP(n7405), .ZN(n8847) );
  NAND2X0 U7013 ( .IN1(n8752), .IN2(n9203), .QN(n7009) );
  OA22X1 U7014 ( .IN1(n8667), .IN2(n7404), .IN3(n8847), .IN4(n7009), .Q(n5501)
         );
  NAND2X0 U7015 ( .IN1(n7033), .IN2(n8041), .QN(n8590) );
  NAND4X0 U7016 ( .IN1(n5502), .IN2(n5501), .IN3(n5500), .IN4(n8590), .QN(
        n5503) );
  NOR4X0 U7017 ( .IN1(n7518), .IN2(n7850), .IN3(n5504), .IN4(n5503), .QN(n5506) );
  NAND2X0 U7018 ( .IN1(n9190), .IN2(n9084), .QN(n7647) );
  AO21X1 U7019 ( .IN1(n8268), .IN2(n8684), .IN3(n8333), .Q(n5505) );
  NAND4X0 U7020 ( .IN1(n5506), .IN2(n7025), .IN3(n7647), .IN4(n5505), .QN(
        \a6/N446 ) );
  OA22X1 U7021 ( .IN1(n7597), .IN2(n9020), .IN3(n8169), .IN4(n6804), .Q(n5515)
         );
  NOR2X0 U7022 ( .IN1(n8649), .IN2(n7647), .QN(n7907) );
  NOR2X0 U7023 ( .IN1(n8531), .IN2(n8527), .QN(n6640) );
  OA21X1 U7024 ( .IN1(n9033), .IN2(n7582), .IN3(n8188), .Q(n5512) );
  NAND2X0 U7025 ( .IN1(n9435), .IN2(n8567), .QN(n8024) );
  NAND2X0 U7026 ( .IN1(n8247), .IN2(n9442), .QN(n5507) );
  OA22X1 U7027 ( .IN1(n8978), .IN2(n8024), .IN3(n5507), .IN4(n8684), .Q(n5510)
         );
  INVX0 U7028 ( .INP(n5708), .ZN(n8782) );
  NAND2X0 U7029 ( .IN1(n7736), .IN2(n8782), .QN(n6863) );
  NAND2X0 U7030 ( .IN1(n7032), .IN2(n6863), .QN(n6500) );
  AO21X1 U7031 ( .IN1(n8043), .IN2(n6500), .IN3(n9434), .Q(n5509) );
  INVX0 U7032 ( .INP(n9155), .ZN(n9131) );
  NOR2X0 U7033 ( .IN1(degrees_tmp2[0]), .IN2(n9131), .QN(n6755) );
  NAND2X0 U7034 ( .IN1(n8186), .IN2(n6755), .QN(n5508) );
  NAND4X0 U7035 ( .IN1(n5510), .IN2(n5509), .IN3(n5520), .IN4(n5508), .QN(
        n5511) );
  NOR4X0 U7036 ( .IN1(n7907), .IN2(n6640), .IN3(n5512), .IN4(n5511), .QN(n5514) );
  NAND2X0 U7037 ( .IN1(n8816), .IN2(n9164), .QN(n6413) );
  NAND2X0 U7038 ( .IN1(degrees_tmp2[0]), .IN2(n8675), .QN(n7143) );
  NAND2X0 U7039 ( .IN1(n8229), .IN2(n7143), .QN(n6085) );
  NAND2X0 U7040 ( .IN1(n6637), .IN2(n6085), .QN(n5513) );
  NAND4X0 U7041 ( .IN1(n5515), .IN2(n5514), .IN3(n6413), .IN4(n5513), .QN(
        \a6/N447 ) );
  AND2X1 U7042 ( .IN1(n7111), .IN2(n9041), .Q(n5954) );
  NOR2X0 U7043 ( .IN1(n6194), .IN2(n5516), .QN(n8881) );
  NAND2X0 U7044 ( .IN1(n6119), .IN2(n6493), .QN(n7251) );
  OA22X1 U7045 ( .IN1(n8881), .IN2(n7876), .IN3(n6369), .IN4(n7251), .Q(n5522)
         );
  NOR2X0 U7046 ( .IN1(n7437), .IN2(n9119), .QN(n5518) );
  NOR2X0 U7047 ( .IN1(n6371), .IN2(n8001), .QN(n6448) );
  NAND2X0 U7048 ( .IN1(n9202), .IN2(n6797), .QN(n8218) );
  INVX0 U7049 ( .INP(n6635), .ZN(n6268) );
  NAND2X0 U7050 ( .IN1(n6268), .IN2(n5547), .QN(n6524) );
  NAND4X0 U7051 ( .IN1(n8218), .IN2(n7838), .IN3(n7099), .IN4(n6524), .QN(
        n5517) );
  NOR4X0 U7052 ( .IN1(n5518), .IN2(n6448), .IN3(n6914), .IN4(n5517), .QN(n5519) );
  OA221X1 U7053 ( .IN1(n9433), .IN2(n6835), .IN3(n9433), .IN4(n5520), .IN5(
        n5519), .Q(n5521) );
  NAND2X0 U7054 ( .IN1(n5913), .IN2(n9442), .QN(n6426) );
  NOR2X0 U7055 ( .IN1(n9437), .IN2(n6426), .QN(n7669) );
  NAND2X0 U7056 ( .IN1(n8883), .IN2(n7669), .QN(n7010) );
  NAND4X0 U7057 ( .IN1(n5954), .IN2(n5522), .IN3(n5521), .IN4(n7010), .QN(
        \a6/N448 ) );
  NOR2X0 U7058 ( .IN1(n8386), .IN2(n8595), .QN(n6124) );
  NAND2X0 U7059 ( .IN1(n8467), .IN2(n6124), .QN(n8906) );
  NOR2X0 U7060 ( .IN1(n7347), .IN2(n8588), .QN(n8654) );
  NAND2X0 U7061 ( .IN1(n8654), .IN2(n9440), .QN(n8364) );
  NAND2X0 U7062 ( .IN1(n8424), .IN2(n6623), .QN(n8801) );
  INVX0 U7063 ( .INP(n8801), .ZN(n7487) );
  NAND2X0 U7064 ( .IN1(degrees_tmp2[5]), .IN2(n7487), .QN(n8055) );
  NAND2X0 U7065 ( .IN1(n8424), .IN2(n8163), .QN(n7165) );
  NAND4X0 U7066 ( .IN1(n8906), .IN2(n8364), .IN3(n8055), .IN4(n7165), .QN(
        n5526) );
  NOR2X0 U7067 ( .IN1(n8883), .IN2(n9073), .QN(n6257) );
  OA22X1 U7068 ( .IN1(n8598), .IN2(n8244), .IN3(n6257), .IN4(n7393), .Q(n5524)
         );
  NAND2X0 U7069 ( .IN1(n9435), .IN2(n8731), .QN(n6728) );
  INVX0 U7070 ( .INP(n6296), .ZN(n7340) );
  OA22X1 U7071 ( .IN1(n6182), .IN2(n6728), .IN3(n9045), .IN4(n7340), .Q(n5523)
         );
  INVX0 U7072 ( .INP(n8310), .ZN(n9200) );
  NAND4X0 U7073 ( .IN1(n5524), .IN2(n5523), .IN3(n9030), .IN4(n9200), .QN(
        n5525) );
  NOR2X0 U7074 ( .IN1(n5526), .IN2(n5525), .QN(n5528) );
  INVX0 U7075 ( .INP(n5722), .ZN(n9067) );
  NAND2X0 U7076 ( .IN1(n8180), .IN2(n6736), .QN(n5607) );
  NAND4X0 U7077 ( .IN1(n5528), .IN2(n9067), .IN3(n5527), .IN4(n5607), .QN(
        \a6/N449 ) );
  NAND2X0 U7078 ( .IN1(n9076), .IN2(n9442), .QN(n8193) );
  INVX0 U7079 ( .INP(n8193), .ZN(n7652) );
  NOR2X0 U7080 ( .IN1(n6919), .IN2(n8317), .QN(n5869) );
  NOR2X0 U7081 ( .IN1(n7652), .IN2(n5869), .QN(n7153) );
  NOR2X0 U7082 ( .IN1(n8597), .IN2(n9023), .QN(n5534) );
  INVX0 U7083 ( .INP(n7954), .ZN(n8655) );
  NAND2X0 U7084 ( .IN1(n6650), .IN2(n8655), .QN(n8701) );
  NAND2X0 U7085 ( .IN1(n8247), .IN2(n5971), .QN(n7773) );
  NAND4X0 U7086 ( .IN1(n7729), .IN2(n8846), .IN3(n8701), .IN4(n7773), .QN(
        n5531) );
  NOR2X0 U7087 ( .IN1(n7717), .IN2(n6967), .QN(n9176) );
  NAND2X0 U7088 ( .IN1(n8995), .IN2(n9176), .QN(n6536) );
  NAND2X0 U7089 ( .IN1(n8723), .IN2(n9149), .QN(n8808) );
  NAND2X0 U7090 ( .IN1(n5529), .IN2(n8760), .QN(n8962) );
  NOR2X0 U7091 ( .IN1(n8531), .IN2(n8707), .QN(n6720) );
  NAND2X0 U7092 ( .IN1(n6720), .IN2(n9445), .QN(n6072) );
  NAND4X0 U7093 ( .IN1(n6536), .IN2(n8808), .IN3(n8962), .IN4(n6072), .QN(
        n5530) );
  NOR2X0 U7094 ( .IN1(n5531), .IN2(n5530), .QN(n5532) );
  NAND3X0 U7095 ( .IN1(degrees_tmp2[0]), .IN2(n9435), .IN3(n8408), .QN(n8892)
         );
  NAND2X0 U7096 ( .IN1(n5532), .IN2(n8892), .QN(n5533) );
  NOR2X0 U7097 ( .IN1(n5534), .IN2(n5533), .QN(n5537) );
  NAND2X0 U7098 ( .IN1(n5843), .IN2(n7405), .QN(n5535) );
  NAND4X0 U7099 ( .IN1(n7153), .IN2(n5537), .IN3(n5536), .IN4(n5535), .QN(
        \a6/N450 ) );
  INVX0 U7100 ( .INP(n6238), .ZN(n6416) );
  AO22X1 U7101 ( .IN1(n8519), .IN2(n8645), .IN3(n8567), .IN4(n8531), .Q(n5542)
         );
  NOR2X0 U7102 ( .IN1(n8529), .IN2(n7936), .QN(n8772) );
  INVX0 U7103 ( .INP(n7700), .ZN(n5795) );
  OA22X1 U7104 ( .IN1(n8772), .IN2(n5795), .IN3(n9197), .IN4(n9003), .Q(n5540)
         );
  NAND2X0 U7105 ( .IN1(n5538), .IN2(n6401), .QN(n8034) );
  INVX0 U7106 ( .INP(n8034), .ZN(n7613) );
  NAND2X0 U7107 ( .IN1(n5832), .IN2(n8816), .QN(n6553) );
  OA21X1 U7108 ( .IN1(n7613), .IN2(n6553), .IN3(n7099), .Q(n5539) );
  INVX0 U7109 ( .INP(n6640), .ZN(n7861) );
  NAND4X0 U7110 ( .IN1(n5540), .IN2(n5539), .IN3(n7495), .IN4(n7861), .QN(
        n5541) );
  NOR4X0 U7111 ( .IN1(n6416), .IN2(n7678), .IN3(n5542), .IN4(n5541), .QN(n5544) );
  INVX0 U7112 ( .INP(n7827), .ZN(n5667) );
  NAND3X0 U7113 ( .IN1(n8249), .IN2(n6758), .IN3(n9166), .QN(n5543) );
  NAND4X0 U7114 ( .IN1(n5544), .IN2(n5667), .IN3(n8563), .IN4(n5543), .QN(
        \a6/N451 ) );
  NAND2X0 U7115 ( .IN1(n5545), .IN2(n5913), .QN(n5768) );
  INVX0 U7116 ( .INP(n5768), .ZN(n6942) );
  NOR2X0 U7117 ( .IN1(n6942), .IN2(n9202), .QN(n5546) );
  NAND3X0 U7118 ( .IN1(degrees_tmp2[5]), .IN2(n9190), .IN3(n9436), .QN(n8276)
         );
  OA22X1 U7119 ( .IN1(n5546), .IN2(n9155), .IN3(n9048), .IN4(n8276), .Q(n5552)
         );
  INVX0 U7120 ( .INP(n9122), .ZN(n8533) );
  INVX0 U7121 ( .INP(n6085), .ZN(n7058) );
  OA22X1 U7122 ( .IN1(n8533), .IN2(n8438), .IN3(n7058), .IN4(n5624), .Q(n5551)
         );
  NOR2X0 U7123 ( .IN1(n7534), .IN2(n6836), .QN(n8982) );
  INVX0 U7124 ( .INP(n8982), .ZN(n8522) );
  NAND2X0 U7125 ( .IN1(n5547), .IN2(n9209), .QN(n6088) );
  NAND2X0 U7126 ( .IN1(n8529), .IN2(n9023), .QN(n5853) );
  AND4X1 U7127 ( .IN1(n8522), .IN2(n8571), .IN3(n6088), .IN4(n5853), .Q(n5549)
         );
  NAND2X0 U7128 ( .IN1(n8180), .IN2(n8710), .QN(n8748) );
  NAND2X0 U7129 ( .IN1(n8534), .IN2(n6067), .QN(n8966) );
  NAND3X0 U7130 ( .IN1(n8697), .IN2(n9436), .IN3(n7736), .QN(n5548) );
  AND4X1 U7131 ( .IN1(n5549), .IN2(n8748), .IN3(n8966), .IN4(n5548), .Q(n5550)
         );
  NOR2X0 U7132 ( .IN1(n8268), .IN2(n8282), .QN(n6974) );
  INVX0 U7133 ( .INP(n6974), .ZN(n7273) );
  NAND4X0 U7134 ( .IN1(n5552), .IN2(n5551), .IN3(n5550), .IN4(n7273), .QN(
        \a6/N452 ) );
  INVX0 U7135 ( .INP(n7518), .ZN(n8067) );
  NOR2X0 U7136 ( .IN1(n8649), .IN2(n8067), .QN(n7077) );
  NOR2X0 U7137 ( .IN1(n6651), .IN2(n5757), .QN(n7236) );
  NOR3X0 U7138 ( .IN1(n7236), .IN2(n5709), .IN3(n5553), .QN(n5554) );
  NOR2X0 U7139 ( .IN1(n5554), .IN2(n9061), .QN(n5559) );
  AOI22X1 U7140 ( .IN1(n8282), .IN2(n6668), .IN3(n8630), .IN4(n7843), .QN(
        n5555) );
  NAND2X0 U7141 ( .IN1(n9435), .IN2(n9076), .QN(n8426) );
  NAND4X0 U7142 ( .IN1(n9210), .IN2(degrees_tmp2[3]), .IN3(n8171), .IN4(n8630), 
        .QN(n6450) );
  NAND3X0 U7143 ( .IN1(n5555), .IN2(n8426), .IN3(n6450), .QN(n5558) );
  INVX0 U7144 ( .INP(n6448), .ZN(n8069) );
  NAND2X0 U7145 ( .IN1(n9033), .IN2(n9442), .QN(n8841) );
  NOR2X0 U7146 ( .IN1(degrees_tmp2[3]), .IN2(n8841), .QN(n7849) );
  NAND2X0 U7147 ( .IN1(n7849), .IN2(n9440), .QN(n7924) );
  NAND4X0 U7148 ( .IN1(n8846), .IN2(n5556), .IN3(n8069), .IN4(n7924), .QN(
        n5557) );
  NOR4X0 U7149 ( .IN1(n7077), .IN2(n5559), .IN3(n5558), .IN4(n5557), .QN(n5560) );
  NAND3X0 U7150 ( .IN1(n8186), .IN2(n8185), .IN3(n9442), .QN(n8633) );
  NAND4X0 U7151 ( .IN1(n5560), .IN2(n8748), .IN3(n8633), .IN4(n7738), .QN(
        \a6/N454 ) );
  NOR2X0 U7152 ( .IN1(n9434), .IN2(n6311), .QN(n8606) );
  NAND3X0 U7153 ( .IN1(n9435), .IN2(n6698), .IN3(n7784), .QN(n7475) );
  NOR2X0 U7154 ( .IN1(n9213), .IN2(n7035), .QN(n9075) );
  NAND2X0 U7155 ( .IN1(n9075), .IN2(n7945), .QN(n6950) );
  NAND2X0 U7156 ( .IN1(n7615), .IN2(n8640), .QN(n6254) );
  NAND4X0 U7157 ( .IN1(n7475), .IN2(n7446), .IN3(n6950), .IN4(n6254), .QN(
        n5568) );
  INVX0 U7158 ( .INP(n7989), .ZN(n6365) );
  NAND2X0 U7159 ( .IN1(n6365), .IN2(n7784), .QN(n8834) );
  NAND2X0 U7160 ( .IN1(n8533), .IN2(n9172), .QN(n8668) );
  AND2X1 U7161 ( .IN1(n8834), .IN2(n8668), .Q(n6818) );
  NAND2X0 U7162 ( .IN1(degrees_tmp2[2]), .IN2(n6417), .QN(n7465) );
  NOR2X0 U7163 ( .IN1(n8940), .IN2(n7465), .QN(n8144) );
  NAND2X0 U7164 ( .IN1(n8760), .IN2(n8144), .QN(n5562) );
  NAND3X0 U7165 ( .IN1(n9210), .IN2(n7179), .IN3(n8780), .QN(n5561) );
  NAND4X0 U7166 ( .IN1(n6818), .IN2(n6567), .IN3(n5562), .IN4(n5561), .QN(
        n5567) );
  NAND3X0 U7167 ( .IN1(n6100), .IN2(n7760), .IN3(n7233), .QN(n6402) );
  NOR2X0 U7168 ( .IN1(n9080), .IN2(n6243), .QN(n8321) );
  NAND2X0 U7169 ( .IN1(n9190), .IN2(n8198), .QN(n8859) );
  OA22X1 U7170 ( .IN1(n8321), .IN2(n8859), .IN3(n8171), .IN4(n7009), .Q(n5563)
         );
  OA21X1 U7171 ( .IN1(n9436), .IN2(n6402), .IN3(n5563), .Q(n5565) );
  NAND2X0 U7172 ( .IN1(n5716), .IN2(n9442), .QN(n7881) );
  NOR2X0 U7173 ( .IN1(n9441), .IN2(n7881), .QN(n5788) );
  INVX0 U7174 ( .INP(n5788), .ZN(n7018) );
  NAND2X0 U7175 ( .IN1(n7050), .IN2(n5913), .QN(n7538) );
  INVX0 U7176 ( .INP(n7538), .ZN(n7500) );
  NAND3X0 U7177 ( .IN1(degrees_tmp2[2]), .IN2(n7500), .IN3(n8282), .QN(n5564)
         );
  NAND4X0 U7178 ( .IN1(n5565), .IN2(n7018), .IN3(n8624), .IN4(n5564), .QN(
        n5566) );
  OR4X1 U7179 ( .IN1(n8606), .IN2(n5568), .IN3(n5567), .IN4(n5566), .Q(
        \a6/N455 ) );
  NOR2X0 U7180 ( .IN1(n8489), .IN2(n8729), .QN(n6901) );
  NOR2X0 U7181 ( .IN1(n8041), .IN2(n6634), .QN(n5569) );
  NOR2X0 U7182 ( .IN1(n6901), .IN2(n5569), .QN(n8644) );
  INVX0 U7183 ( .INP(n8131), .ZN(n8786) );
  INVX0 U7184 ( .INP(n8566), .ZN(n7004) );
  AOI21X1 U7185 ( .IN1(n7004), .IN2(n5615), .IN3(n9060), .QN(n5575) );
  NOR3X0 U7186 ( .IN1(degrees_tmp2[5]), .IN2(n8639), .IN3(n7566), .QN(n5574)
         );
  NOR2X0 U7187 ( .IN1(n7585), .IN2(n9435), .QN(n5571) );
  NAND2X0 U7188 ( .IN1(n6155), .IN2(n7784), .QN(n8905) );
  NAND2X0 U7189 ( .IN1(n8706), .IN2(n8905), .QN(n5570) );
  NOR2X0 U7190 ( .IN1(n5571), .IN2(n5570), .QN(n5572) );
  NOR2X0 U7191 ( .IN1(n9433), .IN2(n8004), .QN(n6699) );
  NAND2X0 U7192 ( .IN1(n8534), .IN2(n6699), .QN(n7998) );
  NAND4X0 U7193 ( .IN1(n5572), .IN2(n7998), .IN3(n8892), .IN4(n9058), .QN(
        n5573) );
  NOR4X0 U7194 ( .IN1(n8786), .IN2(n5575), .IN3(n5574), .IN4(n5573), .QN(n5576) );
  NAND4X0 U7195 ( .IN1(n8644), .IN2(n5576), .IN3(n7308), .IN4(n8701), .QN(
        \a6/N456 ) );
  INVX0 U7196 ( .INP(n9075), .ZN(n8708) );
  OA22X1 U7197 ( .IN1(n9082), .IN2(n7011), .IN3(n8710), .IN4(n8708), .Q(n5583)
         );
  NAND2X0 U7198 ( .IN1(n7195), .IN2(n8883), .QN(n7721) );
  NAND4X0 U7199 ( .IN1(n8817), .IN2(n9178), .IN3(n7721), .IN4(n6786), .QN(
        n5581) );
  NOR2X0 U7200 ( .IN1(n8282), .IN2(n7288), .QN(n5578) );
  NAND2X0 U7201 ( .IN1(n5931), .IN2(n6017), .QN(n8100) );
  NAND2X0 U7202 ( .IN1(n8840), .IN2(n8100), .QN(n5577) );
  NOR2X0 U7203 ( .IN1(n5578), .IN2(n5577), .QN(n5579) );
  NAND2X0 U7204 ( .IN1(n9183), .IN2(n5949), .QN(n8316) );
  NAND3X0 U7205 ( .IN1(n9437), .IN2(n8188), .IN3(n6697), .QN(n5742) );
  NAND4X0 U7206 ( .IN1(n5579), .IN2(n8316), .IN3(n8156), .IN4(n5742), .QN(
        n5580) );
  NOR4X0 U7207 ( .IN1(n7077), .IN2(n8855), .IN3(n5581), .IN4(n5580), .QN(n5582) );
  NAND2X0 U7208 ( .IN1(n5673), .IN2(n8282), .QN(n8049) );
  INVX0 U7209 ( .INP(n7875), .ZN(n8948) );
  NAND2X0 U7210 ( .IN1(n8188), .IN2(n8948), .QN(n6305) );
  NAND4X0 U7211 ( .IN1(n5583), .IN2(n5582), .IN3(n8049), .IN4(n6305), .QN(
        \a6/N457 ) );
  NAND2X0 U7212 ( .IN1(n8119), .IN2(n5936), .QN(n6823) );
  INVX0 U7213 ( .INP(n6823), .ZN(n6086) );
  NAND2X0 U7214 ( .IN1(n6086), .IN2(n7784), .QN(n8819) );
  NOR2X0 U7215 ( .IN1(n9440), .IN2(n8819), .QN(n7408) );
  NOR2X0 U7216 ( .IN1(n9438), .IN2(n8578), .QN(n7972) );
  AO22X1 U7217 ( .IN1(n7032), .IN2(n8484), .IN3(n7972), .IN4(n7800), .Q(n5587)
         );
  NAND2X0 U7218 ( .IN1(n6392), .IN2(n6136), .QN(n8514) );
  OA21X1 U7219 ( .IN1(n7184), .IN2(n7721), .IN3(n8514), .Q(n5585) );
  NOR2X0 U7220 ( .IN1(n9435), .IN2(n7168), .QN(n7142) );
  NAND2X0 U7221 ( .IN1(n7142), .IN2(n9436), .QN(n6142) );
  NAND2X0 U7222 ( .IN1(n9182), .IN2(n9080), .QN(n6591) );
  INVX0 U7223 ( .INP(n7378), .ZN(n6055) );
  NOR2X0 U7224 ( .IN1(n6055), .IN2(n8179), .QN(n8211) );
  OA221X1 U7225 ( .IN1(degrees_tmp2[3]), .IN2(n6142), .IN3(degrees_tmp2[3]), 
        .IN4(n6591), .IN5(n8211), .Q(n5584) );
  NAND2X0 U7226 ( .IN1(n7517), .IN2(n6124), .QN(n7082) );
  NAND4X0 U7227 ( .IN1(n5585), .IN2(n5584), .IN3(n6312), .IN4(n7082), .QN(
        n5586) );
  NOR4X0 U7228 ( .IN1(n5606), .IN2(n7408), .IN3(n5587), .IN4(n5586), .QN(n5590) );
  NOR2X0 U7229 ( .IN1(n5588), .IN2(n6574), .QN(n5876) );
  INVX0 U7230 ( .INP(n5876), .ZN(n7943) );
  NAND3X0 U7231 ( .IN1(degrees_tmp2[5]), .IN2(n8163), .IN3(n8947), .QN(n5589)
         );
  NAND4X0 U7232 ( .IN1(n5590), .IN2(n7940), .IN3(n7943), .IN4(n5589), .QN(
        \a6/N458 ) );
  NOR2X0 U7233 ( .IN1(n7686), .IN2(n7649), .QN(n8985) );
  NOR2X0 U7234 ( .IN1(n5788), .IN2(n8985), .QN(n8082) );
  NAND2X0 U7235 ( .IN1(n8186), .IN2(n9440), .QN(n8294) );
  NOR2X0 U7236 ( .IN1(n9188), .IN2(n8468), .QN(n5591) );
  OA22X1 U7237 ( .IN1(n8752), .IN2(n8294), .IN3(n5591), .IN4(n7686), .Q(n5598)
         );
  NAND2X0 U7238 ( .IN1(n8188), .IN2(n6449), .QN(n7245) );
  NAND4X0 U7239 ( .IN1(n6312), .IN2(n7730), .IN3(n8668), .IN4(n7245), .QN(
        n5595) );
  OA22X1 U7240 ( .IN1(n9205), .IN2(n6833), .IN3(n7954), .IN4(n7914), .Q(n5593)
         );
  NAND2X0 U7241 ( .IN1(n8883), .IN2(n6637), .QN(n6131) );
  NAND2X0 U7242 ( .IN1(n9105), .IN2(n6699), .QN(n7118) );
  NAND2X0 U7243 ( .IN1(n8534), .IN2(n7438), .QN(n5592) );
  NAND4X0 U7244 ( .IN1(n5593), .IN2(n6131), .IN3(n7118), .IN4(n5592), .QN(
        n5594) );
  NOR2X0 U7245 ( .IN1(n5595), .IN2(n5594), .QN(n5597) );
  INVX0 U7246 ( .INP(n7873), .ZN(n7728) );
  NAND2X0 U7247 ( .IN1(n7728), .IN2(n9433), .QN(n7519) );
  AO21X1 U7248 ( .IN1(n6286), .IN2(n7519), .IN3(n9073), .Q(n5596) );
  NAND4X0 U7249 ( .IN1(n8082), .IN2(n5598), .IN3(n5597), .IN4(n5596), .QN(
        \a6/N460 ) );
  NOR2X0 U7250 ( .IN1(n8240), .IN2(n9073), .QN(n7895) );
  OA22X1 U7251 ( .IN1(n7895), .IN2(n6832), .IN3(n7402), .IN4(n8979), .Q(n5605)
         );
  NAND2X0 U7252 ( .IN1(n9190), .IN2(n8188), .QN(n7608) );
  NOR2X0 U7253 ( .IN1(n9436), .IN2(n7608), .QN(n7727) );
  OA21X1 U7254 ( .IN1(n6086), .IN2(n8640), .IN3(n7169), .Q(n5603) );
  NOR2X0 U7255 ( .IN1(n9440), .IN2(n6205), .QN(n6504) );
  NOR2X0 U7256 ( .IN1(n6504), .IN2(n7358), .QN(n7926) );
  OR2X1 U7257 ( .IN1(n7926), .IN2(n9445), .Q(n5601) );
  NAND2X0 U7258 ( .IN1(n8890), .IN2(n6756), .QN(n6903) );
  INVX0 U7259 ( .INP(n9202), .ZN(n6568) );
  NAND3X0 U7260 ( .IN1(n6568), .IN2(n8268), .IN3(n8495), .QN(n5599) );
  NAND2X0 U7261 ( .IN1(n5599), .IN2(n9082), .QN(n5600) );
  NAND4X0 U7262 ( .IN1(n8135), .IN2(n5601), .IN3(n6903), .IN4(n5600), .QN(
        n5602) );
  NOR4X0 U7263 ( .IN1(n6771), .IN2(n7727), .IN3(n5603), .IN4(n5602), .QN(n5604) );
  INVX0 U7264 ( .INP(n6283), .ZN(n8226) );
  NAND4X0 U7265 ( .IN1(n5605), .IN2(n5604), .IN3(n8167), .IN4(n8226), .QN(
        \a6/N461 ) );
  NOR2X0 U7266 ( .IN1(n9435), .IN2(n8438), .QN(n7412) );
  NOR3X0 U7267 ( .IN1(n7077), .IN2(n5606), .IN3(n7412), .QN(n5614) );
  NAND2X0 U7268 ( .IN1(n8000), .IN2(n9190), .QN(n8453) );
  OA22X1 U7269 ( .IN1(n9031), .IN2(n8453), .IN3(n7800), .IN4(n6337), .Q(n5613)
         );
  NAND2X0 U7270 ( .IN1(n8572), .IN2(n8823), .QN(n8743) );
  NAND4X0 U7271 ( .IN1(n8891), .IN2(n8069), .IN3(n6903), .IN4(n8743), .QN(
        n5611) );
  OA22X1 U7272 ( .IN1(n8796), .IN2(n5607), .IN3(n8978), .IN4(n8592), .Q(n5609)
         );
  NAND2X0 U7273 ( .IN1(degrees_tmp2[0]), .IN2(n6220), .QN(n5608) );
  NAND3X0 U7274 ( .IN1(n6620), .IN2(n9437), .IN3(n7597), .QN(n6188) );
  NAND4X0 U7275 ( .IN1(n5609), .IN2(n7981), .IN3(n5608), .IN4(n6188), .QN(
        n5610) );
  NOR4X0 U7276 ( .IN1(n6896), .IN2(n6213), .IN3(n5611), .IN4(n5610), .QN(n5612) );
  NAND4X0 U7277 ( .IN1(n5614), .IN2(n5613), .IN3(n5612), .IN4(n7764), .QN(
        \a6/N462 ) );
  NAND2X0 U7278 ( .IN1(n5757), .IN2(n6921), .QN(n8494) );
  OA22X1 U7279 ( .IN1(n9023), .IN2(n8550), .IN3(n8494), .IN4(n8578), .Q(n5622)
         );
  NOR2X0 U7280 ( .IN1(n7808), .IN2(n6322), .QN(n7281) );
  INVX0 U7281 ( .INP(n7281), .ZN(n6727) );
  NOR2X0 U7282 ( .IN1(n8431), .IN2(n6727), .QN(n7374) );
  AND3X1 U7283 ( .IN1(n8875), .IN2(n9433), .IN3(n8787), .Q(n7434) );
  NOR2X0 U7284 ( .IN1(n5615), .IN2(n6836), .QN(n5619) );
  NOR2X0 U7285 ( .IN1(n8001), .IN2(n5616), .QN(n8287) );
  INVX0 U7286 ( .INP(n8287), .ZN(n8689) );
  INVX0 U7287 ( .INP(n7552), .ZN(n6214) );
  NAND2X0 U7288 ( .IN1(n6214), .IN2(n6173), .QN(n7824) );
  NOR2X0 U7289 ( .IN1(n6649), .IN2(n6699), .QN(n7424) );
  NAND2X0 U7290 ( .IN1(n8220), .IN2(n8890), .QN(n6059) );
  OR2X1 U7291 ( .IN1(n7424), .IN2(n6059), .Q(n8388) );
  NOR2X0 U7292 ( .IN1(n8883), .IN2(n9080), .QN(n6895) );
  NAND3X0 U7293 ( .IN1(n6698), .IN2(n9183), .IN3(n6895), .QN(n5617) );
  NAND4X0 U7294 ( .IN1(n8689), .IN2(n7824), .IN3(n8388), .IN4(n5617), .QN(
        n5618) );
  NOR4X0 U7295 ( .IN1(n7374), .IN2(n7434), .IN3(n5619), .IN4(n5618), .QN(n5621) );
  NAND2X0 U7296 ( .IN1(n7582), .IN2(n9433), .QN(n7812) );
  INVX0 U7297 ( .INP(n9027), .ZN(n5620) );
  NAND2X0 U7298 ( .IN1(n5620), .IN2(n7841), .QN(n7785) );
  NAND4X0 U7299 ( .IN1(n5622), .IN2(n5621), .IN3(n7812), .IN4(n7785), .QN(
        \a6/N463 ) );
  NOR2X0 U7300 ( .IN1(n8692), .IN2(n8597), .QN(n9065) );
  NOR2X0 U7301 ( .IN1(n5624), .IN2(n5623), .QN(n7788) );
  NOR3X0 U7302 ( .IN1(n9065), .IN2(n8982), .IN3(n7788), .QN(n8363) );
  NAND3X0 U7303 ( .IN1(n8363), .IN2(n7010), .IN3(n8214), .QN(n5631) );
  INVX0 U7304 ( .INP(n6308), .ZN(n9025) );
  NAND2X0 U7305 ( .IN1(n9025), .IN2(n8947), .QN(n5625) );
  NAND2X0 U7306 ( .IN1(n8728), .IN2(n6296), .QN(n8236) );
  NAND3X0 U7307 ( .IN1(degrees_tmp2[3]), .IN2(n7184), .IN3(n7582), .QN(n6767)
         );
  NAND4X0 U7308 ( .IN1(n6135), .IN2(n5625), .IN3(n8236), .IN4(n6767), .QN(
        n5630) );
  OA22X1 U7309 ( .IN1(n9054), .IN2(n9003), .IN3(n6836), .IN4(n8761), .Q(n5628)
         );
  NAND2X0 U7310 ( .IN1(n5626), .IN2(n7213), .QN(n5627) );
  NAND4X0 U7311 ( .IN1(n5628), .IN2(n5646), .IN3(n7981), .IN4(n5627), .QN(
        n5629) );
  OR4X1 U7312 ( .IN1(n6034), .IN2(n5631), .IN3(n5630), .IN4(n5629), .Q(
        \a6/N464 ) );
  OA22X1 U7313 ( .IN1(n9445), .IN2(n7608), .IN3(n7035), .IN4(n5632), .Q(n5639)
         );
  NOR2X0 U7314 ( .IN1(degrees_tmp2[2]), .IN2(n7011), .QN(n6541) );
  AND3X1 U7315 ( .IN1(n6637), .IN2(n9440), .IN3(n8947), .Q(n5637) );
  NAND2X0 U7316 ( .IN1(n8447), .IN2(n7760), .QN(n5844) );
  OA22X1 U7317 ( .IN1(n8876), .IN2(n7510), .IN3(n6464), .IN4(n9155), .Q(n5633)
         );
  OA221X1 U7318 ( .IN1(n6919), .IN2(n7679), .IN3(n6919), .IN4(n5844), .IN5(
        n5633), .Q(n5635) );
  NAND2X0 U7319 ( .IN1(n8675), .IN2(n5761), .QN(n7953) );
  OA22X1 U7320 ( .IN1(n8816), .IN2(n7548), .IN3(n7953), .IN4(n7233), .Q(n5634)
         );
  NAND3X0 U7321 ( .IN1(n8188), .IN2(n8163), .IN3(n9440), .QN(n7771) );
  INVX0 U7322 ( .INP(n7908), .ZN(n8765) );
  NAND4X0 U7323 ( .IN1(n5635), .IN2(n5634), .IN3(n7771), .IN4(n8765), .QN(
        n5636) );
  NOR4X0 U7324 ( .IN1(n6541), .IN2(n8723), .IN3(n5637), .IN4(n5636), .QN(n5638) );
  NAND2X0 U7325 ( .IN1(n9031), .IN2(n6978), .QN(n8477) );
  NAND4X0 U7326 ( .IN1(n5639), .IN2(n5638), .IN3(n8477), .IN4(n7377), .QN(
        \a6/N465 ) );
  NOR2X0 U7327 ( .IN1(n9204), .IN2(n8229), .QN(n5642) );
  NAND2X0 U7328 ( .IN1(n5640), .IN2(n9442), .QN(n8292) );
  NAND2X0 U7329 ( .IN1(n9047), .IN2(n6327), .QN(n8851) );
  NAND2X0 U7330 ( .IN1(n8292), .IN2(n8851), .QN(n5641) );
  NOR2X0 U7331 ( .IN1(n5642), .IN2(n5641), .QN(n5650) );
  NOR2X0 U7332 ( .IN1(n9442), .IN2(n7471), .QN(n8077) );
  OA21X1 U7333 ( .IN1(n7297), .IN2(n7964), .IN3(n9434), .Q(n5645) );
  NAND2X0 U7334 ( .IN1(n8534), .IN2(n9155), .QN(n8612) );
  INVX0 U7335 ( .INP(n8024), .ZN(n6489) );
  NAND2X0 U7336 ( .IN1(n8699), .IN2(n6489), .QN(n7587) );
  NAND4X0 U7337 ( .IN1(n8612), .IN2(n7729), .IN3(n7257), .IN4(n7587), .QN(
        n5644) );
  NAND2X0 U7338 ( .IN1(n5643), .IN2(n7589), .QN(n8928) );
  NAND2X0 U7339 ( .IN1(n8928), .IN2(n7288), .QN(n7147) );
  NOR4X0 U7340 ( .IN1(n8077), .IN2(n5645), .IN3(n5644), .IN4(n7147), .QN(n5649) );
  NAND3X0 U7341 ( .IN1(n8193), .IN2(n5646), .IN3(n8996), .QN(n5647) );
  NAND2X0 U7342 ( .IN1(n5647), .IN2(n9436), .QN(n5648) );
  NAND2X0 U7343 ( .IN1(n8180), .IN2(n7169), .QN(n8893) );
  NAND4X0 U7344 ( .IN1(n5650), .IN2(n5649), .IN3(n5648), .IN4(n8893), .QN(
        \a6/N466 ) );
  NOR2X0 U7345 ( .IN1(n6487), .IN2(n6720), .QN(n6834) );
  NOR2X0 U7346 ( .IN1(n6401), .IN2(n5651), .QN(n9091) );
  NOR2X0 U7347 ( .IN1(n8847), .IN2(n6373), .QN(n8430) );
  NOR2X0 U7348 ( .IN1(n8876), .IN2(n6150), .QN(n6993) );
  NAND2X0 U7349 ( .IN1(degrees_tmp2[2]), .IN2(n9060), .QN(n6966) );
  NOR2X0 U7350 ( .IN1(n8024), .IN2(n6966), .QN(n5652) );
  NOR4X0 U7351 ( .IN1(n9091), .IN2(n8430), .IN3(n6993), .IN4(n5652), .QN(n5660) );
  INVX0 U7352 ( .INP(n9195), .ZN(n8204) );
  NOR2X0 U7353 ( .IN1(n7035), .IN2(n8204), .QN(n7759) );
  NOR2X0 U7354 ( .IN1(n8349), .IN2(n8494), .QN(n5656) );
  NAND2X0 U7355 ( .IN1(n7654), .IN2(n6678), .QN(n7991) );
  NOR2X0 U7356 ( .IN1(n5653), .IN2(n6369), .QN(n7754) );
  NAND2X0 U7357 ( .IN1(n6614), .IN2(n7754), .QN(n7494) );
  NOR2X0 U7358 ( .IN1(n8489), .IN2(n6427), .QN(n7108) );
  NAND2X0 U7359 ( .IN1(n7108), .IN2(n8282), .QN(n5654) );
  NAND4X0 U7360 ( .IN1(n7991), .IN2(n7812), .IN3(n7494), .IN4(n5654), .QN(
        n5655) );
  NOR4X0 U7361 ( .IN1(n7984), .IN2(n7759), .IN3(n5656), .IN4(n5655), .QN(n5659) );
  NAND2X0 U7362 ( .IN1(n5657), .IN2(n7918), .QN(n5658) );
  NAND4X0 U7363 ( .IN1(n6834), .IN2(n5660), .IN3(n5659), .IN4(n5658), .QN(
        \a6/N467 ) );
  NAND2X0 U7364 ( .IN1(n8760), .IN2(n7035), .QN(n6070) );
  OA22X1 U7365 ( .IN1(n8495), .IN2(n6509), .IN3(n8268), .IN4(n6070), .Q(n5666)
         );
  NOR2X0 U7366 ( .IN1(n8489), .IN2(n6205), .QN(n5703) );
  NAND2X0 U7367 ( .IN1(n9208), .IN2(n9195), .QN(n6949) );
  OAI21X1 U7368 ( .IN1(n8595), .IN2(n6949), .IN3(n7789), .QN(n5664) );
  NAND2X0 U7369 ( .IN1(n8978), .IN2(n7121), .QN(n8028) );
  NAND2X0 U7370 ( .IN1(n8875), .IN2(n8572), .QN(n7845) );
  NAND4X0 U7371 ( .IN1(n7730), .IN2(n6305), .IN3(n8028), .IN4(n7845), .QN(
        n5663) );
  INVX0 U7372 ( .INP(n9156), .ZN(n8084) );
  NAND3X0 U7373 ( .IN1(degrees_tmp2[3]), .IN2(n7735), .IN3(n9023), .QN(n6662)
         );
  NAND2X0 U7374 ( .IN1(degrees_tmp2[5]), .IN2(n8848), .QN(n5926) );
  NAND3X0 U7375 ( .IN1(n8475), .IN2(n9445), .IN3(n9060), .QN(n5661) );
  NAND4X0 U7376 ( .IN1(n8084), .IN2(n6662), .IN3(n5926), .IN4(n5661), .QN(
        n5662) );
  NOR4X0 U7377 ( .IN1(n5703), .IN2(n5664), .IN3(n5663), .IN4(n5662), .QN(n5665) );
  NAND2X0 U7378 ( .IN1(n9437), .IN2(n6412), .QN(n6187) );
  INVX0 U7379 ( .INP(n6353), .ZN(n8039) );
  NAND2X0 U7380 ( .IN1(n6187), .IN2(n8039), .QN(n7221) );
  NAND2X0 U7381 ( .IN1(n8598), .IN2(n7221), .QN(n6555) );
  NAND4X0 U7382 ( .IN1(n5666), .IN2(n5665), .IN3(n8737), .IN4(n6555), .QN(
        \a6/N468 ) );
  NOR2X0 U7383 ( .IN1(n6257), .IN2(n8684), .QN(n5672) );
  INVX0 U7384 ( .INP(n5971), .ZN(n6961) );
  NOR2X0 U7385 ( .IN1(n9166), .IN2(n6961), .QN(n7146) );
  INVX0 U7386 ( .INP(n7146), .ZN(n8900) );
  NAND4X0 U7387 ( .IN1(n8778), .IN2(n5667), .IN3(n8399), .IN4(n8900), .QN(
        n5671) );
  INVX0 U7388 ( .INP(n9091), .ZN(n8913) );
  NOR2X0 U7389 ( .IN1(n8331), .IN2(n7914), .QN(n8698) );
  NAND2X0 U7390 ( .IN1(n9082), .IN2(n8698), .QN(n5669) );
  INVX0 U7391 ( .INP(n8276), .ZN(n7870) );
  NAND2X0 U7392 ( .IN1(n7870), .IN2(n7760), .QN(n5668) );
  NAND4X0 U7393 ( .IN1(n8524), .IN2(n8913), .IN3(n5669), .IN4(n5668), .QN(
        n5670) );
  OR4X1 U7394 ( .IN1(n6068), .IN2(n5672), .IN3(n5671), .IN4(n5670), .Q(
        \a6/N469 ) );
  NAND2X0 U7395 ( .IN1(n9182), .IN2(n7438), .QN(n6849) );
  OA22X1 U7396 ( .IN1(degrees_tmp2[3]), .IN2(n6949), .IN3(n6849), .IN4(n9442), 
        .Q(n5680) );
  NOR2X0 U7397 ( .IN1(degrees_tmp2[2]), .IN2(n8772), .QN(n9145) );
  AOI22X1 U7398 ( .IN1(n7169), .IN2(n9145), .IN3(n5673), .IN4(n7706), .QN(
        n5679) );
  NAND2X0 U7399 ( .IN1(n9434), .IN2(n8848), .QN(n8137) );
  INVX0 U7400 ( .INP(n8137), .ZN(n5677) );
  NAND2X0 U7401 ( .IN1(n9080), .IN2(n5949), .QN(n8412) );
  NAND3X0 U7402 ( .IN1(n7861), .IN2(n8962), .IN3(n8412), .QN(n5676) );
  NAND2X0 U7403 ( .IN1(n6946), .IN2(n6979), .QN(n7842) );
  NAND3X0 U7404 ( .IN1(n9434), .IN2(n7843), .IN3(n7842), .QN(n5674) );
  NAND4X0 U7405 ( .IN1(n8592), .IN2(n8167), .IN3(n6402), .IN4(n5674), .QN(
        n5675) );
  NOR4X0 U7406 ( .IN1(n8638), .IN2(n5677), .IN3(n5676), .IN4(n5675), .QN(n5678) );
  NAND4X0 U7407 ( .IN1(n5680), .IN2(n5679), .IN3(n5678), .IN4(n8817), .QN(
        \a6/N471 ) );
  NOR2X0 U7408 ( .IN1(n9213), .IN2(n5795), .QN(n6737) );
  NOR2X0 U7409 ( .IN1(n8432), .IN2(n7678), .QN(n8693) );
  NOR2X0 U7410 ( .IN1(n8693), .IN2(n8822), .QN(n7753) );
  NOR2X0 U7411 ( .IN1(n9440), .IN2(n8591), .QN(n6153) );
  NOR4X0 U7412 ( .IN1(n5788), .IN2(n5722), .IN3(n8674), .IN4(n6153), .QN(n5682) );
  NAND2X0 U7413 ( .IN1(n9210), .IN2(n9183), .QN(n8170) );
  OA22X1 U7414 ( .IN1(degrees_tmp2[5]), .IN2(n5894), .IN3(n8170), .IN4(n8588), 
        .Q(n5681) );
  NAND2X0 U7415 ( .IN1(n8728), .IN2(n7678), .QN(n7131) );
  INVX0 U7416 ( .INP(n8905), .ZN(n7973) );
  NAND2X0 U7417 ( .IN1(n7973), .IN2(n9438), .QN(n7563) );
  NAND4X0 U7418 ( .IN1(n5682), .IN2(n5681), .IN3(n7131), .IN4(n7563), .QN(
        n5683) );
  NOR4X0 U7419 ( .IN1(n7521), .IN2(n6737), .IN3(n7753), .IN4(n5683), .QN(n5684) );
  NAND4X0 U7420 ( .IN1(n5684), .IN2(n6534), .IN3(n6535), .IN4(n6249), .QN(
        \a6/N472 ) );
  NOR2X0 U7421 ( .IN1(n7405), .IN2(n6510), .QN(n5686) );
  NAND2X0 U7422 ( .IN1(n8968), .IN2(n6187), .QN(n5685) );
  NOR2X0 U7423 ( .IN1(n5686), .IN2(n5685), .QN(n5687) );
  NOR2X0 U7424 ( .IN1(n5687), .IN2(n8041), .QN(n5693) );
  NAND2X0 U7425 ( .IN1(n8467), .IN2(n7121), .QN(n7856) );
  NAND2X0 U7426 ( .IN1(n8697), .IN2(n6207), .QN(n7787) );
  NAND2X0 U7427 ( .IN1(n6360), .IN2(n9442), .QN(n5726) );
  NAND3X0 U7428 ( .IN1(n7856), .IN2(n7787), .IN3(n5726), .QN(n5692) );
  NAND2X0 U7429 ( .IN1(n9105), .IN2(n8978), .QN(n9079) );
  INVX0 U7430 ( .INP(n5688), .ZN(n7547) );
  OA22X1 U7431 ( .IN1(n9031), .IN2(n8705), .IN3(n9079), .IN4(n7547), .Q(n5690)
         );
  NAND3X0 U7432 ( .IN1(n9435), .IN2(n5949), .IN3(n8073), .QN(n5689) );
  NAND2X0 U7433 ( .IN1(n8728), .IN2(n7936), .QN(n9126) );
  NAND4X0 U7434 ( .IN1(n5690), .IN2(n6051), .IN3(n5689), .IN4(n9126), .QN(
        n5691) );
  NOR4X0 U7435 ( .IN1(n8359), .IN2(n5693), .IN3(n5692), .IN4(n5691), .QN(n5694) );
  NAND2X0 U7436 ( .IN1(n9190), .IN2(n6268), .QN(n8253) );
  NAND4X0 U7437 ( .IN1(n5694), .IN2(n8100), .IN3(n8524), .IN4(n8253), .QN(
        \a6/N473 ) );
  NAND2X0 U7438 ( .IN1(n6649), .IN2(n6613), .QN(n6441) );
  OA22X1 U7439 ( .IN1(n7437), .IN2(n8905), .IN3(n6441), .IN4(n6979), .Q(n5701)
         );
  NAND2X0 U7440 ( .IN1(n7517), .IN2(n5695), .QN(n7636) );
  NOR2X0 U7441 ( .IN1(n9442), .IN2(n7636), .QN(n8742) );
  OA22X1 U7442 ( .IN1(n8760), .IN2(n7824), .IN3(n8467), .IN4(n6727), .Q(n5698)
         );
  NAND2X0 U7443 ( .IN1(n5696), .IN2(n8073), .QN(n5774) );
  INVX0 U7444 ( .INP(n7412), .ZN(n7458) );
  NOR2X0 U7445 ( .IN1(n7945), .IN2(n6427), .QN(n7321) );
  OAI21X1 U7446 ( .IN1(n8888), .IN2(n7321), .IN3(n8886), .QN(n5697) );
  NAND4X0 U7447 ( .IN1(n5698), .IN2(n5774), .IN3(n7458), .IN4(n5697), .QN(
        n5699) );
  NOR4X0 U7448 ( .IN1(n6416), .IN2(n7077), .IN3(n8742), .IN4(n5699), .QN(n5700) );
  NAND2X0 U7449 ( .IN1(n8731), .IN2(n9071), .QN(n9006) );
  NAND4X0 U7450 ( .IN1(n5701), .IN2(n5700), .IN3(n7856), .IN4(n9006), .QN(
        \a6/N474 ) );
  INVX0 U7451 ( .INP(n6320), .ZN(n5822) );
  OA22X1 U7452 ( .IN1(n9189), .IN2(n5822), .IN3(n6614), .IN4(n8866), .Q(n5707)
         );
  NAND2X0 U7453 ( .IN1(n9190), .IN2(n9073), .QN(n9168) );
  NAND2X0 U7454 ( .IN1(n8796), .IN2(n7936), .QN(n6669) );
  OA22X1 U7455 ( .IN1(n8675), .IN2(n8470), .IN3(n8752), .IN4(n6669), .Q(n5702)
         );
  OA21X1 U7456 ( .IN1(n8249), .IN2(n9168), .IN3(n5702), .Q(n5706) );
  NAND2X0 U7457 ( .IN1(n8995), .IN2(n7735), .QN(n8487) );
  INVX0 U7458 ( .INP(n8487), .ZN(n6058) );
  INVX0 U7459 ( .INP(n5703), .ZN(n8803) );
  NAND4X0 U7460 ( .IN1(n8673), .IN2(n8043), .IN3(n8055), .IN4(n8803), .QN(
        n5704) );
  NOR4X0 U7461 ( .IN1(n7832), .IN2(n8319), .IN3(n6058), .IN4(n5704), .QN(n5705) );
  NAND4X0 U7462 ( .IN1(n5707), .IN2(n5706), .IN3(n5705), .IN4(n6131), .QN(
        \a6/N475 ) );
  INVX0 U7463 ( .INP(n8055), .ZN(n5715) );
  NAND2X0 U7464 ( .IN1(n9190), .IN2(n5708), .QN(n6118) );
  NAND2X0 U7465 ( .IN1(n6365), .IN2(n8947), .QN(n8802) );
  AND4X1 U7466 ( .IN1(n8689), .IN2(n8799), .IN3(n6118), .IN4(n8802), .Q(n5713)
         );
  NOR2X0 U7467 ( .IN1(n9084), .IN2(n8262), .QN(n6532) );
  AO22X1 U7468 ( .IN1(n5863), .IN2(n5709), .IN3(n6392), .IN4(n8588), .Q(n5710)
         );
  NOR4X0 U7469 ( .IN1(n7033), .IN2(n6532), .IN3(n6448), .IN4(n5710), .QN(n5712) );
  NAND2X0 U7470 ( .IN1(n9105), .IN2(n8675), .QN(n8845) );
  NAND2X0 U7471 ( .IN1(n8071), .IN2(n8845), .QN(n6556) );
  NAND2X0 U7472 ( .IN1(n9208), .IN2(n6556), .QN(n5711) );
  NAND4X0 U7473 ( .IN1(n5713), .IN2(n5712), .IN3(n9212), .IN4(n5711), .QN(
        n5714) );
  AO221X1 U7474 ( .IN1(n9183), .IN2(n7669), .IN3(n9183), .IN4(n5715), .IN5(
        n5714), .Q(\a6/N476 ) );
  INVX0 U7475 ( .INP(n8043), .ZN(n8994) );
  NOR2X0 U7476 ( .IN1(n8889), .IN2(n8494), .QN(n5721) );
  INVX0 U7477 ( .INP(n6414), .ZN(n8718) );
  INVX0 U7478 ( .INP(n5716), .ZN(n8726) );
  NOR2X0 U7479 ( .IN1(n8073), .IN2(n8726), .QN(n8178) );
  NOR2X0 U7480 ( .IN1(n8718), .IN2(n8178), .QN(n7351) );
  OA21X1 U7481 ( .IN1(n9073), .IN2(n9029), .IN3(n7943), .Q(n5847) );
  NOR2X0 U7482 ( .IN1(n8067), .IN2(n8995), .QN(n5718) );
  NAND2X0 U7483 ( .IN1(n5936), .IN2(n7589), .QN(n8967) );
  NAND2X0 U7484 ( .IN1(n8967), .IN2(n8885), .QN(n5717) );
  NOR2X0 U7485 ( .IN1(n5718), .IN2(n5717), .QN(n5719) );
  NAND4X0 U7486 ( .IN1(n7351), .IN2(n5847), .IN3(n5719), .IN4(n7060), .QN(
        n5720) );
  NOR4X0 U7487 ( .IN1(n8994), .IN2(n5722), .IN3(n5721), .IN4(n5720), .QN(n5724) );
  NAND2X0 U7488 ( .IN1(n9183), .IN2(n6274), .QN(n5723) );
  NAND4X0 U7489 ( .IN1(n5724), .IN2(n8292), .IN3(n6286), .IN4(n5723), .QN(
        \a6/N477 ) );
  INVX0 U7490 ( .INP(n6231), .ZN(n6266) );
  AND4X1 U7491 ( .IN1(n6150), .IN2(n8906), .IN3(n6266), .IN4(n8799), .Q(n5731)
         );
  NOR2X0 U7492 ( .IN1(n8386), .IN2(n6013), .QN(n8105) );
  NAND2X0 U7493 ( .IN1(n8890), .IN2(n6034), .QN(n8546) );
  NAND2X0 U7494 ( .IN1(n9075), .IN2(n8171), .QN(n5725) );
  NAND4X0 U7495 ( .IN1(n5727), .IN2(n5726), .IN3(n8546), .IN4(n5725), .QN(
        n5729) );
  INVX0 U7496 ( .INP(n8494), .ZN(n7668) );
  NOR2X0 U7497 ( .IN1(n7668), .IN2(n6337), .QN(n8142) );
  NOR2X0 U7498 ( .IN1(n8898), .IN2(n9033), .QN(n6256) );
  NOR2X0 U7499 ( .IN1(n6256), .IN2(n7035), .QN(n8415) );
  AO221X1 U7500 ( .IN1(n9434), .IN2(n9154), .IN3(n9434), .IN4(n8142), .IN5(
        n8415), .Q(n5728) );
  NOR4X0 U7501 ( .IN1(n6271), .IN2(n8105), .IN3(n5729), .IN4(n5728), .QN(n5730) );
  NAND4X0 U7502 ( .IN1(n5731), .IN2(n5730), .IN3(n5951), .IN4(n6135), .QN(
        \a6/N480 ) );
  NOR3X0 U7503 ( .IN1(n6124), .IN2(n5895), .IN3(n7645), .QN(n5732) );
  NOR2X0 U7504 ( .IN1(n5732), .IN2(n9061), .QN(n5738) );
  INVX0 U7505 ( .INP(n7751), .ZN(n8219) );
  NAND3X0 U7506 ( .IN1(n8511), .IN2(n5739), .IN3(n8724), .QN(n5733) );
  NAND4X0 U7507 ( .IN1(n5734), .IN2(n8219), .IN3(n6305), .IN4(n5733), .QN(
        n5737) );
  NOR2X0 U7508 ( .IN1(degrees_tmp2[2]), .IN2(n6823), .QN(n7342) );
  NAND2X0 U7509 ( .IN1(n7342), .IN2(n9433), .QN(n8607) );
  NAND2X0 U7510 ( .IN1(n6296), .IN2(n9061), .QN(n6008) );
  NAND2X0 U7511 ( .IN1(n9188), .IN2(n8947), .QN(n5735) );
  NAND4X0 U7512 ( .IN1(n6706), .IN2(n8607), .IN3(n6008), .IN4(n5735), .QN(
        n5736) );
  NOR4X0 U7513 ( .IN1(n9024), .IN2(n5738), .IN3(n5737), .IN4(n5736), .QN(n5741) );
  NOR2X0 U7514 ( .IN1(n9032), .IN2(n8880), .QN(n8257) );
  INVX0 U7515 ( .INP(n8257), .ZN(n5878) );
  NOR2X0 U7516 ( .IN1(n9047), .IN2(n5739), .QN(n8139) );
  INVX0 U7517 ( .INP(n8139), .ZN(n6326) );
  NAND3X0 U7518 ( .IN1(n7784), .IN2(n8978), .IN3(n6326), .QN(n5740) );
  NAND4X0 U7519 ( .IN1(n5741), .IN2(n7998), .IN3(n5878), .IN4(n5740), .QN(
        \a6/N481 ) );
  NAND3X0 U7520 ( .IN1(n6826), .IN2(n8171), .IN3(n8630), .QN(n7567) );
  OA22X1 U7521 ( .IN1(degrees_tmp2[0]), .IN2(n7567), .IN3(n6591), .IN4(n6198), 
        .Q(n5749) );
  OA22X1 U7522 ( .IN1(n6650), .IN2(n7881), .IN3(n8424), .IN4(n8705), .Q(n5748)
         );
  NOR2X0 U7523 ( .IN1(n8727), .IN2(n7463), .QN(n7586) );
  INVX0 U7524 ( .INP(n7842), .ZN(n5899) );
  INVX0 U7525 ( .INP(n6173), .ZN(n9196) );
  NOR2X0 U7526 ( .IN1(n5899), .IN2(n9196), .QN(n8993) );
  OA21X1 U7527 ( .IN1(n7586), .IN2(n8993), .IN3(degrees_tmp2[3]), .Q(n5744) );
  NAND2X0 U7528 ( .IN1(n5931), .IN2(n7784), .QN(n6909) );
  NAND4X0 U7529 ( .IN1(n5742), .IN2(n8737), .IN3(n6249), .IN4(n6909), .QN(
        n5743) );
  NOR4X0 U7530 ( .IN1(n7970), .IN2(n5745), .IN3(n5744), .IN4(n5743), .QN(n5747) );
  NAND2X0 U7531 ( .IN1(n7518), .IN2(n8692), .QN(n5746) );
  NAND4X0 U7532 ( .IN1(n5749), .IN2(n5748), .IN3(n5747), .IN4(n5746), .QN(
        \a6/N482 ) );
  INVX0 U7533 ( .INP(n8319), .ZN(n8809) );
  NAND2X0 U7534 ( .IN1(n8240), .IN2(n5750), .QN(n6130) );
  NAND2X0 U7535 ( .IN1(n8180), .IN2(n7956), .QN(n8152) );
  AND3X1 U7536 ( .IN1(n8809), .IN2(n6130), .IN3(n8152), .Q(n5756) );
  INVX0 U7537 ( .INP(n8244), .ZN(n9013) );
  OA21X1 U7538 ( .IN1(n7033), .IN2(n5751), .IN3(n9037), .Q(n5754) );
  NAND2X0 U7539 ( .IN1(n7861), .IN2(n6814), .QN(n6603) );
  NAND2X0 U7540 ( .IN1(n6942), .IN2(n9084), .QN(n6277) );
  NAND2X0 U7541 ( .IN1(n7198), .IN2(n8171), .QN(n5752) );
  NAND4X0 U7542 ( .IN1(n8708), .IN2(n8267), .IN3(n6277), .IN4(n5752), .QN(
        n5753) );
  NOR4X0 U7543 ( .IN1(n9013), .IN2(n5754), .IN3(n6603), .IN4(n5753), .QN(n5755) );
  NAND2X0 U7544 ( .IN1(n7870), .IN2(n9445), .QN(n7363) );
  INVX0 U7545 ( .INP(n8751), .ZN(n7670) );
  NAND2X0 U7546 ( .IN1(n9037), .IN2(n7670), .QN(n8615) );
  NAND4X0 U7547 ( .IN1(n5756), .IN2(n5755), .IN3(n7363), .IN4(n8615), .QN(
        \a6/N483 ) );
  INVX0 U7548 ( .INP(n8460), .ZN(n8303) );
  NOR2X0 U7549 ( .IN1(n5758), .IN2(n5757), .QN(n6292) );
  NOR2X0 U7550 ( .IN1(n8534), .IN2(n6292), .QN(n5759) );
  OA22X1 U7551 ( .IN1(n8730), .IN2(n8303), .IN3(n5759), .IN4(n7164), .Q(n5765)
         );
  NAND4X0 U7552 ( .IN1(n9437), .IN2(n6412), .IN3(n7945), .IN4(n8026), .QN(
        n7156) );
  OA221X1 U7553 ( .IN1(n8185), .IN2(n8262), .IN3(n8185), .IN4(n8007), .IN5(
        n7156), .Q(n5764) );
  NAND2X0 U7554 ( .IN1(n9436), .IN2(n7686), .QN(n9107) );
  OR2X1 U7555 ( .IN1(n8124), .IN2(n9107), .Q(n5760) );
  AND4X1 U7556 ( .IN1(n8183), .IN2(n7165), .IN3(n6305), .IN4(n5760), .Q(n5763)
         );
  NAND2X0 U7557 ( .IN1(n6936), .IN2(n5761), .QN(n6408) );
  AO221X1 U7558 ( .IN1(n9140), .IN2(n9434), .IN3(n9140), .IN4(n6408), .IN5(
        n7800), .Q(n5762) );
  NAND4X0 U7559 ( .IN1(n5765), .IN2(n5764), .IN3(n5763), .IN4(n5762), .QN(
        \a6/N484 ) );
  NAND2X0 U7560 ( .IN1(n5766), .IN2(n9071), .QN(n7051) );
  NOR2X0 U7561 ( .IN1(n8461), .IN2(n8213), .QN(n7999) );
  NAND2X0 U7562 ( .IN1(n7999), .IN2(n8034), .QN(n8444) );
  OA22X1 U7563 ( .IN1(n6921), .IN2(n7051), .IN3(n8444), .IN4(n6635), .Q(n5776)
         );
  NOR2X0 U7564 ( .IN1(n7437), .IN2(n7251), .QN(n9093) );
  AO22X1 U7565 ( .IN1(n9073), .IN2(n9093), .IN3(n5767), .IN4(n7597), .Q(n5773)
         );
  NAND4X0 U7566 ( .IN1(n8124), .IN2(n8445), .IN3(n8530), .IN4(n5768), .QN(
        n5771) );
  INVX0 U7567 ( .INP(n8893), .ZN(n6503) );
  NAND2X0 U7568 ( .IN1(n6503), .IN2(n9442), .QN(n9077) );
  NAND2X0 U7569 ( .IN1(n6620), .IN2(n8510), .QN(n5769) );
  NAND4X0 U7570 ( .IN1(n9077), .IN2(n9030), .IN3(n6312), .IN4(n5769), .QN(
        n5770) );
  AO22X1 U7571 ( .IN1(n9031), .IN2(n5771), .IN3(n9054), .IN4(n5770), .Q(n5772)
         );
  NOR2X0 U7572 ( .IN1(n5773), .IN2(n5772), .QN(n5775) );
  NAND4X0 U7573 ( .IN1(n5776), .IN2(n5775), .IN3(n7998), .IN4(n5774), .QN(
        \a6/N485 ) );
  OA22X1 U7574 ( .IN1(n8816), .IN2(n7394), .IN3(n9054), .IN4(n6908), .Q(n8216)
         );
  INVX0 U7575 ( .INP(n7445), .ZN(n8983) );
  INVX0 U7576 ( .INP(n6758), .ZN(n8040) );
  NOR2X0 U7577 ( .IN1(n9435), .IN2(n8040), .QN(n5777) );
  INVX0 U7578 ( .INP(n6859), .ZN(n6605) );
  NAND2X0 U7579 ( .IN1(n9023), .IN2(n8026), .QN(n6370) );
  NOR2X0 U7580 ( .IN1(n6605), .IN2(n6370), .QN(n6851) );
  NOR4X0 U7581 ( .IN1(n9074), .IN2(n8983), .IN3(n5777), .IN4(n6851), .QN(n5779) );
  NAND2X0 U7582 ( .IN1(n8468), .IN2(n8282), .QN(n6761) );
  OR2X1 U7583 ( .IN1(n8568), .IN2(n6624), .Q(n5778) );
  NAND4X0 U7584 ( .IN1(n8216), .IN2(n5779), .IN3(n6761), .IN4(n5778), .QN(
        \a6/N488 ) );
  INVX0 U7585 ( .INP(n6512), .ZN(n7472) );
  OA21X1 U7586 ( .IN1(n6342), .IN2(n7472), .IN3(n9213), .Q(n7422) );
  NAND3X0 U7587 ( .IN1(n9437), .IN2(n6620), .IN3(n5780), .QN(n8756) );
  NAND3X0 U7588 ( .IN1(n7422), .IN2(n8756), .IN3(n5781), .QN(\a6/N489 ) );
  AO21X1 U7589 ( .IN1(n9438), .IN2(n5786), .IN3(n6651), .Q(n5784) );
  NAND3X0 U7590 ( .IN1(n5784), .IN2(n5783), .IN3(n5782), .QN(\a6/N490 ) );
  NAND4X0 U7591 ( .IN1(n9212), .IN2(n8422), .IN3(n5785), .IN4(n5784), .QN(
        \a6/N491 ) );
  AND2X1 U7592 ( .IN1(n7699), .IN2(n5786), .Q(\a6/N492 ) );
  NAND2X0 U7593 ( .IN1(n9203), .IN2(n8467), .QN(n8491) );
  NOR2X0 U7594 ( .IN1(n8890), .IN2(n8491), .QN(n5787) );
  NOR2X0 U7595 ( .IN1(n7600), .IN2(n7466), .QN(n8462) );
  NOR4X0 U7596 ( .IN1(n6451), .IN2(n5787), .IN3(n7804), .IN4(n8462), .QN(n5794) );
  AND2X1 U7597 ( .IN1(n8026), .IN2(n8848), .Q(n8256) );
  NOR2X0 U7598 ( .IN1(n8728), .IN2(n7824), .QN(n8130) );
  NOR2X0 U7599 ( .IN1(n6371), .IN2(n7969), .QN(n7997) );
  NOR2X0 U7600 ( .IN1(n9166), .IN2(n9053), .QN(n7003) );
  NOR2X0 U7601 ( .IN1(n7997), .IN2(n7003), .QN(n6273) );
  NAND4X0 U7602 ( .IN1(degrees_tmp2[2]), .IN2(n8534), .IN3(n9054), .IN4(n9436), 
        .QN(n5790) );
  NAND2X0 U7603 ( .IN1(n5788), .IN2(n8004), .QN(n6206) );
  NOR2X0 U7604 ( .IN1(n8724), .IN2(n6059), .QN(n8518) );
  NAND2X0 U7605 ( .IN1(n8518), .IN2(n9440), .QN(n5789) );
  NAND4X0 U7606 ( .IN1(n6273), .IN2(n5790), .IN3(n6206), .IN4(n5789), .QN(
        n5791) );
  NOR4X0 U7607 ( .IN1(n9024), .IN2(n8256), .IN3(n8130), .IN4(n5791), .QN(n5793) );
  NAND4X0 U7608 ( .IN1(n5794), .IN2(n5793), .IN3(n5792), .IN4(n7308), .QN(
        \a5/N436 ) );
  OA22X1 U7609 ( .IN1(n7517), .IN2(n8706), .IN3(n5795), .IN4(n8495), .Q(n5802)
         );
  INVX0 U7610 ( .INP(n7856), .ZN(n8143) );
  NOR2X0 U7611 ( .IN1(n8710), .IN2(n7340), .QN(n5800) );
  NAND2X0 U7612 ( .IN1(n7699), .IN2(n8431), .QN(n7685) );
  NAND4X0 U7613 ( .IN1(n5822), .IN2(n7685), .IN3(n8574), .IN4(n7392), .QN(
        n5796) );
  NAND2X0 U7614 ( .IN1(n8825), .IN2(n5796), .QN(n5798) );
  NOR2X0 U7615 ( .IN1(n8534), .IN2(n6360), .QN(n7211) );
  OA22X1 U7616 ( .IN1(degrees_tmp2[3]), .IN2(n9006), .IN3(n7211), .IN4(n9166), 
        .Q(n5797) );
  NAND3X0 U7617 ( .IN1(n5798), .IN2(n7781), .IN3(n5797), .QN(n5799) );
  NOR4X0 U7618 ( .IN1(n8436), .IN2(n8143), .IN3(n5800), .IN4(n5799), .QN(n5801) );
  NAND2X0 U7619 ( .IN1(n6100), .IN2(n7233), .QN(n6078) );
  NAND4X0 U7620 ( .IN1(n5802), .IN2(n5801), .IN3(n6078), .IN4(n6131), .QN(
        \a5/N437 ) );
  NAND2X0 U7621 ( .IN1(degrees_tmp2[2]), .IN2(n9061), .QN(n8904) );
  AOI22X1 U7622 ( .IN1(n6194), .IN2(n7971), .IN3(n6292), .IN4(n8904), .QN(
        n5808) );
  NOR2X0 U7623 ( .IN1(n9435), .IN2(n9098), .QN(n6781) );
  AO22X1 U7624 ( .IN1(n6697), .IN2(n8630), .IN3(n6365), .IN4(n7656), .Q(n5805)
         );
  NOR2X0 U7625 ( .IN1(n7679), .IN2(n7760), .QN(n6453) );
  NAND2X0 U7626 ( .IN1(n8730), .IN2(n6453), .QN(n9177) );
  NOR2X0 U7627 ( .IN1(n9442), .IN2(n5803), .QN(n7916) );
  NAND2X0 U7628 ( .IN1(degrees_tmp2[5]), .IN2(n7916), .QN(n8719) );
  NOR2X0 U7629 ( .IN1(degrees_tmp2[5]), .IN2(n6832), .QN(n9035) );
  NAND2X0 U7630 ( .IN1(degrees_tmp2[3]), .IN2(n9035), .QN(n8230) );
  NAND3X0 U7631 ( .IN1(n9183), .IN2(n7669), .IN3(n9433), .QN(n8147) );
  NAND4X0 U7632 ( .IN1(n9177), .IN2(n8719), .IN3(n8230), .IN4(n8147), .QN(
        n5804) );
  NOR4X0 U7633 ( .IN1(n8566), .IN2(n6781), .IN3(n5805), .IN4(n5804), .QN(n5807) );
  NAND3X0 U7634 ( .IN1(degrees_tmp2[2]), .IN2(n8534), .IN3(n9054), .QN(n5806)
         );
  NAND4X0 U7635 ( .IN1(n5809), .IN2(n5808), .IN3(n5807), .IN4(n5806), .QN(
        \a5/N438 ) );
  NAND2X0 U7636 ( .IN1(n7236), .IN2(n9436), .QN(n8315) );
  NAND2X0 U7637 ( .IN1(n7347), .IN2(n8315), .QN(n6092) );
  OA22X1 U7638 ( .IN1(n8978), .IN2(n8706), .IN3(n9436), .IN4(n7954), .Q(n5813)
         );
  NOR2X0 U7639 ( .IN1(n9037), .IN2(n8452), .QN(n8378) );
  NAND4X0 U7640 ( .IN1(n9047), .IN2(degrees_tmp2[3]), .IN3(n9131), .IN4(n9032), 
        .QN(n7641) );
  NOR2X0 U7641 ( .IN1(n9436), .IN2(n7641), .QN(n5811) );
  NOR2X0 U7642 ( .IN1(n9213), .IN2(n8531), .QN(n7581) );
  NAND2X0 U7643 ( .IN1(n7581), .IN2(n7473), .QN(n7817) );
  AND3X1 U7644 ( .IN1(n8220), .IN2(n9037), .IN3(n9071), .Q(n7170) );
  NAND2X0 U7645 ( .IN1(n7170), .IN2(n9438), .QN(n6739) );
  NAND2X0 U7646 ( .IN1(n8408), .IN2(n9209), .QN(n6684) );
  NAND4X0 U7647 ( .IN1(n8219), .IN2(n7817), .IN3(n6739), .IN4(n6684), .QN(
        n5810) );
  NOR4X0 U7648 ( .IN1(n6360), .IN2(n8378), .IN3(n5811), .IN4(n5810), .QN(n5812) );
  NOR2X0 U7649 ( .IN1(n7858), .IN2(n6325), .QN(n6454) );
  OR2X1 U7650 ( .IN1(n8909), .IN2(n6454), .Q(n6355) );
  NAND4X0 U7651 ( .IN1(n5813), .IN2(n5812), .IN3(n7519), .IN4(n6355), .QN(
        n5814) );
  AO221X1 U7652 ( .IN1(n8533), .IN2(n6523), .IN3(n8533), .IN4(n6092), .IN5(
        n5814), .Q(\a5/N439 ) );
  NOR2X0 U7653 ( .IN1(n8978), .IN2(n6747), .QN(n8561) );
  NAND2X0 U7654 ( .IN1(n8188), .IN2(n8561), .QN(n7715) );
  NOR2X0 U7655 ( .IN1(degrees_tmp2[0]), .IN2(n7715), .QN(n5841) );
  NAND2X0 U7656 ( .IN1(n6016), .IN2(n6947), .QN(n8839) );
  NOR2X0 U7657 ( .IN1(n8710), .IN2(n9031), .QN(n7084) );
  INVX0 U7658 ( .INP(n7084), .ZN(n5815) );
  NAND4X0 U7659 ( .IN1(n8119), .IN2(degrees_tmp2[2]), .IN3(n8118), .IN4(n5815), 
        .QN(n6372) );
  NAND2X0 U7660 ( .IN1(n7841), .IN2(n6360), .QN(n5966) );
  NAND4X0 U7661 ( .IN1(n6112), .IN2(n8839), .IN3(n6372), .IN4(n5966), .QN(
        n5819) );
  INVX0 U7662 ( .INP(n6034), .ZN(n9072) );
  NAND3X0 U7663 ( .IN1(n9072), .IN2(n7721), .IN3(n9126), .QN(n5818) );
  AO22X1 U7664 ( .IN1(n5816), .IN2(n8598), .IN3(n5949), .IN4(n9001), .Q(n5817)
         );
  NOR4X0 U7665 ( .IN1(n5841), .IN2(n5819), .IN3(n5818), .IN4(n5817), .QN(n5820) );
  NAND4X0 U7666 ( .IN1(n5820), .IN2(n8624), .IN3(n6904), .IN4(n8007), .QN(
        \a5/N440 ) );
  INVX0 U7667 ( .INP(n8324), .ZN(n8338) );
  NAND3X0 U7668 ( .IN1(n5986), .IN2(n8730), .IN3(n5985), .QN(n8314) );
  AND2X1 U7669 ( .IN1(n8338), .IN2(n8314), .Q(n5979) );
  NAND4X0 U7670 ( .IN1(n9210), .IN2(n8699), .IN3(n7169), .IN4(n6946), .QN(
        n5821) );
  NAND2X0 U7671 ( .IN1(n8737), .IN2(n5821), .QN(n6010) );
  NAND2X0 U7672 ( .IN1(n5822), .IN2(n8574), .QN(n7701) );
  OR2X1 U7673 ( .IN1(n9195), .IN2(n6235), .Q(n8734) );
  AO22X1 U7674 ( .IN1(n9189), .IN2(n7701), .IN3(n8825), .IN4(n8734), .Q(n5829)
         );
  NAND2X0 U7675 ( .IN1(degrees_tmp2[3]), .IN2(n9023), .QN(n5824) );
  OA22X1 U7676 ( .IN1(n8890), .IN2(n8763), .IN3(n5824), .IN4(n5823), .Q(n5825)
         );
  NAND2X0 U7677 ( .IN1(n6826), .IN2(n6507), .QN(n6094) );
  NAND3X0 U7678 ( .IN1(n5825), .IN2(n6524), .IN3(n6094), .QN(n5828) );
  NAND2X0 U7679 ( .IN1(n7816), .IN2(n7035), .QN(n8225) );
  NOR2X0 U7680 ( .IN1(n9149), .IN2(n6059), .QN(n6688) );
  INVX0 U7681 ( .INP(n6688), .ZN(n5826) );
  NAND4X0 U7682 ( .IN1(n7738), .IN2(n8668), .IN3(n8225), .IN4(n5826), .QN(
        n5827) );
  NOR4X0 U7683 ( .IN1(n6010), .IN2(n5829), .IN3(n5828), .IN4(n5827), .QN(n5830) );
  NAND4X0 U7684 ( .IN1(n5831), .IN2(n5979), .IN3(n5830), .IN4(n8292), .QN(
        \a5/N441 ) );
  NAND3X0 U7685 ( .IN1(n8034), .IN2(n9209), .IN3(n5832), .QN(n5833) );
  AND2X1 U7686 ( .IN1(n8249), .IN2(n8118), .Q(n8862) );
  NAND2X0 U7687 ( .IN1(n9433), .IN2(n8862), .QN(n7349) );
  OR2X1 U7688 ( .IN1(n8822), .IN2(n7349), .Q(n9015) );
  NAND2X0 U7689 ( .IN1(n5833), .IN2(n9015), .QN(n6289) );
  NAND2X0 U7690 ( .IN1(n8567), .IN2(n7935), .QN(n8762) );
  INVX0 U7691 ( .INP(n8597), .ZN(n5834) );
  NAND2X0 U7692 ( .IN1(n5834), .IN2(n7956), .QN(n5835) );
  NAND4X0 U7693 ( .IN1(n8689), .IN2(n7377), .IN3(n8762), .IN4(n5835), .QN(
        n5840) );
  INVX0 U7694 ( .INP(n6720), .ZN(n8613) );
  NAND2X0 U7695 ( .IN1(n6613), .IN2(n9155), .QN(n6193) );
  OA22X1 U7696 ( .IN1(n7035), .IN2(n8613), .IN3(n7552), .IN4(n6193), .Q(n5838)
         );
  NAND2X0 U7697 ( .IN1(n8876), .IN2(n7093), .QN(n7975) );
  AO221X1 U7698 ( .IN1(n7118), .IN2(n9434), .IN3(n7118), .IN4(n7975), .IN5(
        n8424), .Q(n5836) );
  NAND4X0 U7699 ( .IN1(n5838), .IN2(n8720), .IN3(n5837), .IN4(n5836), .QN(
        n5839) );
  OR4X1 U7700 ( .IN1(n5841), .IN2(n6289), .IN3(n5840), .IN4(n5839), .Q(
        \a5/N442 ) );
  OA22X1 U7701 ( .IN1(n8977), .IN2(n7897), .IN3(n5842), .IN4(n7143), .Q(n5851)
         );
  NAND2X0 U7702 ( .IN1(n8249), .IN2(n5843), .QN(n7577) );
  NOR2X0 U7703 ( .IN1(n6624), .IN2(n8645), .QN(n8273) );
  NAND2X0 U7704 ( .IN1(n8796), .IN2(n8273), .QN(n7154) );
  INVX0 U7705 ( .INP(n7377), .ZN(n6481) );
  NOR2X0 U7706 ( .IN1(n8942), .IN2(n6481), .QN(n6099) );
  INVX0 U7707 ( .INP(n6142), .ZN(n5992) );
  NAND2X0 U7708 ( .IN1(n5992), .IN2(n6919), .QN(n7274) );
  OA22X1 U7709 ( .IN1(n8730), .IN2(n7274), .IN3(n9440), .IN4(n5844), .Q(n5846)
         );
  INVX0 U7710 ( .INP(n6373), .ZN(n6647) );
  NAND2X0 U7711 ( .IN1(n6647), .IN2(n7913), .QN(n5845) );
  AND4X1 U7712 ( .IN1(n5847), .IN2(n6099), .IN3(n5846), .IN4(n5845), .Q(n5848)
         );
  OA221X1 U7713 ( .IN1(n9436), .IN2(n7577), .IN3(n9436), .IN4(n7154), .IN5(
        n5848), .Q(n5850) );
  NAND2X0 U7714 ( .IN1(n9150), .IN2(n9019), .QN(n5849) );
  NAND4X0 U7715 ( .IN1(n5851), .IN2(n5850), .IN3(n8737), .IN4(n5849), .QN(
        \a5/N444 ) );
  NOR2X0 U7716 ( .IN1(n6541), .IN2(n8458), .QN(n8792) );
  NOR2X0 U7717 ( .IN1(n9437), .IN2(n6915), .QN(n6850) );
  INVX0 U7718 ( .INP(n7934), .ZN(n5852) );
  NAND2X0 U7719 ( .IN1(n8754), .IN2(n8674), .QN(n8059) );
  NAND2X0 U7720 ( .IN1(n5852), .IN2(n8059), .QN(n8930) );
  INVX0 U7721 ( .INP(n6220), .ZN(n6474) );
  NAND4X0 U7722 ( .IN1(n8778), .IN2(n7748), .IN3(n6474), .IN4(n6217), .QN(
        n5856) );
  NAND2X0 U7723 ( .IN1(n8485), .IN2(n8947), .QN(n5854) );
  NAND2X0 U7724 ( .IN1(n9435), .IN2(n6108), .QN(n6321) );
  NAND3X0 U7725 ( .IN1(n5854), .IN2(n5853), .IN3(n6321), .QN(n5855) );
  NOR4X0 U7726 ( .IN1(n6850), .IN2(n8930), .IN3(n5856), .IN4(n5855), .QN(n5857) );
  NAND2X0 U7727 ( .IN1(n6698), .IN2(n7784), .QN(n6001) );
  NAND4X0 U7728 ( .IN1(n8792), .IN2(n5857), .IN3(n6001), .IN4(n8591), .QN(
        \a5/N445 ) );
  NAND2X0 U7729 ( .IN1(n9433), .IN2(n9019), .QN(n7550) );
  NOR2X0 U7730 ( .IN1(n7550), .IN2(n8968), .QN(n5859) );
  NAND2X0 U7731 ( .IN1(n8685), .IN2(n8891), .QN(n5858) );
  NOR2X0 U7732 ( .IN1(n5859), .IN2(n5858), .QN(n5862) );
  NAND2X0 U7733 ( .IN1(n8731), .IN2(n8710), .QN(n8202) );
  NAND2X0 U7734 ( .IN1(n6417), .IN2(n8816), .QN(n8939) );
  INVX0 U7735 ( .INP(n8939), .ZN(n6246) );
  NAND2X0 U7736 ( .IN1(n9437), .IN2(n6246), .QN(n7635) );
  NAND4X0 U7737 ( .IN1(n7981), .IN2(n7824), .IN3(n8202), .IN4(n7635), .QN(
        n5860) );
  NOR4X0 U7738 ( .IN1(n8638), .IN2(n6416), .IN3(n6882), .IN4(n5860), .QN(n5861) );
  INVX0 U7739 ( .INP(n6359), .ZN(n7430) );
  NAND4X0 U7740 ( .IN1(n5862), .IN2(n5861), .IN3(n8338), .IN4(n7430), .QN(
        \a5/N446 ) );
  NAND2X0 U7741 ( .IN1(n8188), .IN2(n6697), .QN(n8375) );
  INVX0 U7742 ( .INP(n6781), .ZN(n7823) );
  NAND2X0 U7743 ( .IN1(n6758), .IN2(n5863), .QN(n7498) );
  NAND2X0 U7744 ( .IN1(n6067), .IN2(n8197), .QN(n5864) );
  NAND4X0 U7745 ( .IN1(n8375), .IN2(n7823), .IN3(n7498), .IN4(n5864), .QN(
        n5868) );
  OA21X1 U7746 ( .IN1(n7571), .IN2(n6371), .IN3(n7118), .Q(n5866) );
  NAND2X0 U7747 ( .IN1(n7518), .IN2(n8572), .QN(n6723) );
  NAND3X0 U7748 ( .IN1(n6699), .IN2(n5986), .IN3(n8034), .QN(n5865) );
  NAND4X0 U7749 ( .IN1(n5866), .IN2(n6888), .IN3(n6723), .IN4(n5865), .QN(
        n5867) );
  NOR4X0 U7750 ( .IN1(n5869), .IN2(n8832), .IN3(n5868), .IN4(n5867), .QN(n5871) );
  INVX0 U7751 ( .INP(n8408), .ZN(n8153) );
  NAND2X0 U7752 ( .IN1(n8153), .IN2(n8845), .QN(n6660) );
  NAND2X0 U7753 ( .IN1(n7880), .IN2(n6660), .QN(n5870) );
  NAND4X0 U7754 ( .IN1(n5871), .IN2(n8244), .IN3(n9140), .IN4(n5870), .QN(
        \a5/N448 ) );
  INVX0 U7755 ( .INP(n6311), .ZN(n6766) );
  AO22X1 U7756 ( .IN1(n6766), .IN2(n8978), .IN3(n5872), .IN4(n6326), .Q(n5875)
         );
  NAND2X0 U7757 ( .IN1(n8727), .IN2(n9074), .QN(n5972) );
  NAND4X0 U7758 ( .IN1(n6205), .IN2(n7392), .IN3(n8156), .IN4(n5972), .QN(
        n5874) );
  NAND2X0 U7759 ( .IN1(n6638), .IN2(n8728), .QN(n6437) );
  NAND4X0 U7760 ( .IN1(n8487), .IN2(n8607), .IN3(n8719), .IN4(n6437), .QN(
        n5873) );
  NOR4X0 U7761 ( .IN1(n5876), .IN2(n5875), .IN3(n5874), .IN4(n5873), .QN(n5879) );
  INVX0 U7762 ( .INP(n8968), .ZN(n8320) );
  NAND2X0 U7763 ( .IN1(n8320), .IN2(n9149), .QN(n8224) );
  NAND2X0 U7764 ( .IN1(n8646), .IN2(n7402), .QN(n5877) );
  NAND4X0 U7765 ( .IN1(n5879), .IN2(n5878), .IN3(n8224), .IN4(n5877), .QN(
        \a5/N449 ) );
  OA21X1 U7766 ( .IN1(n6016), .IN2(n8862), .IN3(n8572), .Q(n5883) );
  INVX0 U7767 ( .INP(n9079), .ZN(n7529) );
  NOR2X0 U7768 ( .IN1(n7033), .IN2(n7529), .QN(n7766) );
  NAND2X0 U7769 ( .IN1(n8995), .IN2(n5880), .QN(n5881) );
  NAND4X0 U7770 ( .IN1(n7766), .IN2(n6442), .IN3(n7223), .IN4(n5881), .QN(
        n5882) );
  NOR4X0 U7771 ( .IN1(n7520), .IN2(n8518), .IN3(n5883), .IN4(n5882), .QN(n5889) );
  NAND2X0 U7772 ( .IN1(n9434), .IN2(n7843), .QN(n5884) );
  NAND3X0 U7773 ( .IN1(n7349), .IN2(n5884), .IN3(n7183), .QN(n5885) );
  NAND2X0 U7774 ( .IN1(n5885), .IN2(n6614), .QN(n5888) );
  OAI21X1 U7775 ( .IN1(n7012), .IN2(n8825), .IN3(n7093), .QN(n5887) );
  NAND2X0 U7776 ( .IN1(n8163), .IN2(n8494), .QN(n5886) );
  NAND4X0 U7777 ( .IN1(n5889), .IN2(n5888), .IN3(n5887), .IN4(n5886), .QN(
        \a5/N450 ) );
  NOR2X0 U7778 ( .IN1(n9438), .IN2(n9100), .QN(n8472) );
  INVX0 U7779 ( .INP(n8082), .ZN(n5893) );
  NOR2X0 U7780 ( .IN1(degrees_tmp2[3]), .IN2(n6256), .QN(n5910) );
  NAND2X0 U7781 ( .IN1(n8268), .IN2(n8726), .QN(n7522) );
  OA21X1 U7782 ( .IN1(n5910), .IN2(n7522), .IN3(n8533), .Q(n5892) );
  INVX0 U7783 ( .INP(n7032), .ZN(n7057) );
  NAND2X0 U7784 ( .IN1(n7057), .IN2(n8169), .QN(n5890) );
  AO22X1 U7785 ( .IN1(n5995), .IN2(n5890), .IN3(n8247), .IN4(n7321), .Q(n5891)
         );
  NOR4X0 U7786 ( .IN1(n8472), .IN2(n5893), .IN3(n5892), .IN4(n5891), .QN(n5898) );
  NAND4X0 U7787 ( .IN1(degrees_tmp2[2]), .IN2(n9437), .IN3(n8000), .IN4(n8101), 
        .QN(n9028) );
  AO21X1 U7788 ( .IN1(n9028), .IN2(n5894), .IN3(n8588), .Q(n5896) );
  NAND3X0 U7789 ( .IN1(n5895), .IN2(n9440), .IN3(n8073), .QN(n7837) );
  NAND4X0 U7790 ( .IN1(n5898), .IN2(n5897), .IN3(n5896), .IN4(n7837), .QN(
        \a5/N451 ) );
  NOR2X0 U7791 ( .IN1(n6427), .IN2(n8083), .QN(n7681) );
  OA22X1 U7792 ( .IN1(n5899), .IN2(n8684), .IN3(n8431), .IN4(n6205), .Q(n5900)
         );
  NAND3X0 U7793 ( .IN1(n5900), .IN2(n8380), .IN3(n8737), .QN(n5905) );
  NOR2X0 U7794 ( .IN1(n6322), .IN2(n5901), .QN(n6382) );
  NOR2X0 U7795 ( .IN1(n8282), .IN2(n7465), .QN(n6856) );
  NOR4X0 U7796 ( .IN1(n6584), .IN2(n6451), .IN3(n6382), .IN4(n6856), .QN(n5903) );
  NAND2X0 U7797 ( .IN1(n8942), .IN2(n9445), .QN(n8807) );
  NAND2X0 U7798 ( .IN1(n8317), .IN2(n6187), .QN(n7036) );
  NAND2X0 U7799 ( .IN1(n7169), .IN2(n7036), .QN(n5902) );
  NAND4X0 U7800 ( .IN1(n5903), .IN2(n7225), .IN3(n8807), .IN4(n5902), .QN(
        n5904) );
  NOR4X0 U7801 ( .IN1(n7170), .IN2(n7681), .IN3(n5905), .IN4(n5904), .QN(n5909) );
  NOR2X0 U7802 ( .IN1(n7706), .IN2(n8763), .QN(n9039) );
  INVX0 U7803 ( .INP(n9039), .ZN(n6800) );
  NAND2X0 U7804 ( .IN1(n6766), .IN2(n8978), .QN(n5908) );
  NAND2X0 U7805 ( .IN1(n8118), .IN2(n5906), .QN(n5907) );
  NAND4X0 U7806 ( .IN1(n5909), .IN2(n6800), .IN3(n5908), .IN4(n5907), .QN(
        \a5/N452 ) );
  AND2X1 U7807 ( .IN1(n8533), .IN2(n5910), .Q(n5917) );
  INVX0 U7808 ( .INP(n6668), .ZN(n6773) );
  NAND2X0 U7809 ( .IN1(n9108), .IN2(n6773), .QN(n7161) );
  OA21X1 U7810 ( .IN1(n8181), .IN2(n7161), .IN3(n8816), .Q(n5916) );
  NOR2X0 U7811 ( .IN1(n9075), .IN2(n9025), .QN(n8686) );
  OA22X1 U7812 ( .IN1(n9125), .IN2(n8905), .IN3(n8686), .IN4(n8282), .Q(n5914)
         );
  NAND2X0 U7813 ( .IN1(n6182), .IN2(n7618), .QN(n8974) );
  NAND2X0 U7814 ( .IN1(n5912), .IN2(n5911), .QN(n6611) );
  NAND3X0 U7815 ( .IN1(n5913), .IN2(n9073), .IN3(n6611), .QN(n8818) );
  NAND2X0 U7816 ( .IN1(n9105), .IN2(n7179), .QN(n8265) );
  NAND4X0 U7817 ( .IN1(n5914), .IN2(n8974), .IN3(n8818), .IN4(n8265), .QN(
        n5915) );
  NOR3X0 U7818 ( .IN1(n5917), .IN2(n5916), .IN3(n5915), .QN(n5920) );
  NAND2X0 U7819 ( .IN1(n6412), .IN2(n7179), .QN(n7599) );
  INVX0 U7820 ( .INP(n8904), .ZN(n7515) );
  NAND3X0 U7821 ( .IN1(n9210), .IN2(n8188), .IN3(n7515), .QN(n5919) );
  NAND2X0 U7822 ( .IN1(n6353), .IN2(n8171), .QN(n5918) );
  NAND4X0 U7823 ( .IN1(n5920), .IN2(n7599), .IN3(n5919), .IN4(n5918), .QN(
        \a5/N453 ) );
  INVX0 U7824 ( .INP(n8412), .ZN(n6907) );
  NOR2X0 U7825 ( .IN1(n6163), .IN2(n6907), .QN(n6989) );
  INVX0 U7826 ( .INP(n7494), .ZN(n7222) );
  NOR2X0 U7827 ( .IN1(n8424), .IN2(n6908), .QN(n7775) );
  NOR2X0 U7828 ( .IN1(n9155), .IN2(n8527), .QN(n7366) );
  NOR4X0 U7829 ( .IN1(n7972), .IN2(n7222), .IN3(n7775), .IN4(n7366), .QN(n5924) );
  NOR2X0 U7830 ( .IN1(n8531), .IN2(n8104), .QN(n8628) );
  NOR2X0 U7831 ( .IN1(n9003), .IN2(n8494), .QN(n5922) );
  NAND2X0 U7832 ( .IN1(n9188), .IN2(n9001), .QN(n8860) );
  NAND2X0 U7833 ( .IN1(n7668), .IN2(n6647), .QN(n6655) );
  NAND4X0 U7834 ( .IN1(n7256), .IN2(n7060), .IN3(n8860), .IN4(n6655), .QN(
        n5921) );
  NOR4X0 U7835 ( .IN1(n7483), .IN2(n8628), .IN3(n5922), .IN4(n5921), .QN(n5923) );
  NOR2X0 U7836 ( .IN1(n9437), .IN2(n8996), .QN(n6667) );
  NAND2X0 U7837 ( .IN1(n9434), .IN2(n6667), .QN(n8060) );
  NAND4X0 U7838 ( .IN1(n6989), .IN2(n5924), .IN3(n5923), .IN4(n8060), .QN(
        \a5/N455 ) );
  NAND2X0 U7839 ( .IN1(n6365), .IN2(n6936), .QN(n5925) );
  NAND4X0 U7840 ( .IN1(n7010), .IN2(n5926), .IN3(n8208), .IN4(n5925), .QN(
        n5930) );
  INVX0 U7841 ( .INP(n7809), .ZN(n7070) );
  OA22X1 U7842 ( .IN1(n6182), .IN2(n8224), .IN3(n8675), .IN4(n7070), .Q(n5928)
         );
  INVX0 U7843 ( .INP(n8574), .ZN(n7235) );
  INVX0 U7844 ( .INP(n7895), .ZN(n9173) );
  AOI22X1 U7845 ( .IN1(n8947), .IN2(n7235), .IN3(n9173), .IN4(n5949), .QN(
        n5927) );
  NAND2X0 U7846 ( .IN1(n8512), .IN2(n9131), .QN(n5967) );
  NAND4X0 U7847 ( .IN1(n5928), .IN2(n5927), .IN3(n7378), .IN4(n5967), .QN(
        n5929) );
  NOR2X0 U7848 ( .IN1(n5930), .IN2(n5929), .QN(n5934) );
  INVX0 U7849 ( .INP(n7655), .ZN(n7094) );
  NAND3X0 U7850 ( .IN1(n5931), .IN2(degrees_tmp2[0]), .IN3(n7094), .QN(n5932)
         );
  NAND4X0 U7851 ( .IN1(n5934), .IN2(n5933), .IN3(n6800), .IN4(n5932), .QN(
        \a5/N456 ) );
  NOR2X0 U7852 ( .IN1(n9434), .IN2(n9031), .QN(n8861) );
  INVX0 U7853 ( .INP(n8861), .ZN(n8120) );
  INVX0 U7854 ( .INP(n6449), .ZN(n8545) );
  OA22X1 U7855 ( .IN1(n7679), .IN2(n8120), .IN3(n8568), .IN4(n8545), .Q(n5948)
         );
  INVX0 U7856 ( .INP(n8954), .ZN(n5935) );
  NAND2X0 U7857 ( .IN1(n8730), .IN2(n8728), .QN(n6024) );
  OA22X1 U7858 ( .IN1(n5935), .IN2(n6024), .IN3(n8446), .IN4(n7649), .Q(n5947)
         );
  NAND2X0 U7859 ( .IN1(n5937), .IN2(n5936), .QN(n6965) );
  INVX0 U7860 ( .INP(n6965), .ZN(n8429) );
  NAND2X0 U7861 ( .IN1(n6661), .IN2(n8429), .QN(n8618) );
  INVX0 U7862 ( .INP(n8618), .ZN(n5945) );
  NOR2X0 U7863 ( .IN1(n8947), .IN2(n7989), .QN(n8155) );
  NOR2X0 U7864 ( .IN1(n9001), .IN2(n7485), .QN(n5944) );
  NOR2X0 U7865 ( .IN1(n9155), .IN2(n6371), .QN(n7900) );
  INVX0 U7866 ( .INP(n7900), .ZN(n8299) );
  OA22X1 U7867 ( .IN1(n9434), .IN2(n8299), .IN3(n8730), .IN4(n7638), .Q(n5942)
         );
  NAND2X0 U7868 ( .IN1(n7049), .IN2(n6086), .QN(n7307) );
  NOR2X0 U7869 ( .IN1(n8630), .IN2(n7686), .QN(n5940) );
  NAND2X0 U7870 ( .IN1(n8889), .IN2(n5938), .QN(n5939) );
  NAND2X0 U7871 ( .IN1(n5940), .IN2(n5939), .QN(n5941) );
  NAND4X0 U7872 ( .IN1(n5942), .IN2(n7812), .IN3(n7307), .IN4(n5941), .QN(
        n5943) );
  NOR4X0 U7873 ( .IN1(n5945), .IN2(n8155), .IN3(n5944), .IN4(n5943), .QN(n5946) );
  NAND3X0 U7874 ( .IN1(n5948), .IN2(n5947), .IN3(n5946), .QN(\a5/N457 ) );
  NAND2X0 U7875 ( .IN1(n8001), .IN2(n9128), .QN(n7863) );
  NAND2X0 U7876 ( .IN1(n5949), .IN2(n7863), .QN(n8326) );
  INVX0 U7877 ( .INP(n8527), .ZN(n6543) );
  NAND2X0 U7878 ( .IN1(n8511), .IN2(n6543), .QN(n8998) );
  NAND2X0 U7879 ( .IN1(n6983), .IN2(n7842), .QN(n8355) );
  NAND3X0 U7880 ( .IN1(n8326), .IN2(n8998), .IN3(n8355), .QN(n5957) );
  INVX0 U7881 ( .INP(n7738), .ZN(n6862) );
  NAND2X0 U7882 ( .IN1(n9435), .IN2(n6862), .QN(n7951) );
  NAND2X0 U7883 ( .IN1(n7355), .IN2(n9445), .QN(n7364) );
  NAND2X0 U7884 ( .IN1(n8883), .IN2(n8988), .QN(n6433) );
  NAND2X0 U7885 ( .IN1(n8529), .IN2(n6755), .QN(n5950) );
  NAND4X0 U7886 ( .IN1(n7951), .IN2(n7364), .IN3(n6433), .IN4(n5950), .QN(
        n5956) );
  OA21X1 U7887 ( .IN1(n8886), .IN2(n7839), .IN3(n5951), .Q(n8175) );
  INVX0 U7888 ( .INP(n7521), .ZN(n7316) );
  OA22X1 U7889 ( .IN1(n7656), .IN2(n9027), .IN3(n8575), .IN4(n7316), .Q(n5953)
         );
  NAND3X0 U7890 ( .IN1(n6412), .IN2(n9441), .IN3(n8171), .QN(n5952) );
  NAND4X0 U7891 ( .IN1(n5954), .IN2(n8175), .IN3(n5953), .IN4(n5952), .QN(
        n5955) );
  OR4X1 U7892 ( .IN1(n8379), .IN2(n5957), .IN3(n5956), .IN4(n5955), .Q(
        \a5/N458 ) );
  NOR4X0 U7893 ( .IN1(n7296), .IN2(n9062), .IN3(n5958), .IN4(n8178), .QN(n5963) );
  AND3X1 U7894 ( .IN1(degrees_tmp2[2]), .IN2(n5965), .IN3(n8988), .Q(n7197) );
  NOR2X0 U7895 ( .IN1(n9132), .IN2(n7257), .QN(n5961) );
  NAND2X0 U7896 ( .IN1(n6697), .IN2(n9073), .QN(n8641) );
  NAND2X0 U7897 ( .IN1(n9125), .IN2(n8512), .QN(n8248) );
  NAND4X0 U7898 ( .IN1(n7018), .IN2(n8701), .IN3(n8641), .IN4(n8248), .QN(
        n5960) );
  INVX0 U7899 ( .INP(n7003), .ZN(n7891) );
  NAND2X0 U7900 ( .IN1(n7501), .IN2(n9155), .QN(n6157) );
  NAND4X0 U7901 ( .IN1(n7782), .IN2(n7767), .IN3(n7891), .IN4(n6157), .QN(
        n5959) );
  NOR4X0 U7902 ( .IN1(n7197), .IN2(n5961), .IN3(n5960), .IN4(n5959), .QN(n5962) );
  NAND4X0 U7903 ( .IN1(n5963), .IN2(n5962), .IN3(n9140), .IN4(n8230), .QN(
        \a5/N459 ) );
  NOR3X0 U7904 ( .IN1(n7806), .IN2(n7487), .IN3(n7486), .QN(n5964) );
  OA22X1 U7905 ( .IN1(n7784), .IN2(n5964), .IN3(n9442), .IN4(n6060), .Q(n5974)
         );
  NAND2X0 U7906 ( .IN1(n7501), .IN2(n5965), .QN(n7302) );
  NAND3X0 U7907 ( .IN1(n7485), .IN2(n5966), .IN3(n7302), .QN(n5970) );
  INVX0 U7908 ( .INP(n7850), .ZN(n9102) );
  NAND2X0 U7909 ( .IN1(n9102), .IN2(n5967), .QN(n5968) );
  AO22X1 U7910 ( .IN1(n6736), .IN2(n6805), .IN3(n9440), .IN4(n5968), .Q(n5969)
         );
  NOR4X0 U7911 ( .IN1(n8077), .IN2(n5971), .IN3(n5970), .IN4(n5969), .QN(n5973) );
  NAND2X0 U7912 ( .IN1(n7832), .IN2(n9440), .QN(n7990) );
  NAND4X0 U7913 ( .IN1(n5974), .IN2(n5973), .IN3(n5972), .IN4(n7990), .QN(
        \a5/N460 ) );
  INVX0 U7914 ( .INP(n5975), .ZN(n5976) );
  OA21X1 U7915 ( .IN1(n5976), .IN2(n8273), .IN3(n9125), .Q(n5983) );
  NAND2X0 U7916 ( .IN1(n7678), .IN2(n8026), .QN(n5977) );
  NAND4X0 U7917 ( .IN1(n7862), .IN2(n6433), .IN3(n8514), .IN4(n5977), .QN(
        n5982) );
  AO22X1 U7918 ( .IN1(n7870), .IN2(n8645), .IN3(n9154), .IN4(n8822), .Q(n5981)
         );
  OA22X1 U7919 ( .IN1(n9084), .IN2(n9098), .IN3(n8185), .IN4(n8550), .Q(n5978)
         );
  INVX0 U7920 ( .INP(n7415), .ZN(n8678) );
  NAND4X0 U7921 ( .IN1(n5979), .IN2(n5978), .IN3(n8678), .IN4(n8743), .QN(
        n5980) );
  OR4X1 U7922 ( .IN1(n5983), .IN2(n5982), .IN3(n5981), .IN4(n5980), .Q(
        \a5/N461 ) );
  NOR2X0 U7923 ( .IN1(n9066), .IN2(n5984), .QN(n8116) );
  OA21X1 U7924 ( .IN1(n8431), .IN2(n7431), .IN3(n8592), .Q(n5994) );
  INVX0 U7925 ( .INP(n7093), .ZN(n8903) );
  NOR2X0 U7926 ( .IN1(n8185), .IN2(n8903), .QN(n7250) );
  AO22X1 U7927 ( .IN1(n9031), .IN2(n7582), .IN3(n9080), .IN4(n7754), .Q(n5991)
         );
  OA22X1 U7928 ( .IN1(n7668), .IN2(n6373), .IN3(n8816), .IN4(n8859), .Q(n5989)
         );
  INVX0 U7929 ( .INP(n6891), .ZN(n9087) );
  NAND3X0 U7930 ( .IN1(n5986), .IN2(n7184), .IN3(n5985), .QN(n7330) );
  AND3X1 U7931 ( .IN1(n6312), .IN2(n9087), .IN3(n7330), .Q(n5987) );
  OA22X1 U7932 ( .IN1(n8533), .IN2(n8921), .IN3(n5987), .IN4(n8568), .Q(n5988)
         );
  INVX0 U7933 ( .INP(n6038), .ZN(n7805) );
  NAND2X0 U7934 ( .IN1(n8764), .IN2(n7805), .QN(n7968) );
  NAND4X0 U7935 ( .IN1(n5989), .IN2(n5988), .IN3(n7378), .IN4(n7968), .QN(
        n5990) );
  NOR4X0 U7936 ( .IN1(n5992), .IN2(n7250), .IN3(n5991), .IN4(n5990), .QN(n5993) );
  NAND4X0 U7937 ( .IN1(n8116), .IN2(n5994), .IN3(n5993), .IN4(n8928), .QN(
        \a5/N462 ) );
  INVX0 U7938 ( .INP(n7806), .ZN(n6039) );
  OA22X1 U7939 ( .IN1(n8760), .IN2(n8869), .IN3(n9054), .IN4(n6039), .Q(n6003)
         );
  NAND2X0 U7940 ( .IN1(n5995), .IN2(n8468), .QN(n5996) );
  NAND2X0 U7941 ( .IN1(n9102), .IN2(n5996), .QN(n5999) );
  NAND2X0 U7942 ( .IN1(n9074), .IN2(n7800), .QN(n8044) );
  OR2X1 U7943 ( .IN1(n7638), .IN2(n9054), .Q(n7188) );
  NAND4X0 U7944 ( .IN1(n7223), .IN2(n8044), .IN3(n7587), .IN4(n7188), .QN(
        n5998) );
  NAND2X0 U7945 ( .IN1(n9434), .IN2(n6781), .QN(n8056) );
  NAND2X0 U7946 ( .IN1(n9188), .IN2(n9166), .QN(n6375) );
  NAND4X0 U7947 ( .IN1(n8720), .IN2(n7771), .IN3(n8056), .IN4(n6375), .QN(
        n5997) );
  NOR4X0 U7948 ( .IN1(n6000), .IN2(n5999), .IN3(n5998), .IN4(n5997), .QN(n6002) );
  NAND4X0 U7949 ( .IN1(n6003), .IN2(n6002), .IN3(n8314), .IN4(n6001), .QN(
        \a5/N463 ) );
  NOR2X0 U7950 ( .IN1(n9053), .IN2(n8123), .QN(n6012) );
  OA21X1 U7951 ( .IN1(n6504), .IN2(n7500), .IN3(n7233), .Q(n6011) );
  NOR2X0 U7952 ( .IN1(n6649), .IN2(n8772), .QN(n8305) );
  NAND2X0 U7953 ( .IN1(n8598), .IN2(n8305), .QN(n6007) );
  INVX0 U7954 ( .INP(n7414), .ZN(n6951) );
  NAND3X0 U7955 ( .IN1(n7009), .IN2(n6951), .IN3(n7182), .QN(n6004) );
  NAND2X0 U7956 ( .IN1(n6004), .IN2(n9125), .QN(n6006) );
  NAND2X0 U7957 ( .IN1(n8567), .IN2(n8675), .QN(n7369) );
  NOR2X0 U7958 ( .IN1(n9434), .IN2(n8190), .QN(n8239) );
  INVX0 U7959 ( .INP(n8239), .ZN(n9207) );
  AO221X1 U7960 ( .IN1(n7369), .IN2(n8876), .IN3(n7369), .IN4(n9207), .IN5(
        n7760), .Q(n6005) );
  NAND4X0 U7961 ( .IN1(n6008), .IN2(n6007), .IN3(n6006), .IN4(n6005), .QN(
        n6009) );
  OR4X1 U7962 ( .IN1(n6012), .IN2(n6011), .IN3(n6010), .IN4(n6009), .Q(
        \a5/N464 ) );
  INVX0 U7963 ( .INP(n8461), .ZN(n9147) );
  OA22X1 U7964 ( .IN1(n8495), .IN2(n6013), .IN3(n9147), .IN4(n6728), .Q(n6014)
         );
  OA21X1 U7965 ( .IN1(n6979), .IN2(n8267), .IN3(n6014), .Q(n6023) );
  NOR2X0 U7966 ( .IN1(n9434), .IN2(n7340), .QN(n8660) );
  NAND2X0 U7967 ( .IN1(n7182), .IN2(n7635), .QN(n6594) );
  NOR4X0 U7968 ( .IN1(n9066), .IN2(n8888), .IN3(n8660), .IN4(n6594), .QN(n6022) );
  NOR2X0 U7969 ( .IN1(n8649), .IN2(n7404), .QN(n6037) );
  NOR2X0 U7970 ( .IN1(n9208), .IN2(n7018), .QN(n6393) );
  NAND2X0 U7971 ( .IN1(n6493), .IN2(n8728), .QN(n6015) );
  OA22X1 U7972 ( .IN1(n8754), .IN2(n8423), .IN3(n7613), .IN4(n6015), .Q(n6019)
         );
  NAND2X0 U7973 ( .IN1(n8730), .IN2(n6016), .QN(n6018) );
  NAND2X0 U7974 ( .IN1(n8180), .IN2(n6017), .QN(n7865) );
  NAND4X0 U7975 ( .IN1(n6019), .IN2(n6811), .IN3(n6018), .IN4(n7865), .QN(
        n6020) );
  NOR4X0 U7976 ( .IN1(n6504), .IN2(n6037), .IN3(n6393), .IN4(n6020), .QN(n6021) );
  NAND2X0 U7977 ( .IN1(n8289), .IN2(n9032), .QN(n6520) );
  NAND4X0 U7978 ( .IN1(n6023), .IN2(n6022), .IN3(n6021), .IN4(n6520), .QN(
        \a5/N465 ) );
  OA22X1 U7979 ( .IN1(n8188), .IN2(n8545), .IN3(n6024), .IN4(n6747), .Q(n6033)
         );
  NOR2X0 U7980 ( .IN1(n8124), .IN2(n9037), .QN(n6026) );
  NAND2X0 U7981 ( .IN1(n9025), .IN2(n8595), .QN(n7509) );
  NAND2X0 U7982 ( .IN1(n7509), .IN2(n6835), .QN(n6025) );
  NOR2X0 U7983 ( .IN1(n6026), .IN2(n6025), .QN(n6027) );
  NOR2X0 U7984 ( .IN1(n7784), .IN2(n6027), .QN(n6030) );
  OA221X1 U7985 ( .IN1(n7221), .IN2(n7414), .IN3(n7221), .IN4(n9440), .IN5(
        n8760), .Q(n6029) );
  OA21X1 U7986 ( .IN1(n6859), .IN2(n6983), .IN3(n8727), .Q(n6028) );
  NOR4X0 U7987 ( .IN1(n6031), .IN2(n6030), .IN3(n6029), .IN4(n6028), .QN(n6032) );
  NAND2X0 U7988 ( .IN1(n8710), .IN2(n7428), .QN(n6730) );
  NAND4X0 U7989 ( .IN1(n6033), .IN2(n6032), .IN3(n8426), .IN4(n6730), .QN(
        \a5/N466 ) );
  INVX0 U7990 ( .INP(n7195), .ZN(n8401) );
  OA22X1 U7991 ( .IN1(n9208), .IN2(n6727), .IN3(n8401), .IN4(n8782), .Q(n6046)
         );
  NOR2X0 U7992 ( .IN1(n6771), .IN2(n6034), .QN(n6036) );
  AND3X1 U7993 ( .IN1(n8268), .IN2(n6773), .IN3(n9027), .Q(n6035) );
  OA22X1 U7994 ( .IN1(n8890), .IN2(n6036), .IN3(n6035), .IN4(n7736), .Q(n6045)
         );
  INVX0 U7995 ( .INP(n6037), .ZN(n7205) );
  AND4X1 U7996 ( .IN1(n9129), .IN2(n9102), .IN3(n7636), .IN4(n7205), .Q(n6044)
         );
  NOR2X0 U7997 ( .IN1(n6038), .IN2(n9031), .QN(n6042) );
  NAND2X0 U7998 ( .IN1(n6119), .IN2(n7597), .QN(n8526) );
  OA22X1 U7999 ( .IN1(n8728), .IN2(n6039), .IN3(n8350), .IN4(n8526), .Q(n6040)
         );
  NAND2X0 U8000 ( .IN1(n6040), .IN2(n9140), .QN(n6041) );
  NOR2X0 U8001 ( .IN1(n6042), .IN2(n6041), .QN(n6043) );
  NAND4X0 U8002 ( .IN1(n6046), .IN2(n6045), .IN3(n6044), .IN4(n6043), .QN(
        \a5/N467 ) );
  INVX0 U8003 ( .INP(n7362), .ZN(n7008) );
  NOR2X0 U8004 ( .IN1(n9208), .IN2(n6205), .QN(n6048) );
  NOR2X0 U8005 ( .IN1(n9438), .IN2(n9027), .QN(n7506) );
  NOR2X0 U8006 ( .IN1(n8321), .IN2(n6568), .QN(n6047) );
  NOR4X0 U8007 ( .IN1(n7008), .IN2(n6048), .IN3(n7506), .IN4(n6047), .QN(n6057) );
  NOR2X0 U8008 ( .IN1(n6049), .IN2(n7293), .QN(n8683) );
  NOR2X0 U8009 ( .IN1(n8138), .IN2(n6408), .QN(n6054) );
  OA22X1 U8010 ( .IN1(n8760), .IN2(n8882), .IN3(n8764), .IN4(n9192), .Q(n6052)
         );
  NAND2X0 U8011 ( .IN1(n8534), .IN2(n9054), .QN(n6050) );
  NAND4X0 U8012 ( .IN1(n6052), .IN2(n9110), .IN3(n6051), .IN4(n6050), .QN(
        n6053) );
  NOR4X0 U8013 ( .IN1(n6055), .IN2(n8683), .IN3(n6054), .IN4(n6053), .QN(n6056) );
  NAND2X0 U8014 ( .IN1(n8533), .IN2(n8181), .QN(n7259) );
  NAND4X0 U8015 ( .IN1(n6834), .IN2(n6057), .IN3(n6056), .IN4(n7259), .QN(
        \a5/N468 ) );
  NOR2X0 U8016 ( .IN1(n9437), .IN2(n7070), .QN(n8629) );
  NOR4X0 U8017 ( .IN1(n6163), .IN2(n9091), .IN3(n6058), .IN4(n8629), .QN(n6066) );
  INVX0 U8018 ( .INP(n7213), .ZN(n7462) );
  NOR2X0 U8019 ( .IN1(n6059), .IN2(n7462), .QN(n6064) );
  NOR2X0 U8020 ( .IN1(n9438), .IN2(n6060), .QN(n8066) );
  NAND2X0 U8021 ( .IN1(n6275), .IN2(n9445), .QN(n8281) );
  NAND2X0 U8022 ( .IN1(n7271), .IN2(n7142), .QN(n8410) );
  INVX0 U8023 ( .INP(n8685), .ZN(n6110) );
  NAND2X0 U8024 ( .IN1(n6110), .IN2(n8041), .QN(n6061) );
  NAND4X0 U8025 ( .IN1(n8281), .IN2(n6373), .IN3(n8410), .IN4(n6061), .QN(
        n6063) );
  INVX0 U8026 ( .INP(n7550), .ZN(n8696) );
  NAND2X0 U8027 ( .IN1(n9047), .IN2(n8696), .QN(n6197) );
  NAND4X0 U8028 ( .IN1(n8891), .IN2(n6728), .IN3(n6669), .IN4(n6197), .QN(
        n6062) );
  NOR4X0 U8029 ( .IN1(n6064), .IN2(n8066), .IN3(n6063), .IN4(n6062), .QN(n6065) );
  NAND4X0 U8030 ( .IN1(n6066), .IN2(n6065), .IN3(n6072), .IN4(n8208), .QN(
        \a5/N469 ) );
  OA22X1 U8031 ( .IN1(n8947), .IN2(n9027), .IN3(n7164), .IN4(n7954), .Q(n6077)
         );
  NAND2X0 U8032 ( .IN1(n6067), .IN2(n6920), .QN(n8403) );
  OA22X1 U8033 ( .IN1(degrees_tmp2[2]), .IN2(n8403), .IN3(n6391), .IN4(n9002), 
        .Q(n6074) );
  INVX0 U8034 ( .INP(n6068), .ZN(n6071) );
  OA22X1 U8035 ( .IN1(degrees_tmp2[0]), .IN2(n6071), .IN3(n6070), .IN4(n6069), 
        .Q(n6073) );
  AND4X1 U8036 ( .IN1(n6074), .IN2(n6073), .IN3(n6072), .IN4(n6249), .Q(n6075)
         );
  OA221X1 U8037 ( .IN1(n8730), .IN2(n6811), .IN3(n8730), .IN4(n8587), .IN5(
        n6075), .Q(n6076) );
  NAND2X0 U8038 ( .IN1(n9435), .IN2(n9005), .QN(n8367) );
  NAND4X0 U8039 ( .IN1(n6077), .IN2(n6076), .IN3(n8778), .IN4(n8367), .QN(
        \a5/N470 ) );
  INVX0 U8040 ( .INP(n8518), .ZN(n7872) );
  INVX0 U8041 ( .INP(n7355), .ZN(n6982) );
  NAND2X0 U8042 ( .IN1(n8485), .IN2(n8198), .QN(n6996) );
  NAND4X0 U8043 ( .IN1(n7872), .IN2(n6982), .IN3(n6078), .IN4(n6996), .QN(
        n6080) );
  INVX0 U8044 ( .INP(n8519), .ZN(n6497) );
  NAND4X0 U8045 ( .IN1(n6497), .IN2(n8869), .IN3(n6567), .IN4(n7118), .QN(
        n6079) );
  NOR4X0 U8046 ( .IN1(n6448), .IN2(n7984), .IN3(n6080), .IN4(n6079), .QN(n6084) );
  NAND2X0 U8047 ( .IN1(n8384), .IN2(n8587), .QN(n6081) );
  NAND2X0 U8048 ( .IN1(degrees_tmp2[3]), .IN2(n6081), .QN(n6083) );
  NAND2X0 U8049 ( .IN1(n8710), .IN2(n8241), .QN(n6082) );
  NAND4X0 U8050 ( .IN1(n6084), .IN2(n7259), .IN3(n6083), .IN4(n6082), .QN(
        \a5/N471 ) );
  NOR2X0 U8051 ( .IN1(n8001), .IN2(n8726), .QN(n8369) );
  NAND2X0 U8052 ( .IN1(n6086), .IN2(n6085), .QN(n6087) );
  NAND4X0 U8053 ( .IN1(n8964), .IN2(n8885), .IN3(n6088), .IN4(n6087), .QN(
        n6097) );
  NOR2X0 U8054 ( .IN1(n6728), .IN2(n8461), .QN(n6091) );
  INVX0 U8055 ( .INP(n8106), .ZN(n6089) );
  NOR3X0 U8056 ( .IN1(n6091), .IN2(n6090), .IN3(n6089), .QN(n6095) );
  NAND2X0 U8057 ( .IN1(n6461), .IN2(n9061), .QN(n8941) );
  NAND2X0 U8058 ( .IN1(n8796), .IN2(n6092), .QN(n6093) );
  NAND4X0 U8059 ( .IN1(n6095), .IN2(n6094), .IN3(n8941), .IN4(n6093), .QN(
        n6096) );
  OR4X1 U8060 ( .IN1(n6231), .IN2(n8369), .IN3(n6097), .IN4(n6096), .Q(
        \a5/N472 ) );
  OA22X1 U8061 ( .IN1(n7402), .IN2(n8763), .IN3(n6605), .IN4(n8227), .Q(n6107)
         );
  NAND2X0 U8062 ( .IN1(n6466), .IN2(n8522), .QN(n6098) );
  OA21X1 U8063 ( .IN1(n6213), .IN2(n6098), .IN3(n9073), .Q(n6105) );
  NOR2X0 U8064 ( .IN1(n6099), .IN2(n9445), .QN(n8048) );
  AO22X1 U8065 ( .IN1(n8727), .IN2(n6100), .IN3(n8460), .IN4(n9060), .Q(n6104)
         );
  INVX0 U8066 ( .INP(n8294), .ZN(n7300) );
  NAND2X0 U8067 ( .IN1(n7300), .IN2(n9166), .QN(n7770) );
  NAND2X0 U8068 ( .IN1(n6647), .IN2(n8229), .QN(n6102) );
  NAND2X0 U8069 ( .IN1(n8728), .IN2(n8561), .QN(n6101) );
  NAND4X0 U8070 ( .IN1(n8607), .IN2(n7770), .IN3(n6102), .IN4(n6101), .QN(
        n6103) );
  NOR4X0 U8071 ( .IN1(n6105), .IN2(n8048), .IN3(n6104), .IN4(n6103), .QN(n6106) );
  INVX0 U8072 ( .INP(n7997), .ZN(n7453) );
  NAND4X0 U8073 ( .IN1(n6107), .IN2(n6106), .IN3(n6112), .IN4(n7453), .QN(
        \a5/N473 ) );
  INVX0 U8074 ( .INP(n7816), .ZN(n7822) );
  OA22X1 U8075 ( .IN1(n8876), .IN2(n7822), .IN3(n8550), .IN4(n8904), .Q(n6117)
         );
  NOR2X0 U8076 ( .IN1(n7164), .IN2(n8294), .QN(n6744) );
  INVX0 U8077 ( .INP(n6108), .ZN(n6167) );
  NOR2X0 U8078 ( .IN1(n8531), .IN2(n6120), .QN(n7312) );
  OAI21X1 U8079 ( .IN1(n7354), .IN2(n7312), .IN3(n9189), .QN(n6109) );
  NAND4X0 U8080 ( .IN1(n9200), .IN2(n6167), .IN3(n8202), .IN4(n6109), .QN(
        n6114) );
  NAND2X0 U8081 ( .IN1(n6110), .IN2(n9155), .QN(n6111) );
  NAND4X0 U8082 ( .IN1(n6112), .IN2(n6312), .IN3(n7205), .IN4(n6111), .QN(
        n6113) );
  NOR4X0 U8083 ( .IN1(n6744), .IN2(n6147), .IN3(n6114), .IN4(n6113), .QN(n6116) );
  NAND2X0 U8084 ( .IN1(n9212), .IN2(n8564), .QN(n9036) );
  NAND2X0 U8085 ( .IN1(n9433), .IN2(n9036), .QN(n6115) );
  NAND4X0 U8086 ( .IN1(n6117), .IN2(n6116), .IN3(n8060), .IN4(n6115), .QN(
        \a5/N474 ) );
  OA22X1 U8087 ( .IN1(n8752), .IN2(n8880), .IN3(n8249), .IN4(n6118), .Q(n6129)
         );
  AOI22X1 U8088 ( .IN1(n6119), .IN2(n6983), .IN3(n6392), .IN4(n6863), .QN(
        n6128) );
  NOR2X0 U8089 ( .IN1(n6833), .IN2(n6120), .QN(n6745) );
  NOR2X0 U8090 ( .IN1(n9060), .IN2(n8564), .QN(n6913) );
  NOR2X0 U8091 ( .IN1(n7463), .IN2(n6370), .QN(n6122) );
  INVX0 U8092 ( .INP(n6153), .ZN(n8448) );
  NAND4X0 U8093 ( .IN1(n8800), .IN2(n6985), .IN3(n8448), .IN4(n8546), .QN(
        n6121) );
  NOR4X0 U8094 ( .IN1(n6745), .IN2(n6913), .IN3(n6122), .IN4(n6121), .QN(n6127) );
  NOR3X0 U8095 ( .IN1(n6651), .IN2(n9435), .IN3(n9189), .QN(n6123) );
  OR4X1 U8096 ( .IN1(n6766), .IN2(n6124), .IN3(n7421), .IN4(n6123), .Q(n6125)
         );
  NAND2X0 U8097 ( .IN1(n7169), .IN2(n6125), .QN(n6126) );
  NAND4X0 U8098 ( .IN1(n6129), .IN2(n6128), .IN3(n6127), .IN4(n6126), .QN(
        \a5/N475 ) );
  INVX0 U8099 ( .INP(n7558), .ZN(n6751) );
  NAND4X0 U8100 ( .IN1(n7587), .IN2(n6600), .IN3(n6131), .IN4(n6130), .QN(
        n6141) );
  NOR2X0 U8101 ( .IN1(n9053), .IN2(n9019), .QN(n8986) );
  NAND2X0 U8102 ( .IN1(n9434), .IN2(n8986), .QN(n6924) );
  INVX0 U8103 ( .INP(n8855), .ZN(n6133) );
  INVX0 U8104 ( .INP(n6286), .ZN(n7801) );
  NAND2X0 U8105 ( .IN1(n7801), .IN2(n7736), .QN(n6132) );
  NAND4X0 U8106 ( .IN1(n6134), .IN2(n6924), .IN3(n6133), .IN4(n6132), .QN(
        n6140) );
  OA21X1 U8107 ( .IN1(n8489), .IN2(n6135), .IN3(n8338), .Q(n6138) );
  INVX0 U8108 ( .INP(n7640), .ZN(n6945) );
  NAND2X0 U8109 ( .IN1(n8468), .IN2(n6136), .QN(n6137) );
  NAND4X0 U8110 ( .IN1(n6138), .IN2(n7940), .IN3(n6945), .IN4(n6137), .QN(
        n6139) );
  OR4X1 U8111 ( .IN1(n6751), .IN2(n6141), .IN3(n6140), .IN4(n6139), .Q(
        \a5/N476 ) );
  NOR2X0 U8112 ( .IN1(n6142), .IN2(n8730), .QN(n6145) );
  AO21X1 U8113 ( .IN1(n7169), .IN2(n8119), .IN3(n7589), .Q(n8222) );
  NAND2X0 U8114 ( .IN1(n6143), .IN2(n8222), .QN(n6677) );
  NAND2X0 U8115 ( .IN1(n6677), .IN2(n8522), .QN(n6144) );
  NOR2X0 U8116 ( .IN1(n6145), .IN2(n6144), .QN(n6152) );
  NOR4X0 U8117 ( .IN1(n8888), .IN2(n8144), .IN3(n6147), .IN4(n6146), .QN(n6151) );
  NAND2X0 U8118 ( .IN1(n8461), .IN2(n6148), .QN(n8535) );
  NOR2X0 U8119 ( .IN1(n7529), .IN2(n7727), .QN(n8081) );
  AO221X1 U8120 ( .IN1(n8535), .IN2(n8081), .IN3(n8535), .IN4(n9435), .IN5(
        n9436), .Q(n6149) );
  NAND4X0 U8121 ( .IN1(n6152), .IN2(n6151), .IN3(n6150), .IN4(n6149), .QN(
        \a5/N477 ) );
  NAND2X0 U8122 ( .IN1(n9437), .IN2(n6153), .QN(n8339) );
  OA22X1 U8123 ( .IN1(degrees_tmp2[2]), .IN2(n8339), .IN3(n7668), .IN4(n7392), 
        .Q(n6166) );
  AO22X1 U8124 ( .IN1(n8180), .IN2(n7389), .IN3(n6155), .IN4(n6154), .Q(n6161)
         );
  INVX0 U8125 ( .INP(n6156), .ZN(n7828) );
  AND2X1 U8126 ( .IN1(n7082), .IN2(n7828), .Q(n7853) );
  INVX0 U8127 ( .INP(n8206), .ZN(n8593) );
  OA22X1 U8128 ( .IN1(n9438), .IN2(n6157), .IN3(n9122), .IN4(n8593), .Q(n6159)
         );
  INVX0 U8129 ( .INP(n8986), .ZN(n6158) );
  NAND4X0 U8130 ( .IN1(n7853), .IN2(n6159), .IN3(n8070), .IN4(n6158), .QN(
        n6160) );
  NOR4X0 U8131 ( .IN1(n6163), .IN2(n6162), .IN3(n6161), .IN4(n6160), .QN(n6165) );
  NAND3X0 U8132 ( .IN1(n6461), .IN2(n9440), .IN3(n8649), .QN(n6164) );
  NAND4X0 U8133 ( .IN1(n6166), .IN2(n6165), .IN3(n6535), .IN4(n6164), .QN(
        \a5/N478 ) );
  INVX0 U8134 ( .INP(n6541), .ZN(n8677) );
  NAND2X0 U8135 ( .IN1(n7754), .IN2(n9166), .QN(n8576) );
  NAND4X0 U8136 ( .IN1(n8677), .IN2(n6167), .IN3(n6591), .IN4(n8576), .QN(
        n6172) );
  NAND3X0 U8137 ( .IN1(degrees_tmp2[0]), .IN2(n8198), .IN3(n8197), .QN(n7884)
         );
  NAND4X0 U8138 ( .IN1(n8809), .IN2(n7009), .IN3(n8737), .IN4(n7884), .QN(
        n6171) );
  INVX0 U8139 ( .INP(n8921), .ZN(n7413) );
  NAND2X0 U8140 ( .IN1(n7413), .IN2(n8026), .QN(n6440) );
  INVX0 U8141 ( .INP(n7049), .ZN(n8700) );
  NAND2X0 U8142 ( .IN1(n8700), .IN2(n8004), .QN(n7879) );
  NAND2X0 U8143 ( .IN1(n6261), .IN2(n7879), .QN(n6679) );
  NAND2X0 U8144 ( .IN1(n8566), .IN2(n8675), .QN(n6168) );
  NAND4X0 U8145 ( .IN1(n6169), .IN2(n6440), .IN3(n6679), .IN4(n6168), .QN(
        n6170) );
  OR4X1 U8146 ( .IN1(n8559), .IN2(n6172), .IN3(n6171), .IN4(n6170), .Q(
        \a5/N479 ) );
  OA22X1 U8147 ( .IN1(n8816), .IN2(n9165), .IN3(n8764), .IN4(n7009), .Q(n6181)
         );
  INVX0 U8148 ( .INP(n8292), .ZN(n8972) );
  NOR2X0 U8149 ( .IN1(n9433), .IN2(n7363), .QN(n8094) );
  NAND2X0 U8150 ( .IN1(n7500), .IN2(n8727), .QN(n6174) );
  NAND2X0 U8151 ( .IN1(n6173), .IN2(n8696), .QN(n8844) );
  NAND3X0 U8152 ( .IN1(n6174), .IN2(n8844), .IN3(n8069), .QN(n6175) );
  NOR4X0 U8153 ( .IN1(n8972), .IN2(n7934), .IN3(n8094), .IN4(n6175), .QN(n6180) );
  NAND3X0 U8154 ( .IN1(n8401), .IN2(n8842), .IN3(n6510), .QN(n6176) );
  NAND3X0 U8155 ( .IN1(n9071), .IN2(n9037), .IN3(n6176), .QN(n6179) );
  NAND3X0 U8156 ( .IN1(n8921), .IN2(n7291), .IN3(n9108), .QN(n6177) );
  NAND2X0 U8157 ( .IN1(n6177), .IN2(n9125), .QN(n6178) );
  NAND4X0 U8158 ( .IN1(n6181), .IN2(n6180), .IN3(n6179), .IN4(n6178), .QN(
        \a5/N480 ) );
  NAND2X0 U8159 ( .IN1(n9190), .IN2(n9082), .QN(n7749) );
  NOR2X0 U8160 ( .IN1(n6182), .IN2(n7749), .QN(n6186) );
  OA21X1 U8161 ( .IN1(n9031), .IN2(n6755), .IN3(n9182), .Q(n6185) );
  OAI21X1 U8162 ( .IN1(n8760), .IN2(n8845), .IN3(n8962), .QN(n7217) );
  NAND2X0 U8163 ( .IN1(n9203), .IN2(n7179), .QN(n8532) );
  OR2X1 U8164 ( .IN1(n9073), .IN2(n8453), .Q(n7734) );
  NAND2X0 U8165 ( .IN1(n7355), .IN2(n8073), .QN(n6183) );
  NAND4X0 U8166 ( .IN1(n8819), .IN2(n8532), .IN3(n7734), .IN4(n6183), .QN(
        n6184) );
  NOR4X0 U8167 ( .IN1(n6186), .IN2(n6185), .IN3(n7217), .IN4(n6184), .QN(n6191) );
  INVX0 U8168 ( .INP(n6187), .ZN(n7523) );
  NAND2X0 U8169 ( .IN1(n7523), .IN2(n8026), .QN(n6189) );
  NAND4X0 U8170 ( .IN1(n6191), .IN2(n6190), .IN3(n6189), .IN4(n6188), .QN(
        \a5/N481 ) );
  OA22X1 U8171 ( .IN1(n8825), .IN2(n7316), .IN3(n8564), .IN4(n8431), .Q(n6196)
         );
  NAND2X0 U8172 ( .IN1(n8752), .IN2(n8239), .QN(n7986) );
  AND3X1 U8173 ( .IN1(n9435), .IN2(n8220), .IN3(n8675), .Q(n7611) );
  NAND2X0 U8174 ( .IN1(n7271), .IN2(n7611), .QN(n8172) );
  NAND2X0 U8175 ( .IN1(n7487), .IN2(n9438), .QN(n8838) );
  AND4X1 U8176 ( .IN1(n6800), .IN2(n7377), .IN3(n8172), .IN4(n8838), .Q(n6192)
         );
  OA221X1 U8177 ( .IN1(n7650), .IN2(n6193), .IN3(n7650), .IN4(n7986), .IN5(
        n6192), .Q(n6195) );
  NAND2X0 U8178 ( .IN1(n9105), .IN2(n7784), .QN(n8961) );
  OR2X1 U8179 ( .IN1(n8961), .IN2(n6194), .Q(n6216) );
  NAND4X0 U8180 ( .IN1(n6196), .IN2(n6195), .IN3(n8028), .IN4(n6216), .QN(
        \a5/N482 ) );
  NOR2X0 U8181 ( .IN1(n7168), .IN2(n7800), .QN(n7081) );
  INVX0 U8182 ( .INP(n7081), .ZN(n6381) );
  OA22X1 U8183 ( .IN1(n8675), .IN2(n6485), .IN3(n6936), .IN4(n6381), .Q(n6204)
         );
  AND3X1 U8184 ( .IN1(n6286), .IN2(n8834), .IN3(n8068), .Q(n6203) );
  NOR2X0 U8185 ( .IN1(n7517), .IN2(n6197), .QN(n6200) );
  NOR2X0 U8186 ( .IN1(n9434), .IN2(n8024), .QN(n6648) );
  NOR2X0 U8187 ( .IN1(n9441), .IN2(n7554), .QN(n7119) );
  AO22X1 U8188 ( .IN1(n6648), .IN2(n6198), .IN3(n7119), .IN4(n7035), .Q(n6199)
         );
  NOR4X0 U8189 ( .IN1(n8324), .IN2(n7222), .IN3(n6200), .IN4(n6199), .QN(n6202) );
  NAND4X0 U8190 ( .IN1(n6204), .IN2(n6203), .IN3(n6202), .IN4(n6201), .QN(
        \a5/N483 ) );
  AND2X1 U8191 ( .IN1(n6205), .IN2(n8880), .Q(n8471) );
  OA21X1 U8192 ( .IN1(n8471), .IN2(n8004), .IN3(n6206), .Q(n6211) );
  NAND2X0 U8193 ( .IN1(n9190), .IN2(n6207), .QN(n7334) );
  OA22X1 U8194 ( .IN1(n8667), .IN2(n8204), .IN3(n9438), .IN4(n7334), .Q(n6210)
         );
  NAND2X0 U8195 ( .IN1(n7529), .IN2(n9181), .QN(n6209) );
  NAND2X0 U8196 ( .IN1(n9435), .IN2(n8698), .QN(n6208) );
  NAND4X0 U8197 ( .IN1(n6211), .IN2(n6210), .IN3(n6209), .IN4(n6208), .QN(
        n6212) );
  NOR3X0 U8198 ( .IN1(n8606), .IN2(n6213), .IN3(n6212), .QN(n6215) );
  NAND2X0 U8199 ( .IN1(n6214), .IN2(n8496), .QN(n8965) );
  NAND4X0 U8200 ( .IN1(n6215), .IN2(n6238), .IN3(n6266), .IN4(n8965), .QN(
        \a5/N484 ) );
  OA22X1 U8201 ( .IN1(n9080), .IN2(n9165), .IN3(n9435), .IN4(n6216), .Q(n6224)
         );
  NOR2X0 U8202 ( .IN1(n8649), .IN2(n6811), .QN(n7002) );
  NOR2X0 U8203 ( .IN1(n9001), .IN2(n9029), .QN(n6219) );
  NAND3X0 U8204 ( .IN1(n7445), .IN2(n8747), .IN3(n6217), .QN(n6218) );
  NOR4X0 U8205 ( .IN1(n8855), .IN2(n7002), .IN3(n6219), .IN4(n6218), .QN(n6223) );
  NAND2X0 U8206 ( .IN1(degrees_tmp2[3]), .IN2(n6220), .QN(n7769) );
  NAND2X0 U8207 ( .IN1(n6221), .IN2(n8787), .QN(n6222) );
  NAND4X0 U8208 ( .IN1(n6224), .IN2(n6223), .IN3(n7769), .IN4(n6222), .QN(
        \a5/N485 ) );
  OA21X1 U8209 ( .IN1(n9053), .IN2(n9045), .IN3(n7722), .Q(n6228) );
  NOR2X0 U8210 ( .IN1(n9435), .IN2(n8069), .QN(n8923) );
  AO221X1 U8211 ( .IN1(n9080), .IN2(n8529), .IN3(n9080), .IN4(n6668), .IN5(
        n8923), .Q(n6225) );
  NOR4X0 U8212 ( .IN1(n7645), .IN2(n9066), .IN3(n7408), .IN4(n6225), .QN(n6227) );
  NAND2X0 U8213 ( .IN1(n7858), .IN2(n9099), .QN(n6226) );
  NAND4X0 U8214 ( .IN1(n6228), .IN2(n6227), .IN3(n6321), .IN4(n6226), .QN(
        \a5/N486 ) );
  NAND2X0 U8215 ( .IN1(n7421), .IN2(n8822), .QN(n8382) );
  NAND2X0 U8216 ( .IN1(n8731), .IN2(n7956), .QN(n6229) );
  OR2X1 U8217 ( .IN1(n9061), .IN2(n7431), .Q(n8125) );
  AND4X1 U8218 ( .IN1(n9165), .IN2(n8382), .IN3(n6229), .IN4(n8125), .Q(n6230)
         );
  NAND2X0 U8219 ( .IN1(n8796), .IN2(n6665), .QN(n8776) );
  NAND4X0 U8220 ( .IN1(n6230), .IN2(n6845), .IN3(n8339), .IN4(n8776), .QN(
        \a5/N487 ) );
  NOR3X0 U8221 ( .IN1(n9037), .IN2(n6797), .IN3(n6893), .QN(n6232) );
  NOR2X0 U8222 ( .IN1(n6232), .IN2(n6231), .QN(n7420) );
  INVX0 U8223 ( .INP(n7754), .ZN(n8203) );
  NAND3X0 U8224 ( .IN1(n7420), .IN2(n8203), .IN3(n8217), .QN(\a5/N488 ) );
  NAND2X0 U8225 ( .IN1(degrees_tmp2[3]), .IN2(n7582), .QN(n6233) );
  NAND3X0 U8226 ( .IN1(n8218), .IN2(n6233), .IN3(n8217), .QN(\a5/N489 ) );
  OR2X1 U8227 ( .IN1(\a5/N491 ), .IN2(n8718), .Q(\a5/N490 ) );
  INVX0 U8228 ( .INP(n6234), .ZN(\a3/N492 ) );
  NOR2X0 U8229 ( .IN1(n9054), .IN2(n7534), .QN(n6242) );
  INVX0 U8230 ( .INP(n8748), .ZN(n7889) );
  AO22X1 U8231 ( .IN1(n8822), .IN2(n7858), .IN3(degrees_tmp2[3]), .IN4(n7889), 
        .Q(n6241) );
  NAND2X0 U8232 ( .IN1(n6235), .IN2(n7271), .QN(n8610) );
  INVX0 U8233 ( .INP(n8610), .ZN(n6236) );
  NOR2X0 U8234 ( .IN1(n8288), .IN2(n7009), .QN(n6708) );
  NOR4X0 U8235 ( .IN1(n7653), .IN2(n8257), .IN3(n6236), .IN4(n6708), .QN(n6239) );
  NAND4X0 U8236 ( .IN1(n9190), .IN2(n9438), .IN3(n9436), .IN4(n7597), .QN(
        n7673) );
  AO21X1 U8237 ( .IN1(n7600), .IN2(n6408), .IN3(n7969), .Q(n6237) );
  NAND4X0 U8238 ( .IN1(n6239), .IN2(n6238), .IN3(n7673), .IN4(n6237), .QN(
        n6240) );
  NOR4X0 U8239 ( .IN1(n6352), .IN2(n6242), .IN3(n6241), .IN4(n6240), .QN(n6245) );
  INVX0 U8240 ( .INP(n7063), .ZN(n8551) );
  NAND2X0 U8241 ( .IN1(n6243), .IN2(n7236), .QN(n9139) );
  NAND3X0 U8242 ( .IN1(n8760), .IN2(n8186), .IN3(n8474), .QN(n6244) );
  NAND4X0 U8243 ( .IN1(n6245), .IN2(n8551), .IN3(n9139), .IN4(n6244), .QN(
        \a4/N436 ) );
  OA21X1 U8244 ( .IN1(n6461), .IN2(n7678), .IN3(n8431), .Q(n6253) );
  AND3X1 U8245 ( .IN1(degrees_tmp2[0]), .IN2(n8655), .IN3(n8886), .Q(n6252) );
  NAND2X0 U8246 ( .IN1(n7698), .IN2(n8467), .QN(n6248) );
  NAND2X0 U8247 ( .IN1(n6246), .IN2(n8780), .QN(n6247) );
  NAND4X0 U8248 ( .IN1(n6474), .IN2(n7786), .IN3(n6248), .IN4(n6247), .QN(
        n6251) );
  NAND3X0 U8249 ( .IN1(n8529), .IN2(n8995), .IN3(n7745), .QN(n8280) );
  NAND4X0 U8250 ( .IN1(n8280), .IN2(n8135), .IN3(n6249), .IN4(n8885), .QN(
        n6250) );
  NOR4X0 U8251 ( .IN1(n6253), .IN2(n6252), .IN3(n6251), .IN4(n6250), .QN(n6255) );
  INVX0 U8252 ( .INP(n8077), .ZN(n8231) );
  NAND4X0 U8253 ( .IN1(n6255), .IN2(n8231), .IN3(n7781), .IN4(n6254), .QN(
        \a4/N437 ) );
  INVX0 U8254 ( .INP(n7236), .ZN(n9083) );
  OA22X1 U8255 ( .IN1(n7766), .IN2(n8282), .IN3(n7571), .IN4(n9083), .Q(n6263)
         );
  NOR2X0 U8256 ( .IN1(n6256), .IN2(n8568), .QN(n6287) );
  NAND2X0 U8257 ( .IN1(n6287), .IN2(n6979), .QN(n7368) );
  NOR2X0 U8258 ( .IN1(degrees_tmp2[2]), .IN2(n7368), .QN(n8659) );
  NOR2X0 U8259 ( .IN1(n8572), .IN2(n7834), .QN(n6260) );
  OR2X1 U8260 ( .IN1(n6257), .IN2(n8124), .Q(n6258) );
  NAND4X0 U8261 ( .IN1(n8835), .IN2(n8039), .IN3(n7891), .IN4(n6258), .QN(
        n6259) );
  NOR4X0 U8262 ( .IN1(n8324), .IN2(n8659), .IN3(n6260), .IN4(n6259), .QN(n6262) );
  NAND2X0 U8263 ( .IN1(n6261), .IN2(n7012), .QN(n8117) );
  NAND4X0 U8264 ( .IN1(n6263), .IN2(n6262), .IN3(n7743), .IN4(n8117), .QN(
        \a4/N439 ) );
  OA22X1 U8265 ( .IN1(n8881), .IN2(n8317), .IN3(n9445), .IN4(n6264), .Q(n6267)
         );
  NAND3X0 U8266 ( .IN1(n9435), .IN2(n8675), .IN3(n8354), .QN(n6265) );
  NAND4X0 U8267 ( .IN1(n6267), .IN2(n6266), .IN3(n7118), .IN4(n6265), .QN(
        n6270) );
  NOR2X0 U8268 ( .IN1(n7358), .IN2(n8472), .QN(n7543) );
  NAND2X0 U8269 ( .IN1(n6268), .IN2(n6920), .QN(n7022) );
  INVX0 U8270 ( .INP(n6909), .ZN(n7204) );
  NAND2X0 U8271 ( .IN1(n9435), .IN2(n7204), .QN(n7890) );
  NAND4X0 U8272 ( .IN1(n7543), .IN2(n7862), .IN3(n7022), .IN4(n7890), .QN(
        n6269) );
  NOR2X0 U8273 ( .IN1(n6270), .IN2(n6269), .QN(n6272) );
  NAND2X0 U8274 ( .IN1(n8978), .IN2(n6271), .QN(n9118) );
  NAND4X0 U8275 ( .IN1(n6273), .IN2(n6272), .IN3(n8172), .IN4(n9118), .QN(
        \a4/N440 ) );
  NOR2X0 U8276 ( .IN1(n7736), .IN2(n7168), .QN(n6569) );
  NAND2X0 U8277 ( .IN1(degrees_tmp2[0]), .IN2(n6569), .QN(n6689) );
  NAND2X0 U8278 ( .IN1(n8876), .IN2(n6365), .QN(n7181) );
  NAND4X0 U8279 ( .IN1(n6985), .IN2(n7787), .IN3(n6689), .IN4(n7181), .QN(
        n6282) );
  NAND2X0 U8280 ( .IN1(n6274), .IN2(n8073), .QN(n6278) );
  NAND2X0 U8281 ( .IN1(n7615), .IN2(n6275), .QN(n6276) );
  NAND4X0 U8282 ( .IN1(n6278), .IN2(n8514), .IN3(n6277), .IN4(n6276), .QN(
        n6281) );
  NAND2X0 U8283 ( .IN1(n8727), .IN2(n9005), .QN(n8054) );
  NAND3X0 U8284 ( .IN1(n7208), .IN2(n7389), .IN3(n9442), .QN(n6279) );
  NAND4X0 U8285 ( .IN1(n8183), .IN2(n8590), .IN3(n8054), .IN4(n6279), .QN(
        n6280) );
  NOR4X0 U8286 ( .IN1(n6283), .IN2(n6282), .IN3(n6281), .IN4(n6280), .QN(n6285) );
  NAND2X0 U8287 ( .IN1(n8529), .IN2(n7233), .QN(n8381) );
  NOR2X0 U8288 ( .IN1(n9434), .IN2(n8381), .QN(n7338) );
  NAND2X0 U8289 ( .IN1(n7338), .IN2(n9436), .QN(n6390) );
  NAND3X0 U8290 ( .IN1(n7413), .IN2(n9122), .IN3(n8938), .QN(n6284) );
  NAND3X0 U8291 ( .IN1(n6285), .IN2(n6390), .IN3(n6284), .QN(\a4/N441 ) );
  OA22X1 U8292 ( .IN1(n8825), .IN2(n8610), .IN3(n7174), .IN4(n9099), .Q(n6295)
         );
  NOR2X0 U8293 ( .IN1(n8489), .IN2(n6371), .QN(n7203) );
  NAND2X0 U8294 ( .IN1(n8169), .IN2(n6286), .QN(n6872) );
  NAND2X0 U8295 ( .IN1(n7784), .IN2(n6872), .QN(n8554) );
  INVX0 U8296 ( .INP(n8554), .ZN(n6288) );
  OA21X1 U8297 ( .IN1(n6288), .IN2(n6287), .IN3(n9442), .Q(n6291) );
  AND2X1 U8298 ( .IN1(n8724), .IN2(n9150), .Q(n6290) );
  NOR4X0 U8299 ( .IN1(n7203), .IN2(n6291), .IN3(n6290), .IN4(n6289), .QN(n6294) );
  NAND2X0 U8300 ( .IN1(n8424), .IN2(n6296), .QN(n8857) );
  INVX0 U8301 ( .INP(n6292), .ZN(n8507) );
  AO22X1 U8302 ( .IN1(n8124), .IN2(n9061), .IN3(n7467), .IN4(n8507), .Q(n6293)
         );
  NAND4X0 U8303 ( .IN1(n6295), .IN2(n6294), .IN3(n8857), .IN4(n6293), .QN(
        \a4/N442 ) );
  NAND2X0 U8304 ( .IN1(n6296), .IN2(n8026), .QN(n6931) );
  NOR2X0 U8305 ( .IN1(n8431), .IN2(n6931), .QN(n7139) );
  NOR2X0 U8306 ( .IN1(n7414), .IN2(n7281), .QN(n7023) );
  NOR2X0 U8307 ( .IN1(n7023), .IN2(n8692), .QN(n6302) );
  NAND2X0 U8308 ( .IN1(n9434), .IN2(n6453), .QN(n9160) );
  NAND3X0 U8309 ( .IN1(n6826), .IN2(n9031), .IN3(n8787), .QN(n6297) );
  NAND4X0 U8310 ( .IN1(n9160), .IN2(n9111), .IN3(n8892), .IN4(n6297), .QN(
        n6301) );
  NAND2X0 U8311 ( .IN1(n6649), .IN2(n8534), .QN(n8927) );
  NAND3X0 U8312 ( .IN1(n8699), .IN2(n7169), .IN3(n7093), .QN(n8291) );
  NAND2X0 U8313 ( .IN1(n8786), .IN2(n7800), .QN(n6299) );
  NAND4X0 U8314 ( .IN1(n8927), .IN2(n8291), .IN3(n6299), .IN4(n6298), .QN(
        n6300) );
  NOR4X0 U8315 ( .IN1(n7139), .IN2(n6302), .IN3(n6301), .IN4(n6300), .QN(n6304) );
  NAND2X0 U8316 ( .IN1(degrees_tmp2[0]), .IN2(n7900), .QN(n6303) );
  NAND4X0 U8317 ( .IN1(n7926), .IN2(n6304), .IN3(n6303), .IN4(n7558), .QN(
        \a4/N443 ) );
  AOI22X1 U8318 ( .IN1(n9092), .IN2(n8760), .IN3(n7312), .IN4(n7035), .QN(
        n6319) );
  INVX0 U8319 ( .INP(n6305), .ZN(n6317) );
  NOR2X0 U8320 ( .IN1(n8572), .IN2(n6811), .QN(n6316) );
  NOR2X0 U8321 ( .IN1(n8022), .IN2(n6306), .QN(n6307) );
  NOR2X0 U8322 ( .IN1(n7342), .IN2(n6307), .QN(n6310) );
  NAND2X0 U8323 ( .IN1(n9435), .IN2(n8180), .QN(n9022) );
  AND2X1 U8324 ( .IN1(n6308), .IN2(n9022), .Q(n6309) );
  OA22X1 U8325 ( .IN1(n6310), .IN2(n8568), .IN3(n6309), .IN4(n9149), .Q(n6314)
         );
  NAND2X0 U8326 ( .IN1(n9189), .IN2(n9195), .QN(n7287) );
  OA22X1 U8327 ( .IN1(n8816), .IN2(n7287), .IN3(n7517), .IN4(n6311), .Q(n6313)
         );
  INVX0 U8328 ( .INP(n6835), .ZN(n9010) );
  NAND2X0 U8329 ( .IN1(n6650), .IN2(n9010), .QN(n7345) );
  NAND4X0 U8330 ( .IN1(n6314), .IN2(n6313), .IN3(n6312), .IN4(n7345), .QN(
        n6315) );
  NOR4X0 U8331 ( .IN1(n8972), .IN2(n6317), .IN3(n6316), .IN4(n6315), .QN(n6318) );
  NAND4X0 U8332 ( .IN1(n6319), .IN2(n6318), .IN3(n8821), .IN4(n9050), .QN(
        \a4/N444 ) );
  NOR2X0 U8333 ( .IN1(n8978), .IN2(n8761), .QN(n6332) );
  NAND2X0 U8334 ( .IN1(n6320), .IN2(n9122), .QN(n6955) );
  NAND4X0 U8335 ( .IN1(n7771), .IN2(n7363), .IN3(n6955), .IN4(n6321), .QN(
        n6331) );
  OA22X1 U8336 ( .IN1(n8249), .IN2(n6464), .IN3(n6323), .IN4(n6322), .Q(n6324)
         );
  OA221X1 U8337 ( .IN1(n8728), .IN2(n8104), .IN3(n8728), .IN4(n6996), .IN5(
        n6324), .Q(n6329) );
  NAND2X0 U8338 ( .IN1(n7945), .IN2(n9032), .QN(n7238) );
  NAND2X0 U8339 ( .IN1(n6325), .IN2(n7238), .QN(n7860) );
  NAND2X0 U8340 ( .IN1(n6327), .IN2(n6326), .QN(n6328) );
  NAND4X0 U8341 ( .IN1(n6329), .IN2(n7730), .IN3(n7860), .IN4(n6328), .QN(
        n6330) );
  OR4X1 U8342 ( .IN1(n6333), .IN2(n6332), .IN3(n6331), .IN4(n6330), .Q(
        \a4/N445 ) );
  OA21X1 U8343 ( .IN1(n8575), .IN2(n9129), .IN3(n8799), .Q(n6340) );
  NAND2X0 U8344 ( .IN1(n6623), .IN2(n9147), .QN(n6794) );
  OA22X1 U8345 ( .IN1(n7766), .IN2(n8588), .IN3(n7745), .IN4(n6794), .Q(n6336)
         );
  NAND3X0 U8346 ( .IN1(n8315), .IN2(n8545), .IN3(n8882), .QN(n6334) );
  NAND2X0 U8347 ( .IN1(n6334), .IN2(n8796), .QN(n6335) );
  AND4X1 U8348 ( .IN1(n6336), .IN2(n7981), .IN3(n8226), .IN4(n6335), .Q(n6339)
         );
  AO21X1 U8349 ( .IN1(n9002), .IN2(n6337), .IN3(n8724), .Q(n6338) );
  NAND4X0 U8350 ( .IN1(n6340), .IN2(n6339), .IN3(n8470), .IN4(n6338), .QN(
        \a4/N446 ) );
  OA22X1 U8351 ( .IN1(n6342), .IN2(n8922), .IN3(degrees_tmp2[0]), .IN4(n6341), 
        .Q(n6350) );
  INVX0 U8352 ( .INP(n6343), .ZN(n6351) );
  OA22X1 U8353 ( .IN1(n9053), .IN2(n6351), .IN3(n8527), .IN4(n7238), .Q(n6349)
         );
  NOR2X0 U8354 ( .IN1(n8728), .IN2(n9127), .QN(n8560) );
  INVX0 U8355 ( .INP(n8937), .ZN(n6344) );
  NAND2X0 U8356 ( .IN1(n6344), .IN2(n6403), .QN(n8396) );
  NAND4X0 U8357 ( .IN1(n8336), .IN2(n7499), .IN3(n8776), .IN4(n8396), .QN(
        n6346) );
  AO22X1 U8358 ( .IN1(n8760), .IN2(n6660), .IN3(n7437), .IN4(n6584), .Q(n6345)
         );
  NOR4X0 U8359 ( .IN1(n6347), .IN2(n8560), .IN3(n6346), .IN4(n6345), .QN(n6348) );
  NAND4X0 U8360 ( .IN1(n6350), .IN2(n6349), .IN3(n6348), .IN4(n8292), .QN(
        \a4/N447 ) );
  NOR2X0 U8361 ( .IN1(n7510), .IN2(n6351), .QN(n6354) );
  NOR3X0 U8362 ( .IN1(n6354), .IN2(n6353), .IN3(n6352), .QN(n6364) );
  NOR2X0 U8363 ( .IN1(n7517), .IN2(n8587), .QN(n6358) );
  NOR2X0 U8364 ( .IN1(n9183), .IN2(n8751), .QN(n6357) );
  NOR2X0 U8365 ( .IN1(n7652), .IN2(n8654), .QN(n8296) );
  NAND4X0 U8366 ( .IN1(n8296), .IN2(n9041), .IN3(n6669), .IN4(n6355), .QN(
        n6356) );
  NOR4X0 U8367 ( .IN1(n6359), .IN2(n6358), .IN3(n6357), .IN4(n6356), .QN(n6363) );
  INVX0 U8368 ( .INP(n6360), .ZN(n8815) );
  AO21X1 U8369 ( .IN1(n8815), .IN2(n6361), .IN3(n9435), .Q(n6362) );
  NAND4X0 U8370 ( .IN1(n6364), .IN2(n6363), .IN3(n8099), .IN4(n6362), .QN(
        \a4/N448 ) );
  NAND2X0 U8371 ( .IN1(n6365), .IN2(n7656), .QN(n6368) );
  NAND3X0 U8372 ( .IN1(n7093), .IN2(n6366), .IN3(n7462), .QN(n6367) );
  AND3X1 U8373 ( .IN1(n7099), .IN2(n6368), .IN3(n6367), .Q(n6380) );
  NOR2X0 U8374 ( .IN1(n7168), .IN2(n6369), .QN(n9117) );
  NOR2X0 U8375 ( .IN1(n6371), .IN2(n6370), .QN(n8924) );
  NAND4X0 U8376 ( .IN1(n8314), .IN2(n6372), .IN3(n8807), .IN4(n7330), .QN(
        n6378) );
  NAND2X0 U8377 ( .IN1(n8826), .IN2(n9189), .QN(n6374) );
  OA22X1 U8378 ( .IN1(n8247), .IN2(n6374), .IN3(n7913), .IN4(n6373), .Q(n6376)
         );
  NAND4X0 U8379 ( .IN1(n6376), .IN2(n7107), .IN3(n8889), .IN4(n6375), .QN(
        n6377) );
  NOR4X0 U8380 ( .IN1(n9117), .IN2(n8924), .IN3(n6378), .IN4(n6377), .QN(n6379) );
  NAND4X0 U8381 ( .IN1(n6380), .IN2(n6379), .IN3(n7459), .IN4(n8070), .QN(
        \a4/N449 ) );
  INVX0 U8382 ( .INP(n6936), .ZN(n7878) );
  OA22X1 U8383 ( .IN1(n8978), .IN2(n8939), .IN3(n6381), .IN4(n7878), .Q(n6389)
         );
  INVX0 U8384 ( .INP(n6382), .ZN(n8411) );
  NAND2X0 U8385 ( .IN1(n8866), .IN2(n8411), .QN(n7263) );
  INVX0 U8386 ( .INP(n6914), .ZN(n7851) );
  OA21X1 U8387 ( .IN1(n6606), .IN2(n6635), .IN3(n7851), .Q(n6386) );
  OA22X1 U8388 ( .IN1(n9082), .IN2(n8859), .IN3(n9031), .IN4(n6773), .Q(n6385)
         );
  NAND2X0 U8389 ( .IN1(n7533), .IN2(n7251), .QN(n6383) );
  NAND3X0 U8390 ( .IN1(n6383), .IN2(n7717), .IN3(n8675), .QN(n6384) );
  NAND4X0 U8391 ( .IN1(n6386), .IN2(n6385), .IN3(n8244), .IN4(n6384), .QN(
        n6387) );
  NOR4X0 U8392 ( .IN1(n6745), .IN2(n8654), .IN3(n7263), .IN4(n6387), .QN(n6388) );
  NAND4X0 U8393 ( .IN1(n6389), .IN2(n6388), .IN3(n8613), .IN4(n8571), .QN(
        \a4/N450 ) );
  NAND2X0 U8394 ( .IN1(n6569), .IN2(n8787), .QN(n6883) );
  OA22X1 U8395 ( .IN1(n9438), .IN2(n6883), .IN3(n9128), .IN4(n7596), .Q(n6397)
         );
  AOI22X1 U8396 ( .IN1(n7133), .IN2(n8431), .IN3(n8676), .IN4(n8568), .QN(
        n6396) );
  OA221X1 U8397 ( .IN1(n8229), .IN2(n6908), .IN3(n8229), .IN4(n8410), .IN5(
        n6390), .Q(n6395) );
  AND3X1 U8398 ( .IN1(n6649), .IN2(n9195), .IN3(n9166), .Q(n7160) );
  AND3X1 U8399 ( .IN1(n6392), .IN2(n9435), .IN3(n6391), .Q(n6646) );
  NOR4X0 U8400 ( .IN1(n6771), .IN2(n6393), .IN3(n7160), .IN4(n6646), .QN(n6394) );
  NAND4X0 U8401 ( .IN1(n6397), .IN2(n6396), .IN3(n6395), .IN4(n6394), .QN(
        \a4/N451 ) );
  INVX0 U8402 ( .INP(n9126), .ZN(n6861) );
  NOR2X0 U8403 ( .IN1(n6398), .IN2(n8987), .QN(n7129) );
  AO22X1 U8404 ( .IN1(n8883), .IN2(n7161), .IN3(n6399), .IN4(n7402), .Q(n6400)
         );
  NOR4X0 U8405 ( .IN1(n9014), .IN2(n6861), .IN3(n7129), .IN4(n6400), .QN(n6411) );
  NOR2X0 U8406 ( .IN1(n6401), .IN2(n6553), .QN(n7693) );
  INVX0 U8407 ( .INP(n6402), .ZN(n6407) );
  INVX0 U8408 ( .INP(n7183), .ZN(n6516) );
  AOI22X1 U8409 ( .IN1(n7198), .IN2(n6403), .IN3(n6516), .IN4(n7745), .QN(
        n6405) );
  NAND4X0 U8410 ( .IN1(n6405), .IN2(n6404), .IN3(n6982), .IN4(n8265), .QN(
        n6406) );
  NOR4X0 U8411 ( .IN1(n7693), .IN2(n6407), .IN3(n7681), .IN4(n6406), .QN(n6410) );
  NAND2X0 U8412 ( .IN1(n6667), .IN2(n9440), .QN(n7127) );
  NOR2X0 U8413 ( .IN1(degrees_tmp2[2]), .IN2(n6408), .QN(n8662) );
  NAND2X0 U8414 ( .IN1(n8754), .IN2(n8662), .QN(n6409) );
  NAND4X0 U8415 ( .IN1(n6411), .IN2(n6410), .IN3(n7127), .IN4(n6409), .QN(
        \a4/N452 ) );
  NAND4X0 U8416 ( .IN1(n9437), .IN2(n9435), .IN3(n6412), .IN4(n9440), .QN(
        n8829) );
  NAND2X0 U8417 ( .IN1(n8829), .IN2(n6723), .QN(n7231) );
  NOR2X0 U8418 ( .IN1(n9435), .IN2(n7600), .QN(n7436) );
  NAND2X0 U8419 ( .IN1(n7436), .IN2(n9445), .QN(n7024) );
  NAND4X0 U8420 ( .IN1(n6414), .IN2(n7024), .IN3(n6413), .IN4(n7730), .QN(
        n6415) );
  NOR4X0 U8421 ( .IN1(n6528), .IN2(n6416), .IN3(n7231), .IN4(n6415), .QN(n6424) );
  NOR2X0 U8422 ( .IN1(n9188), .IN2(n7501), .QN(n6419) );
  NAND2X0 U8423 ( .IN1(n8886), .IN2(n6417), .QN(n6418) );
  NAND2X0 U8424 ( .IN1(n6419), .IN2(n6418), .QN(n6420) );
  NAND2X0 U8425 ( .IN1(n8760), .IN2(n6420), .QN(n6423) );
  NAND2X0 U8426 ( .IN1(n8239), .IN2(n8886), .QN(n8781) );
  AO21X1 U8427 ( .IN1(n8922), .IN2(n8781), .IN3(n8282), .Q(n6422) );
  NAND2X0 U8428 ( .IN1(n8710), .IN2(n8305), .QN(n6421) );
  NAND4X0 U8429 ( .IN1(n6424), .IN2(n6423), .IN3(n6422), .IN4(n6421), .QN(
        \a4/N453 ) );
  INVX0 U8430 ( .INP(n7165), .ZN(n6425) );
  NOR2X0 U8431 ( .IN1(n6425), .IN2(n9065), .QN(n8037) );
  INVX0 U8432 ( .INP(n8845), .ZN(n9175) );
  NAND3X0 U8433 ( .IN1(n9175), .IN2(n8004), .IN3(n7473), .QN(n7718) );
  OA21X1 U8434 ( .IN1(n6454), .IN2(n6426), .IN3(n7718), .Q(n6432) );
  NOR2X0 U8435 ( .IN1(n7473), .IN2(n7881), .QN(n6430) );
  NOR2X0 U8436 ( .IN1(n6427), .IN2(n8001), .QN(n8943) );
  NAND2X0 U8437 ( .IN1(n6614), .IN2(n8943), .QN(n6628) );
  NAND4X0 U8438 ( .IN1(n8167), .IN2(n7362), .IN3(n8859), .IN4(n6628), .QN(
        n6429) );
  AO22X1 U8439 ( .IN1(n7654), .IN2(n8692), .IN3(n7033), .IN4(n7800), .Q(n6428)
         );
  NOR4X0 U8440 ( .IN1(n9066), .IN2(n6430), .IN3(n6429), .IN4(n6428), .QN(n6431) );
  NAND2X0 U8441 ( .IN1(n7133), .IN2(n9436), .QN(n7747) );
  NAND4X0 U8442 ( .IN1(n8037), .IN2(n6432), .IN3(n6431), .IN4(n7747), .QN(
        \a4/N454 ) );
  NOR2X0 U8443 ( .IN1(degrees_tmp2[2]), .IN2(n6433), .QN(n7031) );
  NAND2X0 U8444 ( .IN1(n8379), .IN2(n9433), .QN(n7443) );
  NAND2X0 U8445 ( .IN1(n6434), .IN2(n6647), .QN(n7224) );
  INVX0 U8446 ( .INP(n6567), .ZN(n7360) );
  NAND2X0 U8447 ( .IN1(n7360), .IN2(n9122), .QN(n6435) );
  NAND4X0 U8448 ( .IN1(n7509), .IN2(n7443), .IN3(n7224), .IN4(n6435), .QN(
        n6447) );
  NAND2X0 U8449 ( .IN1(n8598), .IN2(n9187), .QN(n6436) );
  NAND4X0 U8450 ( .IN1(n9165), .IN2(n8029), .IN3(n6437), .IN4(n6436), .QN(
        n6446) );
  NOR2X0 U8451 ( .IN1(n6780), .IN2(n6438), .QN(n6439) );
  OA22X1 U8452 ( .IN1(degrees_tmp2[2]), .IN2(n6440), .IN3(n6439), .IN4(n8724), 
        .Q(n6444) );
  OA21X1 U8453 ( .IN1(n6614), .IN2(n6441), .IN3(n7494), .Q(n6443) );
  NAND4X0 U8454 ( .IN1(n6444), .IN2(n6443), .IN3(n6442), .IN4(n6524), .QN(
        n6445) );
  OR4X1 U8455 ( .IN1(n7031), .IN2(n6447), .IN3(n6446), .IN4(n6445), .Q(
        \a4/N455 ) );
  INVX0 U8456 ( .INP(n8410), .ZN(n8393) );
  NOR2X0 U8457 ( .IN1(n7168), .IN2(n9046), .QN(n6460) );
  OA21X1 U8458 ( .IN1(n6449), .IN2(n6448), .IN3(n8531), .Q(n6459) );
  NOR2X0 U8459 ( .IN1(degrees_tmp2[2]), .IN2(n6450), .QN(n6452) );
  NOR2X0 U8460 ( .IN1(n6452), .IN2(n6451), .QN(n6457) );
  INVX0 U8461 ( .INP(n6453), .ZN(n6847) );
  NAND3X0 U8462 ( .IN1(n6454), .IN2(n8384), .IN3(n6847), .QN(n6455) );
  NAND2X0 U8463 ( .IN1(n9440), .IN2(n6455), .QN(n6456) );
  NAND2X0 U8464 ( .IN1(n6457), .IN2(n6456), .QN(n6458) );
  NOR4X0 U8465 ( .IN1(n8393), .IN2(n6460), .IN3(n6459), .IN4(n6458), .QN(n6463) );
  NAND2X0 U8466 ( .IN1(n6461), .IN2(n8649), .QN(n6462) );
  NAND4X0 U8467 ( .IN1(n6463), .IN2(n6739), .IN3(n6462), .IN4(n8926), .QN(
        \a4/N456 ) );
  OA222X1 U8468 ( .IN1(n9122), .IN2(n8071), .IN3(n9122), .IN4(n6464), .IN5(
        n8533), .IN6(n8156), .Q(n6472) );
  NOR3X0 U8469 ( .IN1(n8320), .IN2(n9075), .IN3(n7500), .QN(n6465) );
  OA22X1 U8470 ( .IN1(n8883), .IN2(n7259), .IN3(n6465), .IN4(n9181), .Q(n6471)
         );
  INVX0 U8471 ( .INP(n6814), .ZN(n6467) );
  NOR2X0 U8472 ( .IN1(n7656), .IN2(n6466), .QN(n7264) );
  NOR4X0 U8473 ( .IN1(n6914), .IN2(n6467), .IN3(n7804), .IN4(n7264), .QN(n6470) );
  NAND2X0 U8474 ( .IN1(degrees_tmp2[0]), .IN2(n8408), .QN(n8025) );
  AND2X1 U8475 ( .IN1(n8025), .IN2(n7369), .Q(n8870) );
  NOR2X0 U8476 ( .IN1(n9435), .IN2(n8870), .QN(n6468) );
  NOR4X0 U8477 ( .IN1(n7192), .IN2(n6862), .IN3(n8178), .IN4(n6468), .QN(n6469) );
  NAND4X0 U8478 ( .IN1(n6472), .IN2(n6471), .IN3(n6470), .IN4(n6469), .QN(
        \a4/N457 ) );
  INVX0 U8479 ( .INP(n8163), .ZN(n6473) );
  NOR2X0 U8480 ( .IN1(n6968), .IN2(n6473), .QN(n6719) );
  NOR2X0 U8481 ( .IN1(n9445), .IN2(n6903), .QN(n6480) );
  OR2X1 U8482 ( .IN1(n8979), .IN2(n9073), .Q(n8136) );
  OA22X1 U8483 ( .IN1(n9031), .IN2(n8136), .IN3(degrees_tmp2[3]), .IN4(n6878), 
        .Q(n6478) );
  AO22X1 U8484 ( .IN1(n8693), .IN2(n6497), .IN3(n9436), .IN4(n6474), .Q(n6477)
         );
  NAND3X0 U8485 ( .IN1(degrees_tmp2[3]), .IN2(n7437), .IN3(n7254), .QN(n7104)
         );
  NAND2X0 U8486 ( .IN1(n9437), .IN2(n6475), .QN(n6476) );
  NAND4X0 U8487 ( .IN1(n6478), .IN2(n6477), .IN3(n7104), .IN4(n6476), .QN(
        n6479) );
  NOR4X0 U8488 ( .IN1(n6481), .IN2(n6719), .IN3(n6480), .IN4(n6479), .QN(n6484) );
  INVX0 U8489 ( .INP(n6865), .ZN(n8402) );
  NAND2X0 U8490 ( .IN1(n7921), .IN2(n8041), .QN(n7265) );
  INVX0 U8491 ( .INP(n7417), .ZN(n7403) );
  NAND2X0 U8492 ( .IN1(n9047), .IN2(n7403), .QN(n9109) );
  NAND4X0 U8493 ( .IN1(n8597), .IN2(n8903), .IN3(n8596), .IN4(n9109), .QN(
        n6482) );
  NAND2X0 U8494 ( .IN1(n7169), .IN2(n6482), .QN(n6483) );
  NAND4X0 U8495 ( .IN1(n6484), .IN2(n8402), .IN3(n7265), .IN4(n6483), .QN(
        \a4/N458 ) );
  NOR2X0 U8496 ( .IN1(n8675), .IN2(n6485), .QN(n6486) );
  NAND2X0 U8497 ( .IN1(n6737), .IN2(n9433), .QN(n8856) );
  INVX0 U8498 ( .INP(n8856), .ZN(n8953) );
  NOR4X0 U8499 ( .IN1(n6487), .IN2(n8310), .IN3(n6486), .IN4(n8953), .QN(n6496) );
  NOR2X0 U8500 ( .IN1(n9434), .IN2(n6488), .QN(n7277) );
  NAND3X0 U8501 ( .IN1(n9105), .IN2(n9125), .IN3(n9183), .QN(n8733) );
  NAND4X0 U8502 ( .IN1(n8193), .IN2(n8099), .IN3(n8733), .IN4(n7307), .QN(
        n6491) );
  AO22X1 U8503 ( .IN1(degrees_tmp2[2]), .IN2(n7311), .IN3(n8461), .IN4(n6489), 
        .Q(n6490) );
  NOR4X0 U8504 ( .IN1(n6492), .IN2(n7277), .IN3(n6491), .IN4(n6490), .QN(n6495) );
  NAND3X0 U8505 ( .IN1(n9031), .IN2(n6493), .IN3(n8034), .QN(n6494) );
  NAND4X0 U8506 ( .IN1(n6496), .IN2(n6495), .IN3(n6669), .IN4(n6494), .QN(
        \a4/N460 ) );
  OA22X1 U8507 ( .IN1(n9208), .IN2(n6497), .IN3(n9122), .IN4(n8527), .Q(n6506)
         );
  NOR2X0 U8508 ( .IN1(n8948), .IN2(n6974), .QN(n6498) );
  OA22X1 U8509 ( .IN1(n9084), .IN2(n6498), .IN3(n7766), .IN4(n8649), .Q(n6501)
         );
  NAND3X0 U8510 ( .IN1(n9105), .IN2(n9183), .IN3(n9433), .QN(n6499) );
  NAND4X0 U8511 ( .IN1(n6501), .IN2(n6500), .IN3(n8747), .IN4(n6499), .QN(
        n6502) );
  NOR4X0 U8512 ( .IN1(n7081), .IN2(n6503), .IN3(n9066), .IN4(n6502), .QN(n6505) );
  INVX0 U8513 ( .INP(n6504), .ZN(n8555) );
  NAND3X0 U8514 ( .IN1(n6506), .IN2(n6505), .IN3(n8555), .QN(\a4/N461 ) );
  INVX0 U8515 ( .INP(n7108), .ZN(n8157) );
  OA22X1 U8516 ( .IN1(n9071), .IN2(n8882), .IN3(n6979), .IN4(n8157), .Q(n6519)
         );
  INVX0 U8517 ( .INP(n8819), .ZN(n6791) );
  NOR2X0 U8518 ( .IN1(n8995), .IN2(n8244), .QN(n6515) );
  NOR2X0 U8519 ( .IN1(n6508), .IN2(n6507), .QN(n6511) );
  OA22X1 U8520 ( .IN1(n6511), .IN2(n6510), .IN3(n7679), .IN4(n6509), .Q(n6513)
         );
  NAND2X0 U8521 ( .IN1(n6781), .IN2(n9440), .QN(n7612) );
  NAND2X0 U8522 ( .IN1(n8533), .IN2(n6512), .QN(n6692) );
  NAND4X0 U8523 ( .IN1(n6513), .IN2(n8860), .IN3(n7612), .IN4(n6692), .QN(
        n6514) );
  NOR4X0 U8524 ( .IN1(n8638), .IN2(n6791), .IN3(n6515), .IN4(n6514), .QN(n6518) );
  NAND2X0 U8525 ( .IN1(n9082), .IN2(n6516), .QN(n8366) );
  NAND4X0 U8526 ( .IN1(n6519), .IN2(n6518), .IN3(n6517), .IN4(n8366), .QN(
        \a4/N462 ) );
  NOR2X0 U8527 ( .IN1(n9084), .IN2(n8515), .QN(n9134) );
  NOR2X0 U8528 ( .IN1(n9134), .IN2(n8518), .QN(n7106) );
  OA21X1 U8529 ( .IN1(n9438), .IN2(n6520), .IN3(n6662), .Q(n6530) );
  AND3X1 U8530 ( .IN1(n7437), .IN2(n8640), .IN3(n8282), .Q(n6527) );
  NAND2X0 U8531 ( .IN1(degrees_tmp2[2]), .IN2(n6521), .QN(n6522) );
  NAND3X0 U8532 ( .IN1(n6522), .IN2(n7307), .IN3(n6996), .QN(n6526) );
  INVX0 U8533 ( .INP(n6523), .ZN(n7166) );
  NAND4X0 U8534 ( .IN1(n8421), .IN2(n7166), .IN3(n6524), .IN4(n7968), .QN(
        n6525) );
  NOR4X0 U8535 ( .IN1(n7269), .IN2(n6527), .IN3(n6526), .IN4(n6525), .QN(n6529) );
  INVX0 U8536 ( .INP(n6528), .ZN(n7818) );
  NAND4X0 U8537 ( .IN1(n7106), .IN2(n6530), .IN3(n6529), .IN4(n7818), .QN(
        \a4/N463 ) );
  NAND3X0 U8538 ( .IN1(n9210), .IN2(degrees_tmp2[0]), .IN3(n9099), .QN(n6531)
         );
  NAND4X0 U8539 ( .IN1(n8979), .IN2(n7510), .IN3(n8316), .IN4(n6531), .QN(
        n6533) );
  AO22X1 U8540 ( .IN1(n9073), .IN2(n6533), .IN3(n6532), .IN4(n9099), .Q(n6540)
         );
  OA21X1 U8541 ( .IN1(n7517), .IN2(n8406), .IN3(n6534), .Q(n6538) );
  OA22X1 U8542 ( .IN1(n9122), .IN2(n7685), .IN3(n8431), .IN4(n6951), .Q(n6537)
         );
  NAND4X0 U8543 ( .IN1(n6538), .IN2(n6537), .IN3(n6536), .IN4(n6535), .QN(
        n6539) );
  NOR4X0 U8544 ( .IN1(n6541), .IN2(n6745), .IN3(n6540), .IN4(n6539), .QN(n6542) );
  NAND4X0 U8545 ( .IN1(n6542), .IN2(n7577), .IN3(n7156), .IN4(n6696), .QN(
        \a4/N464 ) );
  INVX0 U8546 ( .INP(n8664), .ZN(n6550) );
  OR2X1 U8547 ( .IN1(n9440), .IN2(n8705), .Q(n8609) );
  NAND2X0 U8548 ( .IN1(n9169), .IN2(n8609), .QN(n7477) );
  NOR2X0 U8549 ( .IN1(n6623), .IN2(n6543), .QN(n6544) );
  OA22X1 U8550 ( .IN1(n7841), .IN2(n8281), .IN3(n6544), .IN4(n7945), .Q(n6548)
         );
  OA22X1 U8551 ( .IN1(n9031), .IN2(n8303), .IN3(n8204), .IN4(n8782), .Q(n6547)
         );
  NAND2X0 U8552 ( .IN1(n6545), .IN2(n9032), .QN(n6546) );
  NAND4X0 U8553 ( .IN1(n6548), .IN2(n6547), .IN3(n8820), .IN4(n6546), .QN(
        n6549) );
  NOR4X0 U8554 ( .IN1(n6550), .IN2(n7338), .IN3(n7477), .IN4(n6549), .QN(n6552) );
  NAND2X0 U8555 ( .IN1(n6929), .IN2(n8041), .QN(n6551) );
  NAND4X0 U8556 ( .IN1(n6552), .IN2(n6551), .IN3(n6915), .IN4(n8410), .QN(
        \a4/N465 ) );
  NOR2X0 U8557 ( .IN1(n8533), .IN2(n8262), .QN(n7946) );
  NOR2X0 U8558 ( .IN1(n6554), .IN2(n6553), .QN(n7320) );
  NOR4X0 U8559 ( .IN1(n7934), .IN2(n8985), .IN3(n7946), .IN4(n7320), .QN(n6564) );
  OA22X1 U8560 ( .IN1(n8825), .IN2(n7633), .IN3(n9436), .IN4(n8612), .Q(n6563)
         );
  NAND2X0 U8561 ( .IN1(n9112), .IN2(n6555), .QN(n6560) );
  NAND2X0 U8562 ( .IN1(n8575), .IN2(n6556), .QN(n6558) );
  NAND2X0 U8563 ( .IN1(degrees_tmp2[5]), .IN2(n7693), .QN(n7241) );
  NAND3X0 U8564 ( .IN1(n6558), .IN2(n7241), .IN3(n6557), .QN(n6559) );
  NOR4X0 U8565 ( .IN1(n8077), .IN2(n6561), .IN3(n6560), .IN4(n6559), .QN(n6562) );
  NAND2X0 U8566 ( .IN1(n9156), .IN2(n7745), .QN(n6803) );
  NAND4X0 U8567 ( .IN1(n6564), .IN2(n6563), .IN3(n6562), .IN4(n6803), .QN(
        \a4/N466 ) );
  INVX0 U8568 ( .INP(n8584), .ZN(n8078) );
  NOR2X0 U8569 ( .IN1(n9171), .IN2(n8105), .QN(n6566) );
  NAND2X0 U8570 ( .IN1(n8724), .IN2(n7033), .QN(n6565) );
  NAND2X0 U8571 ( .IN1(n6566), .IN2(n6565), .QN(n6573) );
  OA22X1 U8572 ( .IN1(n7084), .IN2(n8303), .IN3(n8573), .IN4(n8067), .Q(n6571)
         );
  NAND2X0 U8573 ( .IN1(n6568), .IN2(n6567), .QN(n7134) );
  NAND2X0 U8574 ( .IN1(n8533), .IN2(n7134), .QN(n6636) );
  NAND2X0 U8575 ( .IN1(n9023), .IN2(n6569), .QN(n6570) );
  NAND4X0 U8576 ( .IN1(n6571), .IN2(n7022), .IN3(n6636), .IN4(n6570), .QN(
        n6572) );
  NOR4X0 U8577 ( .IN1(n8078), .IN2(n7483), .IN3(n6573), .IN4(n6572), .QN(n6577) );
  NOR2X0 U8578 ( .IN1(n6575), .IN2(n6574), .QN(n8344) );
  NAND2X0 U8579 ( .IN1(n8344), .IN2(n9442), .QN(n6576) );
  NAND4X0 U8580 ( .IN1(n6577), .IN2(n8364), .IN3(n6996), .IN4(n6576), .QN(
        \a4/N467 ) );
  NAND2X0 U8581 ( .IN1(n6859), .IN2(n8533), .QN(n9057) );
  NAND2X0 U8582 ( .IN1(n8730), .IN2(n7214), .QN(n8695) );
  NAND4X0 U8583 ( .IN1(n8928), .IN2(n6588), .IN3(n9057), .IN4(n8695), .QN(
        n6583) );
  INVX0 U8584 ( .INP(n7849), .ZN(n9101) );
  NAND2X0 U8585 ( .IN1(n7484), .IN2(n9048), .QN(n6869) );
  NAND4X0 U8586 ( .IN1(n8817), .IN2(n8720), .IN3(n9101), .IN4(n6869), .QN(
        n6582) );
  OR2X1 U8587 ( .IN1(n7736), .IN2(n6832), .Q(n8775) );
  NAND2X0 U8588 ( .IN1(n8775), .IN2(n6578), .QN(n6871) );
  INVX0 U8589 ( .INP(n6871), .ZN(n6580) );
  NAND2X0 U8590 ( .IN1(n7945), .IN2(n8282), .QN(n8086) );
  NAND3X0 U8591 ( .IN1(n8186), .IN2(degrees_tmp2[2]), .IN3(n8086), .QN(n6579)
         );
  NAND3X0 U8592 ( .IN1(n6580), .IN2(n8135), .IN3(n6579), .QN(n6581) );
  NOR4X0 U8593 ( .IN1(n7964), .IN2(n6583), .IN3(n6582), .IN4(n6581), .QN(n6586) );
  INVX0 U8594 ( .INP(n6584), .ZN(n6585) );
  NAND2X0 U8595 ( .IN1(n8519), .IN2(n9183), .QN(n8441) );
  NAND4X0 U8596 ( .IN1(n6586), .IN2(n6585), .IN3(n7302), .IN4(n8441), .QN(
        \a4/N468 ) );
  INVX0 U8597 ( .INP(n6587), .ZN(n6592) );
  NAND3X0 U8598 ( .IN1(n6588), .IN2(n8317), .IN3(n7404), .QN(n6589) );
  NAND2X0 U8599 ( .IN1(n6589), .IN2(n8825), .QN(n6590) );
  NAND4X0 U8600 ( .IN1(n6592), .IN2(n8817), .IN3(n6591), .IN4(n6590), .QN(
        n6593) );
  NOR4X0 U8601 ( .IN1(n7520), .IN2(n8358), .IN3(n6594), .IN4(n6593), .QN(n6596) );
  NAND2X0 U8602 ( .IN1(n8640), .IN2(n7945), .QN(n6595) );
  NAND4X0 U8603 ( .IN1(n6597), .IN2(n6596), .IN3(n6595), .IN4(n6696), .QN(
        \a4/N469 ) );
  NOR2X0 U8604 ( .IN1(n6797), .IN2(n8685), .QN(n6598) );
  NOR4X0 U8605 ( .IN1(n6599), .IN2(n8660), .IN3(n8369), .IN4(n6598), .QN(n6610) );
  NAND4X0 U8606 ( .IN1(n8384), .IN2(n8820), .IN3(n8412), .IN4(n8068), .QN(
        n6604) );
  AO22X1 U8607 ( .IN1(n7236), .IN2(n8086), .IN3(n8496), .IN4(n7808), .Q(n6602)
         );
  NOR2X0 U8608 ( .IN1(n9445), .IN2(n6600), .QN(n8755) );
  AO22X1 U8609 ( .IN1(n8755), .IN2(n8692), .IN3(n6782), .IN4(n8780), .Q(n6601)
         );
  NOR4X0 U8610 ( .IN1(n6604), .IN2(n6603), .IN3(n6602), .IN4(n6601), .QN(n6609) );
  NAND3X0 U8611 ( .IN1(n6606), .IN2(n6605), .IN3(n8401), .QN(n6607) );
  NAND2X0 U8612 ( .IN1(n6607), .IN2(n8816), .QN(n6608) );
  NAND2X0 U8613 ( .IN1(n8699), .IN2(n7669), .QN(n8189) );
  NAND4X0 U8614 ( .IN1(n6610), .IN2(n6609), .IN3(n6608), .IN4(n8189), .QN(
        \a4/N471 ) );
  INVX0 U8615 ( .INP(n6611), .ZN(n8103) );
  NAND2X0 U8616 ( .IN1(n9131), .IN2(n7784), .QN(n8385) );
  OA22X1 U8617 ( .IN1(n8103), .IN2(n6612), .IN3(n8268), .IN4(n8385), .Q(n6622)
         );
  NAND4X0 U8618 ( .IN1(n7340), .IN2(n7965), .IN3(n7131), .IN4(n7583), .QN(
        n6618) );
  NAND2X0 U8619 ( .IN1(n8978), .IN2(n6613), .QN(n8264) );
  INVX0 U8620 ( .INP(n7581), .ZN(n8508) );
  OA22X1 U8621 ( .IN1(n6614), .IN2(n8264), .IN3(n8752), .IN4(n8508), .Q(n6616)
         );
  AO221X1 U8622 ( .IN1(n7463), .IN2(n6747), .IN3(n7463), .IN4(n8938), .IN5(
        n8724), .Q(n6615) );
  NAND4X0 U8623 ( .IN1(n6616), .IN2(n6892), .IN3(n8514), .IN4(n6615), .QN(
        n6617) );
  NOR2X0 U8624 ( .IN1(n6618), .IN2(n6617), .QN(n6621) );
  NAND2X0 U8625 ( .IN1(n6620), .IN2(n6619), .QN(n7240) );
  NAND4X0 U8626 ( .IN1(n6622), .IN2(n6621), .IN3(n7789), .IN4(n7240), .QN(
        \a4/N472 ) );
  NAND2X0 U8627 ( .IN1(n6623), .IN2(n7233), .QN(n8228) );
  NAND2X0 U8628 ( .IN1(n8445), .IN2(n8228), .QN(n6625) );
  NOR2X0 U8629 ( .IN1(n6624), .IN2(n7745), .QN(n6824) );
  AO22X1 U8630 ( .IN1(n8675), .IN2(n6625), .IN3(n6824), .IN4(n8034), .Q(n6632)
         );
  NOR2X0 U8631 ( .IN1(n7577), .IN2(n8598), .QN(n6627) );
  NAND2X0 U8632 ( .IN1(n7700), .IN2(n9033), .QN(n8263) );
  NAND2X0 U8633 ( .IN1(n8263), .IN2(n8927), .QN(n6626) );
  NOR2X0 U8634 ( .IN1(n6627), .IN2(n6626), .QN(n6630) );
  OA22X1 U8635 ( .IN1(n9442), .IN2(n8846), .IN3(n7463), .IN4(n7897), .Q(n6629)
         );
  NAND2X0 U8636 ( .IN1(n9123), .IN2(n9155), .QN(n6785) );
  NAND4X0 U8637 ( .IN1(n6630), .IN2(n6629), .IN3(n6628), .IN4(n6785), .QN(
        n6631) );
  NOR2X0 U8638 ( .IN1(n6632), .IN2(n6631), .QN(n6633) );
  NAND4X0 U8639 ( .IN1(n6633), .IN2(n8380), .IN3(n7738), .IN4(n7721), .QN(
        \a4/N473 ) );
  NOR2X0 U8640 ( .IN1(n6635), .IN2(n6634), .QN(n6645) );
  NOR2X0 U8641 ( .IN1(n7425), .IN2(n7908), .QN(n7605) );
  OA21X1 U8642 ( .IN1(n9441), .IN2(n6636), .IN3(n7605), .Q(n6643) );
  OA22X1 U8643 ( .IN1(n8728), .IN2(n9165), .IN3(n7668), .IN4(n8349), .Q(n6642)
         );
  NOR2X0 U8644 ( .IN1(n6638), .IN2(n6637), .QN(n6639) );
  OA22X1 U8645 ( .IN1(n8760), .IN2(n8968), .IN3(n6639), .IN4(n8782), .Q(n6641)
         );
  NAND2X0 U8646 ( .IN1(n9437), .IN2(n6640), .QN(n7797) );
  NAND4X0 U8647 ( .IN1(n6643), .IN2(n6642), .IN3(n6641), .IN4(n7797), .QN(
        n6644) );
  OR4X1 U8648 ( .IN1(n6647), .IN2(n6646), .IN3(n6645), .IN4(n6644), .Q(
        \a4/N474 ) );
  INVX0 U8649 ( .INP(n6648), .ZN(n8540) );
  OA22X1 U8650 ( .IN1(n6649), .IN2(n8540), .IN3(n8804), .IN4(n9436), .Q(n6664)
         );
  OA21X1 U8651 ( .IN1(n6668), .IN2(n7934), .IN3(n8588), .Q(n6659) );
  NOR2X0 U8652 ( .IN1(n9437), .IN2(n8461), .QN(n7707) );
  AO22X1 U8653 ( .IN1(n9182), .IN2(n6736), .IN3(n6697), .IN4(n7707), .Q(n6658)
         );
  OA21X1 U8654 ( .IN1(n6650), .IN2(n8996), .IN3(n8966), .Q(n6656) );
  NOR2X0 U8655 ( .IN1(n6651), .IN2(n8588), .QN(n6653) );
  NAND2X0 U8656 ( .IN1(n8846), .IN2(n8904), .QN(n6652) );
  NAND2X0 U8657 ( .IN1(n6653), .IN2(n6652), .QN(n6654) );
  NAND4X0 U8658 ( .IN1(n6656), .IN2(n6655), .IN3(n7307), .IN4(n6654), .QN(
        n6657) );
  NOR3X0 U8659 ( .IN1(n6659), .IN2(n6658), .IN3(n6657), .QN(n6663) );
  NAND2X0 U8660 ( .IN1(n6661), .IN2(n6660), .QN(n9055) );
  NAND4X0 U8661 ( .IN1(n6664), .IN2(n6663), .IN3(n6662), .IN4(n9055), .QN(
        \a4/N475 ) );
  NOR2X0 U8662 ( .IN1(n7077), .IN2(n8855), .QN(n6676) );
  OA21X1 U8663 ( .IN1(n8753), .IN2(n6665), .IN3(n8730), .Q(n6666) );
  NOR4X0 U8664 ( .IN1(n8994), .IN2(n6667), .IN3(n6974), .IN4(n6666), .QN(n6675) );
  AO22X1 U8665 ( .IN1(n8696), .IN2(n8239), .IN3(n6668), .IN4(n8649), .Q(n6671)
         );
  NAND4X0 U8666 ( .IN1(n8338), .IN2(n6669), .IN3(n8056), .IN4(n7633), .QN(
        n6670) );
  NOR4X0 U8667 ( .IN1(n8458), .IN2(n6672), .IN3(n6671), .IN4(n6670), .QN(n6674) );
  NAND2X0 U8668 ( .IN1(n8566), .IN2(n6836), .QN(n6673) );
  NAND4X0 U8669 ( .IN1(n6676), .IN2(n6675), .IN3(n6674), .IN4(n6673), .QN(
        \a4/N477 ) );
  NOR2X0 U8670 ( .IN1(n8022), .IN2(n8411), .QN(n8658) );
  NAND2X0 U8671 ( .IN1(n8432), .IN2(n8171), .QN(n7855) );
  NAND4X0 U8672 ( .IN1(n7111), .IN2(n7362), .IN3(n8029), .IN4(n7855), .QN(
        n6683) );
  NAND4X0 U8673 ( .IN1(n8106), .IN2(n8399), .IN3(n6677), .IN4(n8504), .QN(
        n6682) );
  NAND3X0 U8674 ( .IN1(n9442), .IN2(n6678), .IN3(n7208), .QN(n6680) );
  NAND2X0 U8675 ( .IN1(n6680), .IN2(n6679), .QN(n6681) );
  NOR4X0 U8676 ( .IN1(n8658), .IN2(n6683), .IN3(n6682), .IN4(n6681), .QN(n6685) );
  NAND4X0 U8677 ( .IN1(n6685), .IN2(n7764), .IN3(n6701), .IN4(n6684), .QN(
        \a4/N478 ) );
  AND2X1 U8678 ( .IN1(n9140), .IN2(n8230), .Q(n6695) );
  NOR4X0 U8679 ( .IN1(n8359), .IN2(n9009), .IN3(n7754), .IN4(n6719), .QN(n6694) );
  OA21X1 U8680 ( .IN1(n7436), .IN2(n6686), .IN3(n8598), .Q(n6691) );
  NOR2X0 U8681 ( .IN1(n9435), .IN2(n6687), .QN(n8016) );
  OA21X1 U8682 ( .IN1(n8475), .IN2(n6688), .IN3(n9440), .Q(n6690) );
  NAND2X0 U8683 ( .IN1(n6689), .IN2(n6937), .QN(n7492) );
  NOR4X0 U8684 ( .IN1(n6691), .IN2(n8016), .IN3(n6690), .IN4(n7492), .QN(n6693) );
  NAND4X0 U8685 ( .IN1(n6695), .IN2(n6694), .IN3(n6693), .IN4(n6692), .QN(
        \a4/N479 ) );
  INVX0 U8686 ( .INP(n7647), .ZN(n8371) );
  NAND2X0 U8687 ( .IN1(n9037), .IN2(n8371), .QN(n7568) );
  NAND4X0 U8688 ( .IN1(n7729), .IN2(n6696), .IN3(n8411), .IN4(n7568), .QN(
        n6704) );
  INVX0 U8689 ( .INP(n6697), .ZN(n7933) );
  OA22X1 U8690 ( .IN1(n8461), .IN2(n7933), .IN3(n7234), .IN4(n7571), .Q(n6702)
         );
  NAND2X0 U8691 ( .IN1(n6699), .IN2(n6698), .QN(n6700) );
  NAND4X0 U8692 ( .IN1(n6702), .IN2(n6701), .IN3(n7865), .IN4(n6700), .QN(
        n6703) );
  NOR2X0 U8693 ( .IN1(n6704), .IN2(n6703), .QN(n6707) );
  AO21X1 U8694 ( .IN1(n8564), .IN2(n9083), .IN3(n8787), .Q(n6705) );
  NAND4X0 U8695 ( .IN1(n6707), .IN2(n9111), .IN3(n6706), .IN4(n6705), .QN(
        \a4/N480 ) );
  OA22X1 U8696 ( .IN1(n7656), .IN2(n7316), .IN3(n8752), .IN4(n8845), .Q(n6718)
         );
  AO22X1 U8697 ( .IN1(n8242), .IN2(n6709), .IN3(n6708), .IN4(n9442), .Q(n6716)
         );
  NAND2X0 U8698 ( .IN1(n8180), .IN2(n8727), .QN(n7097) );
  OAI22X1 U8699 ( .IN1(n8910), .IN2(n6710), .IN3(n7097), .IN4(degrees_tmp2[3]), 
        .QN(n6715) );
  NAND2X0 U8700 ( .IN1(n9035), .IN2(n8947), .QN(n6963) );
  NOR2X0 U8701 ( .IN1(n8816), .IN2(n7548), .QN(n6711) );
  NAND2X0 U8702 ( .IN1(n6711), .IN2(n9445), .QN(n6713) );
  NAND3X0 U8703 ( .IN1(n7999), .IN2(n9209), .IN3(n8034), .QN(n6712) );
  NAND4X0 U8704 ( .IN1(n8846), .IN2(n6963), .IN3(n6713), .IN4(n6712), .QN(
        n6714) );
  NOR4X0 U8705 ( .IN1(n8786), .IN2(n6716), .IN3(n6715), .IN4(n6714), .QN(n6717) );
  NAND4X0 U8706 ( .IN1(n6718), .IN2(n6717), .IN3(n7245), .IN4(n7494), .QN(
        \a4/N481 ) );
  OA21X1 U8707 ( .IN1(degrees_tmp2[3]), .IN2(n8801), .IN3(n6996), .Q(n6725) );
  INVX0 U8708 ( .INP(n8846), .ZN(n7952) );
  NOR2X0 U8709 ( .IN1(n7952), .IN2(n6719), .QN(n8916) );
  NOR4X0 U8710 ( .IN1(n7333), .IN2(n9014), .IN3(n9039), .IN4(n6720), .QN(n6721) );
  AND4X1 U8711 ( .IN1(n8916), .IN2(n6721), .IN3(n8893), .IN4(n8964), .Q(n6724)
         );
  NAND2X0 U8712 ( .IN1(n9125), .IN2(n7703), .QN(n6722) );
  NAND4X0 U8713 ( .IN1(n6725), .IN2(n6724), .IN3(n6723), .IN4(n6722), .QN(
        \a4/N482 ) );
  OA22X1 U8714 ( .IN1(n8461), .IN2(n8303), .IN3(n9031), .IN4(n8264), .Q(n6735)
         );
  INVX0 U8715 ( .INP(n6726), .ZN(n8473) );
  NOR2X0 U8716 ( .IN1(n8752), .IN2(n6727), .QN(n6733) );
  INVX0 U8717 ( .INP(n8788), .ZN(n8914) );
  OA22X1 U8718 ( .IN1(n8675), .IN2(n6728), .IN3(n7169), .IN4(n8914), .Q(n6731)
         );
  NAND3X0 U8719 ( .IN1(n7806), .IN2(n7736), .IN3(n7686), .QN(n6729) );
  NAND4X0 U8720 ( .IN1(n6731), .IN2(n6730), .IN3(n8125), .IN4(n6729), .QN(
        n6732) );
  NOR4X0 U8721 ( .IN1(n8473), .IN2(n8982), .IN3(n6733), .IN4(n6732), .QN(n6734) );
  NAND4X0 U8722 ( .IN1(n6735), .IN2(n6734), .IN3(n7587), .IN4(n7165), .QN(
        \a4/N483 ) );
  NOR2X0 U8723 ( .IN1(n8268), .IN2(n6804), .QN(n6743) );
  INVX0 U8724 ( .INP(n6736), .ZN(n8168) );
  OA22X1 U8725 ( .IN1(n9131), .IN2(n8491), .IN3(n8168), .IN4(n8204), .Q(n6741)
         );
  INVX0 U8726 ( .INP(n6737), .ZN(n6740) );
  NAND3X0 U8727 ( .IN1(n8816), .IN2(n9105), .IN3(n8909), .QN(n6738) );
  NAND4X0 U8728 ( .IN1(n6741), .IN2(n6740), .IN3(n6739), .IN4(n6738), .QN(
        n6742) );
  NOR4X0 U8729 ( .IN1(n6745), .IN2(n6744), .IN3(n6743), .IN4(n6742), .QN(n6746) );
  INVX0 U8730 ( .INP(n7608), .ZN(n8774) );
  NAND2X0 U8731 ( .IN1(n8774), .IN2(n9445), .QN(n8374) );
  NAND3X0 U8732 ( .IN1(n6746), .IN2(n6945), .IN3(n8374), .QN(\a4/N484 ) );
  OR2X1 U8733 ( .IN1(n6747), .IN2(n8938), .Q(n6748) );
  OA22X1 U8734 ( .IN1(n8883), .IN2(n8349), .IN3(degrees_tmp2[3]), .IN4(n6748), 
        .Q(n6754) );
  INVX0 U8735 ( .INP(n7499), .ZN(n6750) );
  NAND2X0 U8736 ( .IN1(n7517), .IN2(n8529), .QN(n8732) );
  NAND3X0 U8737 ( .IN1(n8555), .IN2(n7334), .IN3(n8732), .QN(n6749) );
  NOR4X0 U8738 ( .IN1(n6751), .IN2(n6750), .IN3(n8472), .IN4(n6749), .QN(n6753) );
  NAND2X0 U8739 ( .IN1(n7179), .IN2(n7236), .QN(n6752) );
  NAND4X0 U8740 ( .IN1(n6754), .IN2(n6753), .IN3(n7498), .IN4(n6752), .QN(
        \a4/N486 ) );
  AOI22X1 U8741 ( .IN1(n8468), .IN2(n9026), .IN3(n6756), .IN4(n6755), .QN(
        n6757) );
  INVX0 U8742 ( .INP(n7759), .ZN(n8759) );
  NAND4X0 U8743 ( .IN1(n6757), .IN2(n7499), .IN3(n8294), .IN4(n8759), .QN(
        \a4/N487 ) );
  NAND2X0 U8744 ( .IN1(n6758), .IN2(n9166), .QN(n6760) );
  NAND3X0 U8745 ( .IN1(n6761), .IN2(n6760), .IN3(n6759), .QN(\a4/N488 ) );
  AND2X1 U8746 ( .IN1(n8220), .IN2(n6762), .Q(\a4/N492 ) );
  NAND2X0 U8747 ( .IN1(n8861), .IN2(n8731), .QN(n6764) );
  NAND3X0 U8748 ( .IN1(n6764), .IN2(n6763), .IN3(n8522), .QN(n6770) );
  AO21X1 U8749 ( .IN1(n8684), .IN2(n7596), .IN3(n8282), .Q(n6765) );
  NAND3X0 U8750 ( .IN1(n9212), .IN2(n7881), .IN3(n6765), .QN(n6769) );
  NAND2X0 U8751 ( .IN1(n6766), .IN2(n8467), .QN(n7187) );
  NAND4X0 U8752 ( .IN1(n8347), .IN2(n6786), .IN3(n6767), .IN4(n7187), .QN(
        n6768) );
  NOR4X0 U8753 ( .IN1(n7203), .IN2(n6770), .IN3(n6769), .IN4(n6768), .QN(n6772) );
  NAND2X0 U8754 ( .IN1(degrees_tmp2[0]), .IN2(n8459), .QN(n7091) );
  INVX0 U8755 ( .INP(n6771), .ZN(n8541) );
  NAND4X0 U8756 ( .IN1(n6772), .IN2(n7730), .IN3(n7091), .IN4(n8541), .QN(
        \a3/N436 ) );
  OA221X1 U8757 ( .IN1(degrees_tmp2[0]), .IN2(n6773), .IN3(degrees_tmp2[0]), 
        .IN4(n8967), .IN5(n8615), .Q(n6779) );
  INVX0 U8758 ( .INP(n8263), .ZN(n8111) );
  NAND2X0 U8759 ( .IN1(n8545), .IN2(n6908), .QN(n8033) );
  AO221X1 U8760 ( .IN1(n9125), .IN2(n7645), .IN3(n9125), .IN4(n8033), .IN5(
        n8048), .Q(n6777) );
  OA22X1 U8761 ( .IN1(n8185), .IN2(n8507), .IN3(n8752), .IN4(n8859), .Q(n6775)
         );
  NOR2X0 U8762 ( .IN1(n7168), .IN2(n7686), .QN(n7894) );
  NAND2X0 U8763 ( .IN1(n7894), .IN2(n8692), .QN(n6774) );
  NAND2X0 U8764 ( .IN1(n9190), .IN2(n9209), .QN(n8850) );
  NAND4X0 U8765 ( .IN1(n6775), .IN2(n8885), .IN3(n6774), .IN4(n8850), .QN(
        n6776) );
  NOR4X0 U8766 ( .IN1(n9024), .IN2(n8111), .IN3(n6777), .IN4(n6776), .QN(n6778) );
  NAND4X0 U8767 ( .IN1(n6779), .IN2(n6778), .IN3(n8231), .IN4(n7818), .QN(
        \a3/N437 ) );
  AOI22X1 U8768 ( .IN1(n8724), .IN2(n8320), .IN3(n8675), .IN4(n7198), .QN(
        n6793) );
  NAND2X0 U8769 ( .IN1(n8020), .IN2(n8571), .QN(n6789) );
  AND3X1 U8770 ( .IN1(n6780), .IN2(n9436), .IN3(n7808), .Q(n6784) );
  AO22X1 U8771 ( .IN1(n6782), .IN2(n8630), .IN3(n8511), .IN4(n6781), .Q(n6783)
         );
  NOR4X0 U8772 ( .IN1(n7611), .IN2(n6784), .IN3(n8923), .IN4(n6783), .QN(n6787) );
  NAND4X0 U8773 ( .IN1(n6787), .IN2(n8292), .IN3(n6786), .IN4(n6785), .QN(
        n6788) );
  NOR4X0 U8774 ( .IN1(n6791), .IN2(n6790), .IN3(n6789), .IN4(n6788), .QN(n6792) );
  INVX0 U8775 ( .INP(n9098), .ZN(n8352) );
  NAND2X0 U8776 ( .IN1(n7517), .IN2(n8352), .QN(n7113) );
  NAND2X0 U8777 ( .IN1(n9074), .IN2(n8041), .QN(n7299) );
  NAND4X0 U8778 ( .IN1(n6793), .IN2(n6792), .IN3(n7113), .IN4(n7299), .QN(
        \a3/N438 ) );
  AND2X1 U8779 ( .IN1(n8922), .IN2(n6794), .Q(n6795) );
  OA22X1 U8780 ( .IN1(n8978), .IN2(n8406), .IN3(n6795), .IN4(n9122), .Q(n6810)
         );
  NOR2X0 U8781 ( .IN1(n8408), .IN2(n6980), .QN(n6796) );
  OA22X1 U8782 ( .IN1(n9183), .IN2(n6965), .IN3(n6796), .IN4(n9155), .Q(n6809)
         );
  AOI22X1 U8783 ( .IN1(n6797), .IN2(n9005), .IN3(n7645), .IN4(n9023), .QN(
        n6801) );
  NAND3X0 U8784 ( .IN1(n8022), .IN2(n6934), .IN3(n8595), .QN(n6798) );
  AND4X1 U8785 ( .IN1(n6801), .IN2(n6800), .IN3(n6799), .IN4(n6798), .Q(n6802)
         );
  OA21X1 U8786 ( .IN1(n9438), .IN2(n6803), .IN3(n6802), .Q(n6808) );
  NAND2X0 U8787 ( .IN1(n9045), .IN2(n6804), .QN(n6806) );
  NAND3X0 U8788 ( .IN1(n6806), .IN2(n8568), .IN3(n6805), .QN(n6807) );
  NAND4X0 U8789 ( .IN1(n6810), .IN2(n6809), .IN3(n6808), .IN4(n6807), .QN(
        \a3/N439 ) );
  OA22X1 U8790 ( .IN1(n6936), .IN2(n8979), .IN3(n9433), .IN4(n6811), .Q(n6815)
         );
  NAND4X0 U8791 ( .IN1(n8914), .IN2(n8574), .IN3(n8868), .IN4(n7183), .QN(
        n6812) );
  NAND2X0 U8792 ( .IN1(n8004), .IN2(n6812), .QN(n6813) );
  AND4X1 U8793 ( .IN1(n6815), .IN2(n8156), .IN3(n6814), .IN4(n6813), .Q(n6817)
         );
  NAND2X0 U8794 ( .IN1(n7523), .IN2(n7945), .QN(n6816) );
  NAND2X0 U8795 ( .IN1(n8519), .IN2(n8649), .QN(n7381) );
  NAND4X0 U8796 ( .IN1(n6818), .IN2(n6817), .IN3(n6816), .IN4(n7381), .QN(
        \a3/N441 ) );
  NOR2X0 U8797 ( .IN1(n6819), .IN2(n9082), .QN(n6822) );
  AO21X1 U8798 ( .IN1(n8678), .IN2(n8596), .IN3(n8185), .Q(n6820) );
  NAND2X0 U8799 ( .IN1(n7437), .IN2(n7894), .QN(n7829) );
  NAND2X0 U8800 ( .IN1(n6820), .IN2(n7829), .QN(n6821) );
  NOR2X0 U8801 ( .IN1(n6822), .IN2(n6821), .QN(n6831) );
  OA221X1 U8802 ( .IN1(n9048), .IN2(n6823), .IN3(n9048), .IN4(n8801), .IN5(
        n7459), .Q(n6830) );
  NOR4X0 U8803 ( .IN1(n8058), .IN2(n7281), .IN3(n7342), .IN4(n6824), .QN(n6825) );
  NOR2X0 U8804 ( .IN1(n6825), .IN2(n6836), .QN(n6828) );
  AND3X1 U8805 ( .IN1(n8572), .IN2(n6826), .IN3(n7842), .Q(n7719) );
  OA21X1 U8806 ( .IN1(n9075), .IN2(n7133), .IN3(n8598), .Q(n6827) );
  NOR4X0 U8807 ( .IN1(n6828), .IN2(n9066), .IN3(n7719), .IN4(n6827), .QN(n6829) );
  NAND4X0 U8808 ( .IN1(n6831), .IN2(n6830), .IN3(n6829), .IN4(n8892), .QN(
        \a3/N442 ) );
  OA22X1 U8809 ( .IN1(n9433), .IN2(n8668), .IN3(n6833), .IN4(n6832), .Q(n8238)
         );
  INVX0 U8810 ( .INP(n6834), .ZN(n6843) );
  INVX0 U8811 ( .INP(n8660), .ZN(n6841) );
  NAND3X0 U8812 ( .IN1(n7538), .IN2(n8039), .IN3(n6835), .QN(n6837) );
  NAND2X0 U8813 ( .IN1(n6837), .IN2(n6836), .QN(n6839) );
  NOR2X0 U8814 ( .IN1(n8567), .IN2(n7936), .QN(n7572) );
  AO221X1 U8815 ( .IN1(n8937), .IN2(n7572), .IN3(n8937), .IN4(n9440), .IN5(
        n9122), .Q(n6838) );
  NAND4X0 U8816 ( .IN1(n6841), .IN2(n6840), .IN3(n6839), .IN4(n6838), .QN(
        n6842) );
  NOR4X0 U8817 ( .IN1(n7850), .IN2(n8953), .IN3(n6843), .IN4(n6842), .QN(n6846) );
  NAND2X0 U8818 ( .IN1(n8727), .IN2(n8320), .QN(n6844) );
  NAND4X0 U8819 ( .IN1(n8238), .IN2(n6846), .IN3(n6845), .IN4(n6844), .QN(
        \a3/N443 ) );
  OA21X1 U8820 ( .IN1(n6893), .IN2(n8385), .IN3(n6847), .Q(n6848) );
  AND4X1 U8821 ( .IN1(n6848), .IN2(n8669), .IN3(n8803), .IN4(n7820), .Q(n6858)
         );
  NOR2X0 U8822 ( .IN1(n9436), .IN2(n7990), .QN(n8343) );
  NAND4X0 U8823 ( .IN1(n8193), .IN2(n7872), .IN3(n8613), .IN4(n6849), .QN(
        n6855) );
  NOR2X0 U8824 ( .IN1(n6851), .IN2(n6850), .QN(n6853) );
  NAND2X0 U8825 ( .IN1(n8924), .IN2(n9445), .QN(n6852) );
  NAND2X0 U8826 ( .IN1(n6853), .IN2(n6852), .QN(n6854) );
  NOR4X0 U8827 ( .IN1(n6856), .IN2(n8343), .IN3(n6855), .IN4(n6854), .QN(n6857) );
  NAND4X0 U8828 ( .IN1(n6858), .IN2(n6857), .IN3(n7480), .IN4(n8532), .QN(
        \a3/N444 ) );
  AO221X1 U8829 ( .IN1(n6859), .IN2(n8467), .IN3(n6859), .IN4(n7935), .IN5(
        n8855), .Q(n6860) );
  NOR4X0 U8830 ( .IN1(n7192), .IN2(n6862), .IN3(n6861), .IN4(n6860), .QN(n6868) );
  NAND2X0 U8831 ( .IN1(n7018), .IN2(n7245), .QN(n6918) );
  AO22X1 U8832 ( .IN1(n8468), .IN2(n6863), .IN3(n7700), .IN4(n7699), .Q(n6864)
         );
  NOR4X0 U8833 ( .IN1(n6865), .IN2(n7775), .IN3(n6918), .IN4(n6864), .QN(n6867) );
  NAND2X0 U8834 ( .IN1(n7916), .IN2(n8494), .QN(n6866) );
  NAND4X0 U8835 ( .IN1(n6868), .IN2(n6867), .IN3(n7747), .IN4(n6866), .QN(
        \a3/N445 ) );
  OA22X1 U8836 ( .IN1(n8727), .IN2(n6951), .IN3(n9442), .IN4(n6869), .Q(n6876)
         );
  OA22X1 U8837 ( .IN1(n9031), .IN2(n7638), .IN3(n8909), .IN4(n9126), .Q(n6875)
         );
  NAND2X0 U8838 ( .IN1(n8432), .IN2(n9071), .QN(n8038) );
  NAND4X0 U8839 ( .IN1(n8279), .IN2(n7533), .IN3(n7585), .IN4(n8038), .QN(
        n6870) );
  NOR4X0 U8840 ( .IN1(n7652), .IN2(n7581), .IN3(n6871), .IN4(n6870), .QN(n6874) );
  NAND2X0 U8841 ( .IN1(n7656), .IN2(n6872), .QN(n6873) );
  NAND4X0 U8842 ( .IN1(n6876), .IN2(n6875), .IN3(n6874), .IN4(n6873), .QN(
        \a3/N446 ) );
  NOR2X0 U8843 ( .IN1(n9213), .IN2(n7164), .QN(n6877) );
  AOI22X1 U8844 ( .IN1(n6877), .IN2(n8730), .IN3(n8395), .IN4(n9438), .QN(
        n6885) );
  INVX0 U8845 ( .INP(n8668), .ZN(n6881) );
  NOR2X0 U8846 ( .IN1(n7800), .IN2(n6878), .QN(n6880) );
  INVX0 U8847 ( .INP(n7727), .ZN(n8417) );
  NAND4X0 U8848 ( .IN1(n7862), .IN2(n8417), .IN3(n7287), .IN4(n7096), .QN(
        n6879) );
  NOR4X0 U8849 ( .IN1(n6882), .IN2(n6881), .IN3(n6880), .IN4(n6879), .QN(n6884) );
  NAND2X0 U8850 ( .IN1(n7656), .IN2(n6978), .QN(n7073) );
  NAND4X0 U8851 ( .IN1(n6885), .IN2(n6884), .IN3(n6883), .IN4(n7073), .QN(
        n6886) );
  OR4X1 U8852 ( .IN1(n8097), .IN2(n9092), .IN3(n7408), .IN4(n6886), .Q(
        \a3/N447 ) );
  NOR2X0 U8853 ( .IN1(n6887), .IN2(n6966), .QN(n6890) );
  OAI22X1 U8854 ( .IN1(n8754), .IN2(n6888), .IN3(n8188), .IN4(n9027), .QN(
        n6889) );
  NOR4X0 U8855 ( .IN1(n6891), .IN2(n8654), .IN3(n6890), .IN4(n6889), .QN(n6906) );
  INVX0 U8856 ( .INP(n6892), .ZN(n6902) );
  NOR2X0 U8857 ( .IN1(n7842), .IN2(n7812), .QN(n6900) );
  NAND2X0 U8858 ( .IN1(n9073), .IN2(n8780), .QN(n6894) );
  OA22X1 U8859 ( .IN1(n6895), .IN2(n8268), .IN3(n6894), .IN4(n6893), .Q(n6898)
         );
  INVX0 U8860 ( .INP(n6896), .ZN(n6897) );
  NAND4X0 U8861 ( .IN1(n6898), .IN2(n9088), .IN3(n7172), .IN4(n6897), .QN(
        n6899) );
  NOR4X0 U8862 ( .IN1(n6902), .IN2(n6901), .IN3(n6900), .IN4(n6899), .QN(n6905) );
  NAND4X0 U8863 ( .IN1(n6906), .IN2(n6905), .IN3(n6904), .IN4(n6903), .QN(
        \a3/N448 ) );
  NOR2X0 U8864 ( .IN1(degrees_tmp2[0]), .IN2(n8748), .QN(n8098) );
  NOR4X0 U8865 ( .IN1(n9176), .IN2(n8983), .IN3(n6907), .IN4(n8098), .QN(n6911) );
  OA22X1 U8866 ( .IN1(n8461), .IN2(n6908), .IN3(n9122), .IN4(n8084), .Q(n6910)
         );
  INVX0 U8867 ( .INP(n8358), .ZN(n8158) );
  NAND4X0 U8868 ( .IN1(n6911), .IN2(n6910), .IN3(n6909), .IN4(n8158), .QN(
        n6912) );
  NOR4X0 U8869 ( .IN1(n7355), .IN2(n6914), .IN3(n6913), .IN4(n6912), .QN(n6917) );
  OR2X1 U8870 ( .IN1(n7035), .IN2(n7685), .Q(n7791) );
  NAND4X0 U8871 ( .IN1(n6917), .IN2(n6916), .IN3(n6915), .IN4(n7791), .QN(
        \a3/N449 ) );
  INVX0 U8872 ( .INP(n6918), .ZN(n7960) );
  OA21X1 U8873 ( .IN1(n6919), .IN2(n8470), .IN3(n7960), .Q(n6933) );
  INVX0 U8874 ( .INP(n8850), .ZN(n6928) );
  NOR2X0 U8875 ( .IN1(n6920), .IN2(n7889), .QN(n6922) );
  OA22X1 U8876 ( .IN1(n6922), .IN2(n9149), .IN3(n6921), .IN4(n7749), .Q(n6926)
         );
  NAND3X0 U8877 ( .IN1(n9150), .IN2(n8649), .IN3(n9149), .QN(n6923) );
  NAND4X0 U8878 ( .IN1(n6926), .IN2(n6925), .IN3(n6924), .IN4(n6923), .QN(
        n6927) );
  NOR4X0 U8879 ( .IN1(n6930), .IN2(n6929), .IN3(n6928), .IN4(n6927), .QN(n6932) );
  NAND4X0 U8880 ( .IN1(n6933), .IN2(n6932), .IN3(n6931), .IN4(n8607), .QN(
        \a3/N450 ) );
  NAND2X0 U8881 ( .IN1(n6934), .IN2(n9442), .QN(n8509) );
  OA22X1 U8882 ( .IN1(n8667), .IN2(n8509), .IN3(n9166), .IN4(n7824), .Q(n6939)
         );
  INVX0 U8883 ( .INP(n7921), .ZN(n7123) );
  NOR2X0 U8884 ( .IN1(n8073), .IN2(n8171), .QN(n6935) );
  OA22X1 U8885 ( .IN1(n6936), .IN2(n7123), .IN3(n6935), .IN4(n8977), .Q(n6938)
         );
  NAND4X0 U8886 ( .IN1(n6939), .IN2(n6938), .IN3(n7856), .IN4(n6937), .QN(
        n6940) );
  NOR4X0 U8887 ( .IN1(n6942), .IN2(n6941), .IN3(n8629), .IN4(n6940), .QN(n6944) );
  AO221X1 U8888 ( .IN1(n9127), .IN2(n6968), .IN3(n9127), .IN4(n6967), .IN5(
        n8816), .Q(n6943) );
  NAND3X0 U8889 ( .IN1(n6944), .IN2(n8131), .IN3(n6943), .QN(\a3/N451 ) );
  NAND2X0 U8890 ( .IN1(n7973), .IN2(n9440), .QN(n7854) );
  NAND4X0 U8891 ( .IN1(n6945), .IN2(n7862), .IN3(n7951), .IN4(n7854), .QN(
        n6958) );
  NAND4X0 U8892 ( .IN1(n9210), .IN2(n6947), .IN3(n9019), .IN4(n6946), .QN(
        n6948) );
  NAND4X0 U8893 ( .IN1(n7111), .IN2(n6950), .IN3(n6949), .IN4(n6948), .QN(
        n6957) );
  NAND3X0 U8894 ( .IN1(n6952), .IN2(n6951), .IN3(n7746), .QN(n6953) );
  NAND2X0 U8895 ( .IN1(n6953), .IN2(n9155), .QN(n6954) );
  NAND4X0 U8896 ( .IN1(n7749), .IN2(n6955), .IN3(n9057), .IN4(n6954), .QN(
        n6956) );
  OR3X1 U8897 ( .IN1(n6958), .IN2(n6957), .IN3(n6956), .Q(\a3/N452 ) );
  INVX0 U8898 ( .INP(n7707), .ZN(n6960) );
  OA22X1 U8899 ( .IN1(n7184), .IN2(n6961), .IN3(n6960), .IN4(n6959), .Q(n6977)
         );
  NOR2X0 U8900 ( .IN1(n8574), .IN2(n7403), .QN(n7928) );
  INVX0 U8901 ( .INP(n8349), .ZN(n7896) );
  NAND2X0 U8902 ( .IN1(n7896), .IN2(n8494), .QN(n6964) );
  NAND3X0 U8903 ( .IN1(degrees_tmp2[5]), .IN2(n8485), .IN3(n8484), .QN(n6962)
         );
  NAND3X0 U8904 ( .IN1(n6964), .IN2(n6963), .IN3(n6962), .QN(n6973) );
  OA22X1 U8905 ( .IN1(n9149), .IN2(n6965), .IN3(n8229), .IN4(n9087), .Q(n6971)
         );
  NAND2X0 U8906 ( .IN1(n8567), .IN2(n9442), .QN(n7474) );
  OA22X1 U8907 ( .IN1(n6968), .IN2(n6967), .IN3(n6966), .IN4(n7474), .Q(n6970)
         );
  OA22X1 U8908 ( .IN1(n8471), .IN2(n8073), .IN3(n7679), .IN4(n8595), .Q(n6969)
         );
  NAND4X0 U8909 ( .IN1(n6971), .IN2(n6970), .IN3(n6969), .IN4(n8263), .QN(
        n6972) );
  NOR4X0 U8910 ( .IN1(n8066), .IN2(n7928), .IN3(n6973), .IN4(n6972), .QN(n6976) );
  NAND2X0 U8911 ( .IN1(n9189), .IN2(n6974), .QN(n7385) );
  NAND4X0 U8912 ( .IN1(n6977), .IN2(n6976), .IN3(n6975), .IN4(n7385), .QN(
        \a3/N453 ) );
  AOI22X1 U8913 ( .IN1(n6980), .IN2(n6979), .IN3(n6978), .IN4(n8588), .QN(
        n6995) );
  NOR2X0 U8914 ( .IN1(n9147), .IN2(n8563), .QN(n6992) );
  NAND2X0 U8915 ( .IN1(n7784), .IN2(n8496), .QN(n6981) );
  NAND4X0 U8916 ( .IN1(n6982), .IN2(n6981), .IN3(n7851), .IN4(n8248), .QN(
        n6991) );
  INVX0 U8917 ( .INP(n6983), .ZN(n6984) );
  NOR2X0 U8918 ( .IN1(n6984), .IN2(n9080), .QN(n6987) );
  NAND2X0 U8919 ( .IN1(n6985), .IN2(n7785), .QN(n6986) );
  NOR2X0 U8920 ( .IN1(n6987), .IN2(n6986), .QN(n6988) );
  NAND4X0 U8921 ( .IN1(n6989), .IN2(n6988), .IN3(n8657), .IN4(n7940), .QN(
        n6990) );
  NOR4X0 U8922 ( .IN1(n6993), .IN2(n6992), .IN3(n6991), .IN4(n6990), .QN(n6994) );
  NAND2X0 U8923 ( .IN1(n9053), .IN2(n7510), .QN(n7258) );
  NAND2X0 U8924 ( .IN1(n9037), .IN2(n7258), .QN(n7682) );
  NAND4X0 U8925 ( .IN1(n6995), .IN2(n6994), .IN3(n7259), .IN4(n7682), .QN(
        \a3/N454 ) );
  OA21X1 U8926 ( .IN1(degrees_tmp2[0]), .IN2(n6996), .IN3(n7240), .Q(n7007) );
  AO22X1 U8927 ( .IN1(degrees_tmp2[3]), .IN2(n7586), .IN3(n7484), .IN4(n7417), 
        .Q(n7001) );
  OA22X1 U8928 ( .IN1(n8876), .IN2(n9029), .IN3(n8169), .IN4(n8947), .Q(n6999)
         );
  INVX0 U8929 ( .INP(n8942), .ZN(n6998) );
  NAND2X0 U8930 ( .IN1(n9092), .IN2(n8041), .QN(n6997) );
  NAND4X0 U8931 ( .IN1(n6999), .IN2(n6998), .IN3(n8845), .IN4(n6997), .QN(
        n7000) );
  NOR4X0 U8932 ( .IN1(n7003), .IN2(n7002), .IN3(n7001), .IN4(n7000), .QN(n7006) );
  AO221X1 U8933 ( .IN1(n7004), .IN2(n9435), .IN3(n7004), .IN4(n8530), .IN5(
        n8229), .Q(n7005) );
  NAND4X0 U8934 ( .IN1(n7007), .IN2(n7006), .IN3(n8889), .IN4(n7005), .QN(
        \a3/N455 ) );
  INVX0 U8935 ( .INP(n9062), .ZN(n8602) );
  NOR2X0 U8936 ( .IN1(n9434), .IN2(n8602), .QN(n7651) );
  NOR2X0 U8937 ( .IN1(n7008), .IN2(n7651), .QN(n7020) );
  INVX0 U8938 ( .INP(n7009), .ZN(n7017) );
  INVX0 U8939 ( .INP(n7010), .ZN(n9133) );
  NOR2X0 U8940 ( .IN1(n7600), .IN2(n7969), .QN(n8006) );
  OA22X1 U8941 ( .IN1(n8598), .IN2(n8903), .IN3(n8533), .IN4(n7011), .Q(n7015)
         );
  INVX0 U8942 ( .INP(n9092), .ZN(n7014) );
  NAND2X0 U8943 ( .IN1(n7012), .IN2(n7142), .QN(n7013) );
  NAND4X0 U8944 ( .IN1(n7015), .IN2(n7014), .IN3(n8961), .IN4(n7013), .QN(
        n7016) );
  NOR4X0 U8945 ( .IN1(n7017), .IN2(n9133), .IN3(n8006), .IN4(n7016), .QN(n7019) );
  NAND4X0 U8946 ( .IN1(n7020), .IN2(n7019), .IN3(n7857), .IN4(n7018), .QN(
        n7021) );
  AO221X1 U8947 ( .IN1(n9434), .IN2(n7698), .IN3(n9434), .IN4(n8674), .IN5(
        n7021), .Q(\a3/N456 ) );
  INVX0 U8948 ( .INP(n7022), .ZN(n7030) );
  NOR2X0 U8949 ( .IN1(n7169), .IN2(n7023), .QN(n7029) );
  OA21X1 U8950 ( .IN1(n7572), .IN2(n7233), .IN3(n7024), .Q(n7027) );
  OA21X1 U8951 ( .IN1(n8444), .IN2(n8004), .IN3(n7364), .Q(n7026) );
  NAND4X0 U8952 ( .IN1(n7027), .IN2(n7026), .IN3(n7025), .IN4(n8845), .QN(
        n7028) );
  OR4X1 U8953 ( .IN1(n7031), .IN2(n7030), .IN3(n7029), .IN4(n7028), .Q(
        \a3/N457 ) );
  AND2X1 U8954 ( .IN1(n7032), .IN2(n8484), .Q(n7047) );
  OA22X1 U8955 ( .IN1(n8446), .IN2(n8707), .IN3(n9155), .IN4(n8977), .Q(n7045)
         );
  INVX0 U8956 ( .INP(n7187), .ZN(n7042) );
  OA21X1 U8957 ( .IN1(n7033), .IN2(n7142), .IN3(n9037), .Q(n7041) );
  NOR2X0 U8958 ( .IN1(n8229), .IN2(n7034), .QN(n7040) );
  NOR2X0 U8959 ( .IN1(n7035), .IN2(n7235), .QN(n7038) );
  NAND2X0 U8960 ( .IN1(n7036), .IN2(n8467), .QN(n7037) );
  NOR2X0 U8961 ( .IN1(n7038), .IN2(n7037), .QN(n7039) );
  NOR4X0 U8962 ( .IN1(n7042), .IN2(n7041), .IN3(n7040), .IN4(n7039), .QN(n7044) );
  NAND3X0 U8963 ( .IN1(n9182), .IN2(degrees_tmp2[0]), .IN3(n7686), .QN(n7043)
         );
  NAND4X0 U8964 ( .IN1(n7045), .IN2(n7044), .IN3(n7288), .IN4(n7043), .QN(
        n7046) );
  OR4X1 U8965 ( .IN1(n8718), .IN2(n9187), .IN3(n7047), .IN4(n7046), .Q(
        \a3/N458 ) );
  INVX0 U8966 ( .INP(n7254), .ZN(n8523) );
  NAND2X0 U8967 ( .IN1(degrees_tmp2[0]), .IN2(n7686), .QN(n7048) );
  OA22X1 U8968 ( .IN1(n8847), .IN2(n8523), .IN3(n8684), .IN4(n7048), .Q(n7056)
         );
  AO21X1 U8969 ( .IN1(n7049), .IN2(n9195), .IN3(n8324), .Q(n7101) );
  NAND2X0 U8970 ( .IN1(n8301), .IN2(n7050), .QN(n9085) );
  AND3X1 U8971 ( .IN1(n9213), .IN2(n8124), .IN3(n7051), .Q(n7052) );
  OA22X1 U8972 ( .IN1(n8533), .IN2(n9085), .IN3(n7052), .IN4(n7800), .Q(n7053)
         );
  NAND4X0 U8973 ( .IN1(n7053), .IN2(n8869), .IN3(n7781), .IN4(n7368), .QN(
        n7054) );
  NOR2X0 U8974 ( .IN1(n7101), .IN2(n7054), .QN(n7055) );
  NAND4X0 U8975 ( .IN1(n7056), .IN2(n7055), .IN3(n8555), .IN4(n8042), .QN(
        \a3/N459 ) );
  NAND2X0 U8976 ( .IN1(n9435), .IN2(n8883), .QN(n7059) );
  OA22X1 U8977 ( .IN1(n7391), .IN2(n7059), .IN3(n7058), .IN4(n7057), .Q(n7068)
         );
  AOI21X1 U8978 ( .IN1(n8823), .IN2(n8861), .IN3(n8985), .QN(n7067) );
  NAND2X0 U8979 ( .IN1(degrees_tmp2[2]), .IN2(n8774), .QN(n8295) );
  NAND2X0 U8980 ( .IN1(n8529), .IN2(n9099), .QN(n7551) );
  NAND4X0 U8981 ( .IN1(n7495), .IN2(n8295), .IN3(n7636), .IN4(n7551), .QN(
        n7062) );
  NAND2X0 U8982 ( .IN1(n7483), .IN2(n7760), .QN(n7449) );
  NAND4X0 U8983 ( .IN1(n7060), .IN2(n9020), .IN3(n8850), .IN4(n7449), .QN(
        n7061) );
  NOR4X0 U8984 ( .IN1(n7064), .IN2(n7063), .IN3(n7062), .IN4(n7061), .QN(n7066) );
  NAND4X0 U8985 ( .IN1(n7068), .IN2(n7067), .IN3(n7066), .IN4(n7065), .QN(
        \a3/N460 ) );
  NOR2X0 U8986 ( .IN1(n7282), .IN2(n8862), .QN(n7069) );
  OA22X1 U8987 ( .IN1(n7069), .IN2(n8588), .IN3(n7913), .IN4(n9119), .Q(n7080)
         );
  NOR2X0 U8988 ( .IN1(n7070), .IN2(n8572), .QN(n7072) );
  NAND2X0 U8989 ( .IN1(n8615), .IN2(n7113), .QN(n7071) );
  NOR2X0 U8990 ( .IN1(n7072), .IN2(n7071), .QN(n7079) );
  NOR2X0 U8991 ( .IN1(n8752), .IN2(n7839), .QN(n8286) );
  NAND2X0 U8992 ( .IN1(n8696), .IN2(n8731), .QN(n7074) );
  NAND3X0 U8993 ( .IN1(n7074), .IN2(n7073), .IN3(n7641), .QN(n7076) );
  OAI22X1 U8994 ( .IN1(n9131), .IN2(n7875), .IN3(n7572), .IN4(n8531), .QN(
        n7075) );
  NOR4X0 U8995 ( .IN1(n8286), .IN2(n7077), .IN3(n7076), .IN4(n7075), .QN(n7078) );
  NAND4X0 U8996 ( .IN1(n7080), .IN2(n7079), .IN3(n7078), .IN4(n8869), .QN(
        \a3/N461 ) );
  NAND2X0 U8997 ( .IN1(degrees_tmp2[5]), .IN2(n7081), .QN(n7992) );
  AND2X1 U8998 ( .IN1(n7992), .IN2(n7943), .Q(n7967) );
  NOR2X0 U8999 ( .IN1(n9031), .IN2(n8968), .QN(n7089) );
  NAND4X0 U9000 ( .IN1(n8504), .IN2(n7241), .IN3(n8100), .IN4(n7082), .QN(
        n7088) );
  OA22X1 U9001 ( .IN1(n7084), .IN2(n7638), .IN3(n7083), .IN4(n7388), .Q(n7086)
         );
  NAND3X0 U9002 ( .IN1(n8788), .IN2(n8474), .IN3(n9032), .QN(n7370) );
  OAI21X1 U9003 ( .IN1(n8058), .IN2(n8330), .IN3(n8467), .QN(n7085) );
  NAND4X0 U9004 ( .IN1(n8116), .IN2(n7086), .IN3(n7370), .IN4(n7085), .QN(
        n7087) );
  NOR4X0 U9005 ( .IN1(n7090), .IN2(n7089), .IN3(n7088), .IN4(n7087), .QN(n7092) );
  NAND4X0 U9006 ( .IN1(n7967), .IN2(n7092), .IN3(n7091), .IN4(n7771), .QN(
        \a3/N462 ) );
  NOR2X0 U9007 ( .IN1(n9436), .IN2(n9099), .QN(n7624) );
  OA21X1 U9008 ( .IN1(n7451), .IN2(n7624), .IN3(n7093), .Q(n7103) );
  NAND2X0 U9009 ( .IN1(n9033), .IN2(n7094), .QN(n7095) );
  NAND4X0 U9010 ( .IN1(n7494), .IN2(n7787), .IN3(n7096), .IN4(n7095), .QN(
        n7102) );
  INVX0 U9011 ( .INP(n8178), .ZN(n7098) );
  NAND4X0 U9012 ( .IN1(n7099), .IN2(n7098), .IN3(n7797), .IN4(n7097), .QN(
        n7100) );
  NOR4X0 U9013 ( .IN1(n7103), .IN2(n7102), .IN3(n7101), .IN4(n7100), .QN(n7105) );
  INVX0 U9014 ( .INP(n8436), .ZN(n9193) );
  NAND4X0 U9015 ( .IN1(n7105), .IN2(n8820), .IN3(n9193), .IN4(n7104), .QN(
        \a3/N463 ) );
  OA221X1 U9016 ( .IN1(n8787), .IN2(n8693), .IN3(n8787), .IN4(n8564), .IN5(
        n7106), .Q(n7117) );
  NOR2X0 U9017 ( .IN1(n9437), .IN2(n7107), .QN(n7692) );
  OA21X1 U9018 ( .IN1(n7108), .IN2(n7692), .IN3(n7298), .Q(n7115) );
  AO21X1 U9019 ( .IN1(n9212), .IN2(n7657), .IN3(n8787), .Q(n9016) );
  OA22X1 U9020 ( .IN1(n9195), .IN2(n7109), .IN3(n9441), .IN4(n9438), .Q(n7110)
         );
  NAND2X0 U9021 ( .IN1(n9208), .IN2(n7110), .QN(n7112) );
  NAND4X0 U9022 ( .IN1(n9016), .IN2(n7113), .IN3(n7112), .IN4(n7111), .QN(
        n7114) );
  NOR4X0 U9023 ( .IN1(n8786), .IN2(n7115), .IN3(n7795), .IN4(n7114), .QN(n7116) );
  INVX0 U9024 ( .INP(n7296), .ZN(n8911) );
  NAND4X0 U9025 ( .IN1(n7117), .IN2(n7116), .IN3(n8183), .IN4(n8911), .QN(
        \a3/N464 ) );
  INVX0 U9026 ( .INP(n7118), .ZN(n7120) );
  NOR2X0 U9027 ( .IN1(n7120), .IN2(n7119), .QN(n8373) );
  NOR2X0 U9028 ( .IN1(n8977), .IN2(n9045), .QN(n8944) );
  OA21X1 U9029 ( .IN1(n8753), .IN2(n7121), .IN3(n9099), .Q(n7126) );
  OA22X1 U9030 ( .IN1(n8752), .IN2(n7538), .IN3(n7252), .IN4(n7234), .Q(n7124)
         );
  NAND2X0 U9031 ( .IN1(n8567), .IN2(n9173), .QN(n7122) );
  NAND4X0 U9032 ( .IN1(n7124), .IN2(n7123), .IN3(n8819), .IN4(n7122), .QN(
        n7125) );
  NOR4X0 U9033 ( .IN1(n8953), .IN2(n8944), .IN3(n7126), .IN4(n7125), .QN(n7128) );
  NAND4X0 U9034 ( .IN1(n8373), .IN2(n7128), .IN3(n8406), .IN4(n7127), .QN(
        \a3/N465 ) );
  AOI22X1 U9035 ( .IN1(n8731), .IN2(n7451), .IN3(n7436), .IN4(n8431), .QN(
        n7141) );
  NAND2X0 U9036 ( .IN1(n9182), .IN2(n9084), .QN(n8672) );
  NAND2X0 U9037 ( .IN1(n8268), .IN2(n8672), .QN(n7130) );
  AO22X1 U9038 ( .IN1(n9037), .IN2(n7130), .IN3(n7129), .IN4(n9445), .Q(n7138)
         );
  NAND3X0 U9039 ( .IN1(n7394), .IN2(n7131), .IN3(n8265), .QN(n7137) );
  NOR2X0 U9040 ( .IN1(n8816), .IN2(n8859), .QN(n7132) );
  NOR2X0 U9041 ( .IN1(n8622), .IN2(n7132), .QN(n7983) );
  NAND2X0 U9042 ( .IN1(n9434), .IN2(n7133), .QN(n7811) );
  NAND2X0 U9043 ( .IN1(degrees_tmp2[2]), .IN2(n7134), .QN(n7135) );
  NAND4X0 U9044 ( .IN1(n7983), .IN2(n8720), .IN3(n7811), .IN4(n7135), .QN(
        n7136) );
  NOR4X0 U9045 ( .IN1(n7139), .IN2(n7138), .IN3(n7137), .IN4(n7136), .QN(n7140) );
  NAND4X0 U9046 ( .IN1(n7141), .IN2(n7140), .IN3(n8778), .IN4(n8541), .QN(
        \a3/N466 ) );
  INVX0 U9047 ( .INP(n7142), .ZN(n7144) );
  OA22X1 U9048 ( .IN1(n9183), .IN2(n8880), .IN3(n7144), .IN4(n7143), .Q(n7152)
         );
  NAND2X0 U9049 ( .IN1(n8875), .IN2(n8987), .QN(n7145) );
  NAND4X0 U9050 ( .IN1(n8866), .IN2(n7828), .IN3(n8618), .IN4(n7145), .QN(
        n7149) );
  AO21X1 U9051 ( .IN1(n9436), .IN2(n7147), .IN3(n7146), .Q(n7148) );
  NOR4X0 U9052 ( .IN1(n7692), .IN2(n8953), .IN3(n7149), .IN4(n7148), .QN(n7151) );
  NAND3X0 U9053 ( .IN1(n8788), .IN2(n9061), .IN3(n8692), .QN(n7150) );
  NAND4X0 U9054 ( .IN1(n7153), .IN2(n7152), .IN3(n7151), .IN4(n7150), .QN(
        \a3/N467 ) );
  NAND2X0 U9055 ( .IN1(n9087), .IN2(n8410), .QN(n8949) );
  INVX0 U9056 ( .INP(n7528), .ZN(n9004) );
  OAI22X1 U9057 ( .IN1(n8401), .IN2(n9004), .IN3(n7890), .IN4(n9434), .QN(
        n7159) );
  OA21X1 U9058 ( .IN1(n7155), .IN2(n9442), .IN3(n7154), .Q(n7157) );
  NAND4X0 U9059 ( .IN1(n7157), .IN2(n7156), .IN3(n8820), .IN4(n8747), .QN(
        n7158) );
  NOR4X0 U9060 ( .IN1(n7160), .IN2(n8949), .IN3(n7159), .IN4(n7158), .QN(n7163) );
  NAND2X0 U9061 ( .IN1(n9080), .IN2(n7161), .QN(n7162) );
  NAND4X0 U9062 ( .IN1(n7163), .IN2(n8713), .IN3(n9118), .IN4(n7162), .QN(
        \a3/N468 ) );
  NAND2X0 U9063 ( .IN1(n7816), .IN2(n8645), .QN(n7687) );
  OA22X1 U9064 ( .IN1(n9438), .IN2(n7165), .IN3(n7164), .IN4(n7687), .Q(n7178)
         );
  NAND3X0 U9065 ( .IN1(n7167), .IN2(n8675), .IN3(n9181), .QN(n8114) );
  OA22X1 U9066 ( .IN1(n8816), .IN2(n8114), .IN3(n7166), .IN4(n7233), .Q(n7177)
         );
  INVX0 U9067 ( .INP(n7167), .ZN(n7553) );
  OA22X1 U9068 ( .IN1(n8876), .IN2(n7168), .IN3(n7650), .IN4(n7553), .Q(n7175)
         );
  OR2X1 U9069 ( .IN1(n8246), .IN2(n7169), .Q(n8383) );
  NAND2X0 U9070 ( .IN1(degrees_tmp2[5]), .IN2(n7170), .QN(n7171) );
  AND4X1 U9071 ( .IN1(n9111), .IN2(n7172), .IN3(n8383), .IN4(n7171), .Q(n7173)
         );
  OA221X1 U9072 ( .IN1(n8026), .IN2(n7175), .IN3(n8026), .IN4(n7174), .IN5(
        n7173), .Q(n7176) );
  NAND4X0 U9073 ( .IN1(n7178), .IN2(n7177), .IN3(n7176), .IN4(n8202), .QN(
        \a3/N469 ) );
  INVX0 U9074 ( .INP(n7179), .ZN(n7180) );
  OA22X1 U9075 ( .IN1(degrees_tmp2[5]), .IN2(n7181), .IN3(n9083), .IN4(n7180), 
        .Q(n7194) );
  NAND2X0 U9076 ( .IN1(n8996), .IN2(n8452), .QN(n7191) );
  OA22X1 U9077 ( .IN1(n7184), .IN2(n7183), .IN3(n8531), .IN4(n7182), .Q(n7185)
         );
  OA21X1 U9078 ( .IN1(degrees_tmp2[3]), .IN2(n8705), .IN3(n7185), .Q(n7189) );
  NAND2X0 U9079 ( .IN1(n8171), .IN2(n8033), .QN(n7186) );
  NAND4X0 U9080 ( .IN1(n7189), .IN2(n7188), .IN3(n7187), .IN4(n7186), .QN(
        n7190) );
  NOR4X0 U9081 ( .IN1(n7192), .IN2(n7728), .IN3(n7191), .IN4(n7190), .QN(n7193) );
  NAND4X0 U9082 ( .IN1(n7194), .IN2(n7193), .IN3(n7587), .IN4(n7224), .QN(
        \a3/N471 ) );
  OA22X1 U9083 ( .IN1(n7736), .IN2(n8204), .IN3(n7234), .IN4(n9099), .Q(n7207)
         );
  NAND2X0 U9084 ( .IN1(n7195), .IN2(n9026), .QN(n8867) );
  NAND4X0 U9085 ( .IN1(n8851), .IN2(n9110), .IN3(n8265), .IN4(n8867), .QN(
        n7202) );
  INVX0 U9086 ( .INP(n8641), .ZN(n7196) );
  NOR2X0 U9087 ( .IN1(n7197), .IN2(n7196), .QN(n7200) );
  NAND3X0 U9088 ( .IN1(degrees_tmp2[5]), .IN2(n7198), .IN3(n8171), .QN(n7199)
         );
  NAND4X0 U9089 ( .IN1(n7200), .IN2(n8007), .IN3(n7968), .IN4(n7199), .QN(
        n7201) );
  NOR4X0 U9090 ( .IN1(n7204), .IN2(n7203), .IN3(n7202), .IN4(n7201), .QN(n7206) );
  NAND4X0 U9091 ( .IN1(n7207), .IN2(n7206), .IN3(n7787), .IN4(n7205), .QN(
        \a3/N472 ) );
  INVX0 U9092 ( .INP(n7208), .ZN(n7210) );
  OA22X1 U9093 ( .IN1(n7211), .IN2(n8282), .IN3(n7210), .IN4(n7209), .Q(n7220)
         );
  INVX0 U9094 ( .INP(n7408), .ZN(n7212) );
  OA21X1 U9095 ( .IN1(n8883), .IN2(n9002), .IN3(n7212), .Q(n7219) );
  AO22X1 U9096 ( .IN1(n9182), .IN2(n7879), .IN3(n7214), .IN4(n7213), .Q(n7216)
         );
  NAND2X0 U9097 ( .IN1(n7294), .IN2(n9006), .QN(n7215) );
  NOR4X0 U9098 ( .IN1(n8111), .IN2(n7217), .IN3(n7216), .IN4(n7215), .QN(n7218) );
  NAND4X0 U9099 ( .IN1(n7220), .IN2(n7219), .IN3(n7218), .IN4(n8126), .QN(
        \a3/N473 ) );
  OA21X1 U9100 ( .IN1(n7222), .IN2(n7221), .IN3(degrees_tmp2[0]), .Q(n7232) );
  OR2X1 U9101 ( .IN1(n7223), .IN2(n9437), .Q(n7396) );
  NAND4X0 U9102 ( .IN1(n7225), .IN2(n7458), .IN3(n7224), .IN4(n7396), .QN(
        n7230) );
  OA22X1 U9103 ( .IN1(n8510), .IN2(n7714), .IN3(n8760), .IN4(n8815), .Q(n7228)
         );
  INVX0 U9104 ( .INP(n8162), .ZN(n7226) );
  AND4X1 U9105 ( .IN1(n7226), .IN2(n8835), .IN3(n8412), .IN4(n8967), .Q(n7227)
         );
  NAND4X0 U9106 ( .IN1(n7228), .IN2(n7227), .IN3(n8053), .IN4(n7245), .QN(
        n7229) );
  OR4X1 U9107 ( .IN1(n7232), .IN2(n7231), .IN3(n7230), .IN4(n7229), .Q(
        \a3/N474 ) );
  OA22X1 U9108 ( .IN1(n8598), .IN2(n8550), .IN3(n7234), .IN4(n7233), .Q(n7247)
         );
  NAND2X0 U9109 ( .IN1(n9175), .IN2(n9166), .QN(n8547) );
  NAND2X0 U9110 ( .IN1(n7235), .IN2(n7686), .QN(n8503) );
  NAND4X0 U9111 ( .IN1(n8922), .IN2(n8547), .IN3(n8503), .IN4(n7839), .QN(
        n7237) );
  OA221X1 U9112 ( .IN1(n7237), .IN2(n8710), .IN3(n7237), .IN4(n7236), .IN5(
        degrees_tmp2[2]), .Q(n7244) );
  INVX0 U9113 ( .INP(n7238), .ZN(n8140) );
  OA22X1 U9114 ( .IN1(n8140), .IN2(n8921), .IN3(n9147), .IN4(n8303), .Q(n7242)
         );
  NAND2X0 U9115 ( .IN1(n7735), .IN2(n7239), .QN(n8736) );
  NAND4X0 U9116 ( .IN1(n7242), .IN2(n7241), .IN3(n7240), .IN4(n8736), .QN(
        n7243) );
  NOR2X0 U9117 ( .IN1(n7244), .IN2(n7243), .QN(n7246) );
  NAND4X0 U9118 ( .IN1(n7247), .IN2(n7246), .IN3(n7245), .IN4(n8412), .QN(
        \a3/N475 ) );
  NOR2X0 U9119 ( .IN1(n9442), .IN2(n8651), .QN(n7249) );
  NAND2X0 U9120 ( .IN1(n7474), .IN2(n8576), .QN(n7248) );
  NOR2X0 U9121 ( .IN1(n7249), .IN2(n7248), .QN(n7268) );
  OA221X1 U9122 ( .IN1(n7250), .IN2(n8753), .IN3(n7250), .IN4(n8489), .IN5(
        n9433), .Q(n7253) );
  NAND2X0 U9123 ( .IN1(n8289), .IN2(n9438), .QN(n8702) );
  NOR2X0 U9124 ( .IN1(n7252), .IN2(n7251), .QN(n9144) );
  INVX0 U9125 ( .INP(n9144), .ZN(n8003) );
  NAND2X0 U9126 ( .IN1(n8702), .IN2(n8003), .QN(n9174) );
  NOR2X0 U9127 ( .IN1(n7253), .IN2(n9174), .QN(n7267) );
  NAND2X0 U9128 ( .IN1(degrees_tmp2[3]), .IN2(n7254), .QN(n7255) );
  NAND3X0 U9129 ( .IN1(n7257), .IN2(n7256), .IN3(n7255), .QN(n7262) );
  NAND2X0 U9130 ( .IN1(n8883), .IN2(n7258), .QN(n7260) );
  NAND3X0 U9131 ( .IN1(n7260), .IN2(n7259), .IN3(n8743), .QN(n7261) );
  NOR4X0 U9132 ( .IN1(n7264), .IN2(n7263), .IN3(n7262), .IN4(n7261), .QN(n7266) );
  NAND4X0 U9133 ( .IN1(n7268), .IN2(n7267), .IN3(n7266), .IN4(n7265), .QN(
        \a3/N476 ) );
  INVX0 U9134 ( .INP(n7269), .ZN(n8021) );
  NAND2X0 U9135 ( .IN1(n7654), .IN2(n9147), .QN(n7270) );
  AND4X1 U9136 ( .IN1(n8021), .IN2(n7302), .IN3(n7287), .IN4(n7270), .Q(n7280)
         );
  OA22X1 U9137 ( .IN1(n7880), .IN2(n8967), .IN3(n7736), .IN4(n7510), .Q(n7279)
         );
  INVX0 U9138 ( .INP(n7771), .ZN(n7541) );
  OA21X1 U9139 ( .IN1(n8823), .IN2(n7506), .IN3(n8595), .Q(n7276) );
  NAND3X0 U9140 ( .IN1(n9125), .IN2(n8640), .IN3(n7271), .QN(n7272) );
  NAND4X0 U9141 ( .IN1(n7274), .IN2(n7330), .IN3(n7273), .IN4(n7272), .QN(
        n7275) );
  NOR4X0 U9142 ( .IN1(n7541), .IN2(n7277), .IN3(n7276), .IN4(n7275), .QN(n7278) );
  NAND4X0 U9143 ( .IN1(n7280), .IN2(n7279), .IN3(n7278), .IN4(n8292), .QN(
        \a3/N477 ) );
  OA22X1 U9144 ( .IN1(n8511), .IN2(n8880), .IN3(n8073), .IN4(n8422), .Q(n7290)
         );
  NOR3X0 U9145 ( .IN1(n7391), .IN2(n7945), .IN3(n7800), .QN(n7286) );
  OA21X1 U9146 ( .IN1(n7281), .IN2(n8718), .IN3(n8692), .Q(n7285) );
  INVX0 U9147 ( .INP(n8156), .ZN(n7339) );
  AO21X1 U9148 ( .IN1(n7282), .IN2(n8764), .IN3(n7339), .Q(n7826) );
  INVX0 U9149 ( .INP(n7425), .ZN(n7283) );
  NAND4X0 U9150 ( .IN1(n7558), .IN2(n7283), .IN3(n8578), .IN4(n8747), .QN(
        n7284) );
  NOR4X0 U9151 ( .IN1(n7286), .IN2(n7285), .IN3(n7826), .IN4(n7284), .QN(n7289) );
  NAND4X0 U9152 ( .IN1(n7290), .IN2(n7289), .IN3(n7288), .IN4(n7287), .QN(
        \a3/N478 ) );
  NOR2X0 U9153 ( .IN1(n7437), .IN2(n8947), .QN(n7292) );
  OA22X1 U9154 ( .IN1(n8995), .IN2(n7293), .IN3(n7292), .IN4(n7291), .Q(n7310)
         );
  INVX0 U9155 ( .INP(n7294), .ZN(n7295) );
  OA21X1 U9156 ( .IN1(n7295), .IN2(n7582), .IN3(n8188), .Q(n7306) );
  NOR4X0 U9157 ( .IN1(n8379), .IN2(n7297), .IN3(n7296), .IN4(n8483), .QN(n7304) );
  OA22X1 U9158 ( .IN1(n9433), .IN2(n7299), .IN3(n7298), .IN4(n8695), .Q(n7303)
         );
  NAND2X0 U9159 ( .IN1(n8727), .IN2(n7300), .QN(n7301) );
  NAND4X0 U9160 ( .IN1(n7304), .IN2(n7303), .IN3(n7302), .IN4(n7301), .QN(
        n7305) );
  NOR3X0 U9161 ( .IN1(n8094), .IN2(n7306), .IN3(n7305), .QN(n7309) );
  NAND4X0 U9162 ( .IN1(n7310), .IN2(n7309), .IN3(n7308), .IN4(n7307), .QN(
        \a3/N479 ) );
  OA22X1 U9163 ( .IN1(n9080), .IN2(n7510), .IN3(n8262), .IN4(n9032), .Q(n7319)
         );
  NOR2X0 U9164 ( .IN1(n8883), .IN2(n8800), .QN(n7315) );
  NAND2X0 U9165 ( .IN1(n7311), .IN2(n8004), .QN(n8617) );
  NAND2X0 U9166 ( .IN1(n7668), .IN2(n7312), .QN(n7323) );
  NAND4X0 U9167 ( .IN1(n8571), .IN2(n8366), .IN3(n8617), .IN4(n7323), .QN(
        n7314) );
  NAND2X0 U9168 ( .IN1(n9203), .IN2(n9208), .QN(n7840) );
  NAND4X0 U9169 ( .IN1(n8069), .IN2(n9140), .IN3(n8410), .IN4(n7840), .QN(
        n7313) );
  NOR4X0 U9170 ( .IN1(n8407), .IN2(n7315), .IN3(n7314), .IN4(n7313), .QN(n7318) );
  AO221X1 U9171 ( .IN1(n7316), .IN2(degrees_tmp2[0]), .IN3(n7316), .IN4(n8772), 
        .IN5(n9442), .Q(n7317) );
  OR2X1 U9172 ( .IN1(n7721), .IN2(n9437), .Q(n8973) );
  NAND4X0 U9173 ( .IN1(n7319), .IN2(n7318), .IN3(n7317), .IN4(n8973), .QN(
        \a3/N480 ) );
  INVX0 U9174 ( .INP(n7320), .ZN(n7658) );
  NAND4X0 U9175 ( .IN1(n8677), .IN2(n7829), .IN3(n7658), .IN4(n8790), .QN(
        n7329) );
  NAND2X0 U9176 ( .IN1(n7321), .IN2(n7473), .QN(n7324) );
  NAND3X0 U9177 ( .IN1(n7324), .IN2(n7323), .IN3(n7322), .QN(n7328) );
  NAND2X0 U9178 ( .IN1(n7806), .IN2(n7686), .QN(n7325) );
  NAND2X0 U9179 ( .IN1(degrees_tmp2[3]), .IN2(n7477), .QN(n7603) );
  NAND3X0 U9180 ( .IN1(n7326), .IN2(n7325), .IN3(n7603), .QN(n7327) );
  NOR4X0 U9181 ( .IN1(n7804), .IN2(n7329), .IN3(n7328), .IN4(n7327), .QN(n7332) );
  OR2X1 U9182 ( .IN1(n8026), .IN2(n7840), .Q(n8865) );
  NAND4X0 U9183 ( .IN1(n7332), .IN2(n7331), .IN3(n7330), .IN4(n8865), .QN(
        \a3/N481 ) );
  AOI21X1 U9184 ( .IN1(n8778), .IN2(n8315), .IN3(n9082), .QN(n7337) );
  INVX0 U9185 ( .INP(n7333), .ZN(n8625) );
  NAND4X0 U9186 ( .IN1(n8625), .IN2(n7335), .IN3(n8503), .IN4(n7334), .QN(
        n7336) );
  NOR4X0 U9187 ( .IN1(n7339), .IN2(n7338), .IN3(n7337), .IN4(n7336), .QN(n7346) );
  NAND3X0 U9188 ( .IN1(n8701), .IN2(n7558), .IN3(n7340), .QN(n7341) );
  NAND2X0 U9189 ( .IN1(n7341), .IN2(n8041), .QN(n7344) );
  NAND2X0 U9190 ( .IN1(n7342), .IN2(n9060), .QN(n7343) );
  NAND4X0 U9191 ( .IN1(n7346), .IN2(n7345), .IN3(n7344), .IN4(n7343), .QN(
        \a3/N482 ) );
  OA21X1 U9192 ( .IN1(n8978), .IN2(n7347), .IN3(n8937), .Q(n7348) );
  OA22X1 U9193 ( .IN1(n8796), .IN2(n7349), .IN3(n7348), .IN4(n7736), .Q(n7357)
         );
  OAI21X1 U9194 ( .IN1(n8424), .IN2(n8303), .IN3(n8381), .QN(n7353) );
  NAND2X0 U9195 ( .IN1(n8753), .IN2(n8675), .QN(n7350) );
  NAND4X0 U9196 ( .IN1(n7351), .IN2(n9002), .IN3(n7771), .IN4(n7350), .QN(
        n7352) );
  NOR4X0 U9197 ( .IN1(n7355), .IN2(n7354), .IN3(n7353), .IN4(n7352), .QN(n7356) );
  NAND4X0 U9198 ( .IN1(n7357), .IN2(n7356), .IN3(n8664), .IN4(n8263), .QN(
        \a3/N483 ) );
  NOR3X0 U9199 ( .IN1(n7360), .IN2(n7359), .IN3(n7358), .QN(n7361) );
  NOR2X0 U9200 ( .IN1(n7361), .IN2(n7745), .QN(n7375) );
  OA21X1 U9201 ( .IN1(n9131), .IN2(n9192), .IN3(n7362), .Q(n7365) );
  NAND4X0 U9202 ( .IN1(n7365), .IN2(n7364), .IN3(n7363), .IN4(n7658), .QN(
        n7373) );
  NOR2X0 U9203 ( .IN1(n7655), .IN2(n9108), .QN(n7367) );
  NOR2X0 U9204 ( .IN1(n7367), .IN2(n7366), .QN(n7371) );
  NAND4X0 U9205 ( .IN1(n7371), .IN2(n7370), .IN3(n7369), .IN4(n7368), .QN(
        n7372) );
  OR4X1 U9206 ( .IN1(n7375), .IN2(n7374), .IN3(n7373), .IN4(n7372), .Q(
        \a3/N484 ) );
  AO21X1 U9207 ( .IN1(n9041), .IN2(n7376), .IN3(n9445), .Q(n8011) );
  NAND4X0 U9208 ( .IN1(n7379), .IN2(n7378), .IN3(n7377), .IN4(n8021), .QN(
        n7384) );
  OA21X1 U9209 ( .IN1(n8710), .IN2(n8281), .IN3(n8702), .Q(n7382) );
  NAND2X0 U9210 ( .IN1(n9080), .IN2(n8305), .QN(n7380) );
  NAND4X0 U9211 ( .IN1(n7382), .IN2(n8747), .IN3(n7381), .IN4(n7380), .QN(
        n7383) );
  NOR2X0 U9212 ( .IN1(n7384), .IN2(n7383), .QN(n7387) );
  NAND4X0 U9213 ( .IN1(n8011), .IN2(n7387), .IN3(n7386), .IN4(n7385), .QN(
        \a3/N485 ) );
  OA221X1 U9214 ( .IN1(n9196), .IN2(n7686), .IN3(n9196), .IN4(n7388), .IN5(
        n8892), .Q(n7401) );
  INVX0 U9215 ( .INP(n7389), .ZN(n7390) );
  OA22X1 U9216 ( .IN1(n8667), .IN2(n7392), .IN3(n7391), .IN4(n7390), .Q(n7400)
         );
  NOR2X0 U9217 ( .IN1(n7393), .IN2(n9073), .QN(n7398) );
  NOR2X0 U9218 ( .IN1(n9438), .IN2(n8349), .QN(n8884) );
  NOR2X0 U9219 ( .IN1(n9445), .IN2(n7823), .QN(n8637) );
  NOR2X0 U9220 ( .IN1(n8884), .IN2(n8637), .QN(n8012) );
  OA221X1 U9221 ( .IN1(n8727), .IN2(n7394), .IN3(n8727), .IN4(n9129), .IN5(
        n8012), .Q(n7395) );
  NAND2X0 U9222 ( .IN1(n7396), .IN2(n7395), .QN(n7397) );
  NOR2X0 U9223 ( .IN1(n7398), .IN2(n7397), .QN(n7399) );
  NAND4X0 U9224 ( .IN1(n7401), .IN2(n7400), .IN3(n7399), .IN4(n7495), .QN(
        \a3/N486 ) );
  OA22X1 U9225 ( .IN1(n7404), .IN2(n7403), .IN3(n7402), .IN4(n8597), .Q(n7410)
         );
  OA21X1 U9226 ( .IN1(n8697), .IN2(n7421), .IN3(n8947), .Q(n7407) );
  AO22X1 U9227 ( .IN1(n8848), .IN2(n7405), .IN3(n8728), .IN4(n9025), .Q(n7406)
         );
  NOR4X0 U9228 ( .IN1(n8407), .IN2(n7408), .IN3(n7407), .IN4(n7406), .QN(n7409) );
  NAND4X0 U9229 ( .IN1(n7410), .IN2(n7409), .IN3(n8851), .IN4(n8546), .QN(
        n7411) );
  AO221X1 U9230 ( .IN1(n9099), .IN2(n7413), .IN3(n9099), .IN4(n7412), .IN5(
        n7411), .Q(\a3/N487 ) );
  NOR2X0 U9231 ( .IN1(n7415), .IN2(n7414), .QN(n9201) );
  NOR2X0 U9232 ( .IN1(n7417), .IN2(n7416), .QN(n7418) );
  NOR4X0 U9233 ( .IN1(n9182), .IN2(n9014), .IN3(n9176), .IN4(n7418), .QN(n7419) );
  NAND4X0 U9234 ( .IN1(n9201), .IN2(n7420), .IN3(n7419), .IN4(n8799), .QN(
        \a3/N488 ) );
  NAND2X0 U9235 ( .IN1(n8598), .IN2(n7421), .QN(n7423) );
  NAND3X0 U9236 ( .IN1(n7423), .IN2(n8209), .IN3(n7422), .QN(\a3/N489 ) );
  OA21X1 U9237 ( .IN1(n8220), .IN2(\a3/N492 ), .IN3(quad[0]), .Q(\a3/N493 ) );
  OA22X1 U9238 ( .IN1(n7424), .IN2(n7822), .IN3(n8947), .IN4(n9020), .Q(n7442)
         );
  NOR2X0 U9239 ( .IN1(n7425), .IN2(n9039), .QN(n7427) );
  NAND2X0 U9240 ( .IN1(degrees_tmp2[0]), .IN2(n8993), .QN(n7426) );
  NAND2X0 U9241 ( .IN1(n7427), .IN2(n7426), .QN(n7433) );
  NAND2X0 U9242 ( .IN1(n7428), .IN2(n9147), .QN(n7429) );
  NAND4X0 U9243 ( .IN1(n8183), .IN2(n7431), .IN3(n7430), .IN4(n7429), .QN(
        n7432) );
  NOR4X0 U9244 ( .IN1(n7435), .IN2(n7434), .IN3(n7433), .IN4(n7432), .QN(n7441) );
  NAND2X0 U9245 ( .IN1(n7437), .IN2(n7436), .QN(n7440) );
  NAND2X0 U9246 ( .IN1(n9184), .IN2(n7438), .QN(n7439) );
  NAND4X0 U9247 ( .IN1(n7442), .IN2(n7441), .IN3(n7440), .IN4(n7439), .QN(
        \a2/N435 ) );
  OA221X1 U9248 ( .IN1(n9442), .IN2(n7445), .IN3(n9442), .IN4(n7444), .IN5(
        n7443), .Q(n7461) );
  NAND2X0 U9249 ( .IN1(n7984), .IN2(n8724), .QN(n7448) );
  NAND2X0 U9250 ( .IN1(n9125), .IN2(n8640), .QN(n7447) );
  NAND3X0 U9251 ( .IN1(n7448), .IN2(n7447), .IN3(n7446), .QN(n7456) );
  NAND4X0 U9252 ( .IN1(n7450), .IN2(n7861), .IN3(n7498), .IN4(n7449), .QN(
        n7455) );
  NAND2X0 U9253 ( .IN1(n8731), .IN2(n7451), .QN(n7452) );
  NAND4X0 U9254 ( .IN1(n7965), .IN2(n7453), .IN3(n8172), .IN4(n7452), .QN(
        n7454) );
  NOR4X0 U9255 ( .IN1(n7457), .IN2(n7456), .IN3(n7455), .IN4(n7454), .QN(n7460) );
  NAND4X0 U9256 ( .IN1(n7461), .IN2(n7460), .IN3(n7459), .IN4(n7458), .QN(
        \a2/N436 ) );
  NOR2X0 U9257 ( .IN1(n7463), .IN2(n7462), .QN(n7470) );
  NAND2X0 U9258 ( .IN1(n8171), .IN2(n8630), .QN(n7464) );
  OA22X1 U9259 ( .IN1(n7467), .IN2(n7466), .IN3(n7465), .IN4(n7464), .Q(n7468)
         );
  NAND2X0 U9260 ( .IN1(n8551), .IN2(n7468), .QN(n7469) );
  NOR2X0 U9261 ( .IN1(n7470), .IN2(n7469), .QN(n7482) );
  NOR2X0 U9262 ( .IN1(n9445), .IN2(n7471), .QN(n7479) );
  NOR2X0 U9263 ( .IN1(n7473), .IN2(n7472), .QN(n7478) );
  NAND4X0 U9264 ( .IN1(n8835), .IN2(n7475), .IN3(n7845), .IN4(n7474), .QN(
        n7476) );
  NOR4X0 U9265 ( .IN1(n7479), .IN2(n7478), .IN3(n7477), .IN4(n7476), .QN(n7481) );
  NAND4X0 U9266 ( .IN1(n7482), .IN2(n7481), .IN3(n8183), .IN4(n7480), .QN(
        \a2/N437 ) );
  INVX0 U9267 ( .INP(n7483), .ZN(n7709) );
  OA22X1 U9268 ( .IN1(n9084), .IN2(n7709), .IN3(n8041), .IN4(n8851), .Q(n7497)
         );
  NOR2X0 U9269 ( .IN1(n8772), .IN2(n8138), .QN(n7493) );
  NAND2X0 U9270 ( .IN1(n7484), .IN2(n8947), .QN(n7591) );
  NAND4X0 U9271 ( .IN1(n7485), .IN2(n7738), .IN3(n8003), .IN4(n7591), .QN(
        n7491) );
  NOR2X0 U9272 ( .IN1(n7487), .IN2(n7486), .QN(n7489) );
  NAND3X0 U9273 ( .IN1(n8468), .IN2(n9442), .IN3(n9001), .QN(n7488) );
  NAND3X0 U9274 ( .IN1(n7489), .IN2(n8056), .IN3(n7488), .QN(n7490) );
  NOR4X0 U9275 ( .IN1(n7493), .IN2(n7492), .IN3(n7491), .IN4(n7490), .QN(n7496) );
  NAND4X0 U9276 ( .IN1(n7497), .IN2(n7496), .IN3(n7495), .IN4(n7494), .QN(
        \a2/N438 ) );
  NAND2X0 U9277 ( .IN1(n7499), .IN2(n7498), .QN(n7505) );
  NOR2X0 U9278 ( .IN1(n7501), .IN2(n7500), .QN(n8057) );
  OA22X1 U9279 ( .IN1(n8471), .IN2(n9436), .IN3(n8057), .IN4(n8041), .Q(n7502)
         );
  NAND4X0 U9280 ( .IN1(n7503), .IN2(n7502), .IN3(n8922), .IN4(n8541), .QN(
        n7504) );
  NOR4X0 U9281 ( .IN1(n7507), .IN2(n7506), .IN3(n7505), .IN4(n7504), .QN(n7508) );
  OA221X1 U9282 ( .IN1(n8188), .IN2(n7510), .IN3(n8188), .IN4(n7509), .IN5(
        n7508), .Q(n7514) );
  NOR2X0 U9283 ( .IN1(n8474), .IN2(n9166), .QN(n7512) );
  NAND2X0 U9284 ( .IN1(n8153), .IN2(n9083), .QN(n7511) );
  NAND2X0 U9285 ( .IN1(n7512), .IN2(n7511), .QN(n7513) );
  NAND4X0 U9286 ( .IN1(n7514), .IN2(n8524), .IN3(n8765), .IN4(n7513), .QN(
        \a2/N439 ) );
  NAND2X0 U9287 ( .IN1(n8220), .IN2(n7515), .QN(n7516) );
  OA22X1 U9288 ( .IN1(n7517), .IN2(n8104), .IN3(n7516), .IN4(n7736), .Q(n7532)
         );
  NOR2X0 U9289 ( .IN1(n7518), .IN2(n7850), .QN(n7527) );
  INVX0 U9290 ( .INP(n7519), .ZN(n8623) );
  INVX0 U9291 ( .INP(n7520), .ZN(n7790) );
  NAND2X0 U9292 ( .IN1(n8699), .IN2(n7521), .QN(n8251) );
  NAND4X0 U9293 ( .IN1(n7790), .IN2(n8891), .IN3(n8477), .IN4(n8251), .QN(
        n7525) );
  AO22X1 U9294 ( .IN1(n8995), .IN2(n7523), .IN3(n9082), .IN4(n7522), .Q(n7524)
         );
  NOR4X0 U9295 ( .IN1(n8623), .IN2(n8637), .IN3(n7525), .IN4(n7524), .QN(n7526) );
  OA21X1 U9296 ( .IN1(n7527), .IN2(n8692), .IN3(n7526), .Q(n7531) );
  NAND2X0 U9297 ( .IN1(n7529), .IN2(n7528), .QN(n7530) );
  NAND4X0 U9298 ( .IN1(n7532), .IN2(n7531), .IN3(n7558), .IN4(n7530), .QN(
        \a2/N441 ) );
  OA22X1 U9299 ( .IN1(n8461), .IN2(n7533), .IN3(n7766), .IN4(n8041), .Q(n7546)
         );
  NOR2X0 U9300 ( .IN1(n7534), .IN2(n8123), .QN(n7537) );
  NAND3X0 U9301 ( .IN1(n8461), .IN2(n8180), .IN3(n9046), .QN(n7535) );
  NAND2X0 U9302 ( .IN1(n7535), .IN2(n7854), .QN(n7536) );
  NOR2X0 U9303 ( .IN1(n7537), .IN2(n7536), .QN(n7545) );
  NOR2X0 U9304 ( .IN1(n8728), .IN2(n7538), .QN(n7540) );
  NOR2X0 U9305 ( .IN1(n7571), .IN2(n8937), .QN(n7539) );
  NOR4X0 U9306 ( .IN1(n7541), .IN2(n7540), .IN3(n8637), .IN4(n7539), .QN(n7542) );
  OA21X1 U9307 ( .IN1(n9435), .IN2(n7543), .IN3(n7542), .Q(n7544) );
  NAND4X0 U9308 ( .IN1(n7546), .IN2(n7545), .IN3(n7544), .IN4(n7922), .QN(
        \a2/N442 ) );
  OA22X1 U9309 ( .IN1(n9181), .IN2(n8444), .IN3(n7547), .IN4(n9029), .Q(n7565)
         );
  NOR2X0 U9310 ( .IN1(n9435), .IN2(n7548), .QN(n7562) );
  INVX0 U9311 ( .INP(n9117), .ZN(n7985) );
  NOR2X0 U9312 ( .IN1(n9436), .IN2(n7985), .QN(n8920) );
  INVX0 U9313 ( .INP(n8181), .ZN(n7549) );
  OA22X1 U9314 ( .IN1(n9084), .IN2(n7551), .IN3(n7550), .IN4(n7549), .Q(n7559)
         );
  NOR2X0 U9315 ( .IN1(n9080), .IN2(n7552), .QN(n7556) );
  NAND2X0 U9316 ( .IN1(n7554), .IN2(n7553), .QN(n7555) );
  NAND2X0 U9317 ( .IN1(n7556), .IN2(n7555), .QN(n7557) );
  NAND4X0 U9318 ( .IN1(n7559), .IN2(n7558), .IN3(n8487), .IN4(n7557), .QN(
        n7560) );
  NOR4X0 U9319 ( .IN1(n7562), .IN2(n7561), .IN3(n8920), .IN4(n7560), .QN(n7564) );
  NAND4X0 U9320 ( .IN1(n7565), .IN2(n7564), .IN3(n7563), .IN4(n8733), .QN(
        \a2/N443 ) );
  OA22X1 U9321 ( .IN1(n9208), .IN2(n8751), .IN3(n8639), .IN4(n7566), .Q(n7580)
         );
  NOR2X0 U9322 ( .IN1(n9001), .IN2(n8684), .QN(n7570) );
  NAND2X0 U9323 ( .IN1(n7568), .IN2(n7567), .QN(n7569) );
  NOR2X0 U9324 ( .IN1(n7570), .IN2(n7569), .QN(n7579) );
  AND2X1 U9325 ( .IN1(n9060), .IN2(n8475), .Q(n7576) );
  INVX0 U9326 ( .INP(n8086), .ZN(n8984) );
  NOR2X0 U9327 ( .IN1(n8984), .IN2(n8977), .QN(n7575) );
  NOR2X0 U9328 ( .IN1(n7650), .IN2(n7714), .QN(n7574) );
  NOR2X0 U9329 ( .IN1(n7572), .IN2(n7571), .QN(n7573) );
  NOR4X0 U9330 ( .IN1(n7576), .IN2(n7575), .IN3(n7574), .IN4(n7573), .QN(n7578) );
  NAND4X0 U9331 ( .IN1(n7580), .IN2(n7579), .IN3(n7578), .IN4(n7577), .QN(
        \a2/N444 ) );
  OA21X1 U9332 ( .IN1(n8862), .IN2(n8698), .IN3(n8188), .Q(n7595) );
  OA21X1 U9333 ( .IN1(n9005), .IN2(n7581), .IN3(n8752), .Q(n7594) );
  NAND2X0 U9334 ( .IN1(n9031), .IN2(n7582), .QN(n7584) );
  NAND4X0 U9335 ( .IN1(n7585), .IN2(n7845), .IN3(n7584), .IN4(n7583), .QN(
        n7593) );
  INVX0 U9336 ( .INP(n7586), .ZN(n8777) );
  AO21X1 U9337 ( .IN1(n7588), .IN2(n7587), .IN3(n8598), .Q(n7590) );
  NAND2X0 U9338 ( .IN1(n8223), .IN2(n7589), .QN(n9146) );
  NAND4X0 U9339 ( .IN1(n8777), .IN2(n7591), .IN3(n7590), .IN4(n9146), .QN(
        n7592) );
  OR4X1 U9340 ( .IN1(n7595), .IN2(n7594), .IN3(n7593), .IN4(n7592), .Q(
        \a2/N445 ) );
  INVX0 U9341 ( .INP(n7596), .ZN(n7957) );
  AOI22X1 U9342 ( .IN1(n8816), .IN2(n8305), .IN3(n9209), .IN4(n7957), .QN(
        n7610) );
  NAND3X0 U9343 ( .IN1(n9190), .IN2(n9436), .IN3(n7597), .QN(n7598) );
  NAND4X0 U9344 ( .IN1(n7829), .IN2(n7599), .IN3(n8265), .IN4(n7598), .QN(
        n7607) );
  NAND2X0 U9345 ( .IN1(n8889), .IN2(n7600), .QN(n7601) );
  NAND3X0 U9346 ( .IN1(n7601), .IN2(n8474), .IN3(n8890), .QN(n7602) );
  NAND4X0 U9347 ( .IN1(n7605), .IN2(n7604), .IN3(n7603), .IN4(n7602), .QN(
        n7606) );
  NOR2X0 U9348 ( .IN1(n7607), .IN2(n7606), .QN(n7609) );
  INVX0 U9349 ( .INP(n8638), .ZN(n8437) );
  NAND4X0 U9350 ( .IN1(n7610), .IN2(n7609), .IN3(n8437), .IN4(n7608), .QN(
        \a2/N446 ) );
  NAND2X0 U9351 ( .IN1(n7611), .IN2(n9438), .QN(n8864) );
  AND3X1 U9352 ( .IN1(n8055), .IN2(n7612), .IN3(n8864), .Q(n7623) );
  NOR2X0 U9353 ( .IN1(n7613), .IN2(n7736), .QN(n7614) );
  OA21X1 U9354 ( .IN1(n7615), .IN2(n7614), .IN3(n8223), .Q(n7620) );
  NAND3X0 U9355 ( .IN1(n7657), .IN2(n8840), .IN3(n7616), .QN(n7617) );
  AO22X1 U9356 ( .IN1(degrees_tmp2[0]), .IN2(n7618), .IN3(n8692), .IN4(n7617), 
        .Q(n7619) );
  NOR4X0 U9357 ( .IN1(n9176), .IN2(n7621), .IN3(n7620), .IN4(n7619), .QN(n7622) );
  NAND4X0 U9358 ( .IN1(n7623), .IN2(n7622), .IN3(n7709), .IN4(n9146), .QN(
        \a2/N447 ) );
  INVX0 U9359 ( .INP(n7854), .ZN(n7631) );
  NAND2X0 U9360 ( .IN1(n7699), .IN2(n7624), .QN(n7628) );
  AO21X1 U9361 ( .IN1(n8294), .IN2(n8410), .IN3(n8533), .Q(n7627) );
  NAND3X0 U9362 ( .IN1(n9100), .IN2(n8203), .IN3(n8261), .QN(n7625) );
  NAND2X0 U9363 ( .IN1(n7625), .IN2(n8816), .QN(n7626) );
  NAND4X0 U9364 ( .IN1(n8857), .IN2(n7628), .IN3(n7627), .IN4(n7626), .QN(
        n7629) );
  NOR4X0 U9365 ( .IN1(n7632), .IN2(n7631), .IN3(n7630), .IN4(n7629), .QN(n7634) );
  NAND4X0 U9366 ( .IN1(n7634), .IN2(n7856), .IN3(n7633), .IN4(n7820), .QN(
        \a2/N448 ) );
  NAND4X0 U9367 ( .IN1(n7637), .IN2(n7636), .IN3(n7635), .IN4(n8641), .QN(
        n7644) );
  NOR2X0 U9368 ( .IN1(n8754), .IN2(n7638), .QN(n7639) );
  NOR4X0 U9369 ( .IN1(n8496), .IN2(n7640), .IN3(n7788), .IN4(n7639), .QN(n7642) );
  NAND4X0 U9370 ( .IN1(n7642), .IN2(n8554), .IN3(n8878), .IN4(n7641), .QN(
        n7643) );
  NOR2X0 U9371 ( .IN1(n7644), .IN2(n7643), .QN(n7648) );
  NAND2X0 U9372 ( .IN1(n8727), .IN2(n7645), .QN(n7646) );
  NAND4X0 U9373 ( .IN1(n7648), .IN2(n7647), .IN3(n8803), .IN4(n7646), .QN(
        \a2/N449 ) );
  NOR2X0 U9374 ( .IN1(n8423), .IN2(n8026), .QN(n9008) );
  NOR2X0 U9375 ( .IN1(n7650), .IN2(n7649), .QN(n8337) );
  NOR4X0 U9376 ( .IN1(n7652), .IN2(n9008), .IN3(n8337), .IN4(n7651), .QN(n7665) );
  INVX0 U9377 ( .INP(n8823), .ZN(n9052) );
  NOR2X0 U9378 ( .IN1(n7654), .IN2(n7653), .QN(n8570) );
  OA22X1 U9379 ( .IN1(n7655), .IN2(n9052), .IN3(n8570), .IN4(n8724), .Q(n7664)
         );
  NOR2X0 U9380 ( .IN1(n9079), .IN2(n9107), .QN(n9064) );
  NOR2X0 U9381 ( .IN1(n7656), .IN2(n8384), .QN(n7661) );
  OA22X1 U9382 ( .IN1(n8728), .IN2(n9146), .IN3(n7657), .IN4(n8431), .Q(n7659)
         );
  NAND4X0 U9383 ( .IN1(n7659), .IN2(n8069), .IN3(n8452), .IN4(n7658), .QN(
        n7660) );
  NOR4X0 U9384 ( .IN1(n9013), .IN2(n9064), .IN3(n7661), .IN4(n7660), .QN(n7663) );
  NAND4X0 U9385 ( .IN1(n7665), .IN2(n7664), .IN3(n7663), .IN4(n7662), .QN(
        \a2/N450 ) );
  NAND2X0 U9386 ( .IN1(n9080), .IN2(n7666), .QN(n8449) );
  NAND2X0 U9387 ( .IN1(n8534), .IN2(n8484), .QN(n7667) );
  NAND4X0 U9388 ( .IN1(n9067), .IN2(n8900), .IN3(n8449), .IN4(n7667), .QN(
        n7676) );
  NAND3X0 U9389 ( .IN1(n7730), .IN2(n8100), .IN3(n8797), .QN(n7675) );
  NAND3X0 U9390 ( .IN1(n7669), .IN2(n7668), .IN3(n8073), .QN(n7672) );
  NAND3X0 U9391 ( .IN1(n7670), .IN2(n9433), .IN3(n8004), .QN(n7671) );
  NAND4X0 U9392 ( .IN1(n8664), .IN2(n7673), .IN3(n7672), .IN4(n7671), .QN(
        n7674) );
  OR4X1 U9393 ( .IN1(n7677), .IN2(n7676), .IN3(n7675), .IN4(n7674), .Q(
        \a2/N452 ) );
  NOR2X0 U9394 ( .IN1(n9440), .IN2(n8939), .QN(n8207) );
  AND2X1 U9395 ( .IN1(n8531), .IN2(n7678), .Q(n8932) );
  NOR2X0 U9396 ( .IN1(n7679), .IN2(n8171), .QN(n7680) );
  NOR4X0 U9397 ( .IN1(n8207), .IN2(n7681), .IN3(n8932), .IN4(n7680), .QN(n7696) );
  NOR2X0 U9398 ( .IN1(n8841), .IN2(n8667), .QN(n7684) );
  NAND2X0 U9399 ( .IN1(n8137), .IN2(n7682), .QN(n7683) );
  NOR2X0 U9400 ( .IN1(n7684), .IN2(n7683), .QN(n7695) );
  NOR2X0 U9401 ( .IN1(n7686), .IN2(n7685), .QN(n7691) );
  NAND2X0 U9402 ( .IN1(n7952), .IN2(n9433), .QN(n7689) );
  NAND2X0 U9403 ( .IN1(n9031), .IN2(n9195), .QN(n7688) );
  NAND3X0 U9404 ( .IN1(n7689), .IN2(n7688), .IN3(n7687), .QN(n7690) );
  NOR4X0 U9405 ( .IN1(n7693), .IN2(n7692), .IN3(n7691), .IN4(n7690), .QN(n7694) );
  NAND4X0 U9406 ( .IN1(n7696), .IN2(n7695), .IN3(n7694), .IN4(n7944), .QN(
        \a2/N453 ) );
  NOR2X0 U9407 ( .IN1(n8185), .IN2(n8190), .QN(n7697) );
  OA21X1 U9408 ( .IN1(n7698), .IN2(n7697), .IN3(n8728), .Q(n7713) );
  AOI22X1 U9409 ( .IN1(n9082), .IN2(n7701), .IN3(n7700), .IN4(n7699), .QN(
        n7711) );
  INVX0 U9410 ( .INP(n7915), .ZN(n7702) );
  AND3X1 U9411 ( .IN1(n8349), .IN2(n9140), .IN3(n7702), .Q(n7705) );
  NOR2X0 U9412 ( .IN1(n7870), .IN2(n7703), .QN(n7704) );
  OA22X1 U9413 ( .IN1(n7705), .IN2(n8724), .IN3(n7704), .IN4(n9122), .Q(n7710)
         );
  NAND3X0 U9414 ( .IN1(n8301), .IN2(n7707), .IN3(n7706), .QN(n7708) );
  NAND4X0 U9415 ( .IN1(n7711), .IN2(n7710), .IN3(n7709), .IN4(n7708), .QN(
        n7712) );
  OR4X1 U9416 ( .IN1(n8207), .IN2(n9154), .IN3(n7713), .IN4(n7712), .Q(
        \a2/N454 ) );
  OA22X1 U9417 ( .IN1(n8667), .IN2(n7714), .IN3(n8760), .IN4(n9146), .Q(n7732)
         );
  NAND4X0 U9418 ( .IN1(n7716), .IN2(n8905), .IN3(n7715), .IN4(n8367), .QN(
        n7726) );
  OA22X1 U9419 ( .IN1(n8727), .IN2(n7718), .IN3(n7717), .IN4(n8597), .Q(n7724)
         );
  NOR2X0 U9420 ( .IN1(n9023), .IN2(n8914), .QN(n7720) );
  NOR2X0 U9421 ( .IN1(n7720), .IN2(n7719), .QN(n7723) );
  NAND4X0 U9422 ( .IN1(n7724), .IN2(n7723), .IN3(n7722), .IN4(n7721), .QN(
        n7725) );
  NOR4X0 U9423 ( .IN1(n7728), .IN2(n7727), .IN3(n7726), .IN4(n7725), .QN(n7731) );
  NAND4X0 U9424 ( .IN1(n7732), .IN2(n7731), .IN3(n7730), .IN4(n7729), .QN(
        \a2/N455 ) );
  NOR2X0 U9425 ( .IN1(n8444), .IN2(n8332), .QN(n7742) );
  NAND2X0 U9426 ( .IN1(n8529), .IN2(n9019), .QN(n7733) );
  NAND4X0 U9427 ( .IN1(n7873), .IN2(n8613), .IN3(n7734), .IN4(n7733), .QN(
        n7741) );
  AO22X1 U9428 ( .IN1(n7735), .IN2(n9001), .IN3(n8354), .IN4(n8955), .Q(n7740)
         );
  NAND3X0 U9429 ( .IN1(n8163), .IN2(n7736), .IN3(n7913), .QN(n7737) );
  NAND4X0 U9430 ( .IN1(n8406), .IN2(n7738), .IN3(n8265), .IN4(n7737), .QN(
        n7739) );
  NOR4X0 U9431 ( .IN1(n7742), .IN2(n7741), .IN3(n7740), .IN4(n7739), .QN(n7744) );
  NAND4X0 U9432 ( .IN1(n7744), .IN2(n7743), .IN3(n9139), .IN4(n8775), .QN(
        \a2/N456 ) );
  NOR2X0 U9433 ( .IN1(n7746), .IN2(n7745), .QN(n8482) );
  NAND4X0 U9434 ( .IN1(n8452), .IN2(n7747), .IN3(n8926), .IN4(n8504), .QN(
        n7758) );
  INVX0 U9435 ( .INP(n7748), .ZN(n7752) );
  NOR2X0 U9436 ( .IN1(n8724), .IN2(n7749), .QN(n7750) );
  NOR4X0 U9437 ( .IN1(n7752), .IN2(n7751), .IN3(n8344), .IN4(n7750), .QN(n7756) );
  NOR2X0 U9438 ( .IN1(n7754), .IN2(n7753), .QN(n7755) );
  NAND4X0 U9439 ( .IN1(n7756), .IN2(n7755), .IN3(n8882), .IN4(n8454), .QN(
        n7757) );
  NOR4X0 U9440 ( .IN1(n7759), .IN2(n8482), .IN3(n7758), .IN4(n7757), .QN(n7765) );
  NAND2X0 U9441 ( .IN1(n7761), .IN2(n7760), .QN(n7762) );
  NAND4X0 U9442 ( .IN1(n7765), .IN2(n7764), .IN3(n7763), .IN4(n7762), .QN(
        \a2/N457 ) );
  INVX0 U9443 ( .INP(n7766), .ZN(n7768) );
  NAND2X0 U9444 ( .IN1(n7767), .IN2(n8609), .QN(n8089) );
  OA21X1 U9445 ( .IN1(n7768), .IN2(n8089), .IN3(n9442), .Q(n7779) );
  NAND4X0 U9446 ( .IN1(n9030), .IN2(n7771), .IN3(n7770), .IN4(n7769), .QN(
        n7778) );
  NAND3X0 U9447 ( .IN1(n8180), .IN2(n9031), .IN3(n8787), .QN(n7772) );
  NAND4X0 U9448 ( .IN1(n7922), .IN2(n8219), .IN3(n8172), .IN4(n7772), .QN(
        n7777) );
  INVX0 U9449 ( .INP(n7773), .ZN(n7774) );
  AO22X1 U9450 ( .IN1(n8531), .IN2(n7775), .IN3(n9435), .IN4(n7774), .Q(n7776)
         );
  NOR4X0 U9451 ( .IN1(n7779), .IN2(n7778), .IN3(n7777), .IN4(n7776), .QN(n7783) );
  OR2X1 U9452 ( .IN1(n8333), .IN2(n9205), .Q(n7780) );
  NAND4X0 U9453 ( .IN1(n7783), .IN2(n7782), .IN3(n7781), .IN4(n7780), .QN(
        \a2/N458 ) );
  OA22X1 U9454 ( .IN1(n7784), .IN2(n9212), .IN3(n9132), .IN4(n9168), .Q(n7799)
         );
  NOR2X0 U9455 ( .IN1(n9437), .IN2(n8114), .QN(n7796) );
  NAND4X0 U9456 ( .IN1(n7787), .IN2(n7786), .IN3(n7785), .IN4(n8807), .QN(
        n7794) );
  INVX0 U9457 ( .INP(n7788), .ZN(n8577) );
  AND4X1 U9458 ( .IN1(n8625), .IN2(n7790), .IN3(n7789), .IN4(n8577), .Q(n7792)
         );
  NAND4X0 U9459 ( .IN1(n7792), .IN2(n8099), .IN3(n8366), .IN4(n7791), .QN(
        n7793) );
  NOR4X0 U9460 ( .IN1(n7796), .IN2(n7795), .IN3(n7794), .IN4(n7793), .QN(n7798) );
  NAND3X0 U9461 ( .IN1(n7799), .IN2(n7798), .IN3(n7797), .QN(\a2/N459 ) );
  NOR2X0 U9462 ( .IN1(n9445), .IN2(n9041), .QN(n8085) );
  NOR2X0 U9463 ( .IN1(n8085), .IN2(n7849), .QN(n7803) );
  NAND2X0 U9464 ( .IN1(n7801), .IN2(n7800), .QN(n7802) );
  NAND2X0 U9465 ( .IN1(n7803), .IN2(n7802), .QN(n7815) );
  INVX0 U9466 ( .INP(n7804), .ZN(n8499) );
  NOR2X0 U9467 ( .IN1(n7806), .IN2(n7805), .QN(n7807) );
  OA22X1 U9468 ( .IN1(n9435), .IN2(n8499), .IN3(n7807), .IN4(n8595), .Q(n7813)
         );
  NAND2X0 U9469 ( .IN1(n7809), .IN2(n7808), .QN(n7810) );
  NAND4X0 U9470 ( .IN1(n7813), .IN2(n7812), .IN3(n7811), .IN4(n7810), .QN(
        n7814) );
  NOR4X0 U9471 ( .IN1(n7816), .IN2(n7997), .IN3(n7815), .IN4(n7814), .QN(n7819) );
  NAND4X0 U9472 ( .IN1(n7819), .IN2(n7818), .IN3(n7817), .IN4(n8136), .QN(
        \a2/N460 ) );
  OA21X1 U9473 ( .IN1(n7821), .IN2(n8692), .IN3(n7820), .Q(n7836) );
  OA21X1 U9474 ( .IN1(n8667), .IN2(n7822), .IN3(n7890), .Q(n7831) );
  NAND4X0 U9475 ( .IN1(n7824), .IN2(n7823), .IN3(n8054), .IN4(n8251), .QN(
        n7825) );
  NOR4X0 U9476 ( .IN1(n8272), .IN2(n7827), .IN3(n7826), .IN4(n7825), .QN(n7830) );
  AND4X1 U9477 ( .IN1(n7831), .IN2(n7830), .IN3(n7829), .IN4(n7828), .Q(n7835)
         );
  NAND2X0 U9478 ( .IN1(n7832), .IN2(n9023), .QN(n7833) );
  NAND4X0 U9479 ( .IN1(n7836), .IN2(n7835), .IN3(n7834), .IN4(n7833), .QN(
        \a2/N461 ) );
  OA21X1 U9480 ( .IN1(n7838), .IN2(n9433), .IN3(n7837), .Q(n7847) );
  OA22X1 U9481 ( .IN1(n7841), .IN2(n7840), .IN3(n9208), .IN4(n7839), .Q(n7846)
         );
  NAND2X0 U9482 ( .IN1(n7843), .IN2(n7842), .QN(n7844) );
  NAND4X0 U9483 ( .IN1(n7847), .IN2(n7846), .IN3(n7845), .IN4(n7844), .QN(
        n7848) );
  NOR4X0 U9484 ( .IN1(n7850), .IN2(n7849), .IN3(n8111), .IN4(n7848), .QN(n7852) );
  NAND2X0 U9485 ( .IN1(n9195), .IN2(n9001), .QN(n8353) );
  NAND4X0 U9486 ( .IN1(n7853), .IN2(n7852), .IN3(n7851), .IN4(n8353), .QN(
        \a2/N462 ) );
  NAND4X0 U9487 ( .IN1(n7857), .IN2(n7856), .IN3(n7855), .IN4(n7854), .QN(
        n7868) );
  NAND2X0 U9488 ( .IN1(n7858), .IN2(n8511), .QN(n7859) );
  NAND4X0 U9489 ( .IN1(n7862), .IN2(n7861), .IN3(n7860), .IN4(n7859), .QN(
        n7867) );
  NAND2X0 U9490 ( .IN1(n8534), .IN2(n7863), .QN(n7864) );
  NAND4X0 U9491 ( .IN1(n8131), .IN2(n7865), .IN3(n8850), .IN4(n7864), .QN(
        n7866) );
  NOR4X0 U9492 ( .IN1(n7869), .IN2(n7868), .IN3(n7867), .IN4(n7866), .QN(n7874) );
  NAND2X0 U9493 ( .IN1(n9054), .IN2(n7870), .QN(n7871) );
  NAND4X0 U9494 ( .IN1(n7874), .IN2(n7873), .IN3(n7872), .IN4(n7871), .QN(
        \a2/N463 ) );
  OA22X1 U9495 ( .IN1(n8796), .IN2(n7876), .IN3(n8645), .IN4(n7875), .Q(n7893)
         );
  NOR2X0 U9496 ( .IN1(n9071), .IN2(n8261), .QN(n7888) );
  NAND2X0 U9497 ( .IN1(n8669), .IN2(n9072), .QN(n7877) );
  AO22X1 U9498 ( .IN1(n8534), .IN2(n7879), .IN3(n7878), .IN4(n7877), .Q(n7887)
         );
  NOR2X0 U9499 ( .IN1(n7881), .IN2(n7880), .QN(n7883) );
  INVX0 U9500 ( .INP(n8701), .ZN(n7882) );
  NOR3X0 U9501 ( .IN1(n7883), .IN2(n8482), .IN3(n7882), .QN(n7885) );
  NAND4X0 U9502 ( .IN1(n7885), .IN2(n7991), .IN3(n8487), .IN4(n7884), .QN(
        n7886) );
  NOR4X0 U9503 ( .IN1(n7889), .IN2(n7888), .IN3(n7887), .IN4(n7886), .QN(n7892) );
  NAND4X0 U9504 ( .IN1(n7893), .IN2(n7892), .IN3(n7891), .IN4(n7890), .QN(
        \a2/N464 ) );
  INVX0 U9505 ( .INP(n7894), .ZN(n8738) );
  OA22X1 U9506 ( .IN1(n8847), .IN2(n8738), .IN3(n7895), .IN4(n9020), .Q(n7912)
         );
  AO22X1 U9507 ( .IN1(n7898), .IN2(n7897), .IN3(n7896), .IN4(n8649), .Q(n7906)
         );
  NOR2X0 U9508 ( .IN1(n8185), .IN2(n8841), .QN(n7899) );
  NOR2X0 U9509 ( .IN1(n7900), .IN2(n7899), .QN(n7904) );
  NAND2X0 U9510 ( .IN1(n7902), .IN2(n7901), .QN(n7903) );
  NAND2X0 U9511 ( .IN1(n7904), .IN2(n7903), .QN(n7905) );
  NOR4X0 U9512 ( .IN1(n7908), .IN2(n7907), .IN3(n7906), .IN4(n7905), .QN(n7909) );
  OA21X1 U9513 ( .IN1(degrees_tmp2[0]), .IN2(n7910), .IN3(n7909), .Q(n7911) );
  NAND4X0 U9514 ( .IN1(n7912), .IN2(n7911), .IN3(n7981), .IN4(n8003), .QN(
        \a2/N465 ) );
  NOR2X0 U9515 ( .IN1(n8228), .IN2(n7913), .QN(n7919) );
  AO22X1 U9516 ( .IN1(n8825), .IN2(n7916), .IN3(n7915), .IN4(n7914), .Q(n7917)
         );
  NOR3X0 U9517 ( .IN1(n7919), .IN2(n7918), .IN3(n7917), .QN(n7932) );
  NAND2X0 U9518 ( .IN1(n7921), .IN2(n7920), .QN(n7931) );
  NOR2X0 U9519 ( .IN1(degrees_tmp2[2]), .IN2(n8339), .QN(n7929) );
  AO21X1 U9520 ( .IN1(n8183), .IN2(n8367), .IN3(degrees_tmp2[0]), .Q(n7925) );
  AO21X1 U9521 ( .IN1(n7922), .IN2(n8156), .IN3(n9084), .Q(n7923) );
  NAND4X0 U9522 ( .IN1(n7926), .IN2(n7925), .IN3(n7924), .IN4(n7923), .QN(
        n7927) );
  NOR4X0 U9523 ( .IN1(n7929), .IN2(n7928), .IN3(n8257), .IN4(n7927), .QN(n7930) );
  NAND4X0 U9524 ( .IN1(n7932), .IN2(n8610), .IN3(n7931), .IN4(n7930), .QN(
        \a2/N466 ) );
  NOR2X0 U9525 ( .IN1(n7933), .IN2(n8528), .QN(n8582) );
  NOR4X0 U9526 ( .IN1(n7934), .IN2(n8683), .IN3(n8066), .IN4(n8582), .QN(n7950) );
  NAND2X0 U9527 ( .IN1(n7936), .IN2(n7935), .QN(n7937) );
  NAND4X0 U9528 ( .IN1(n7940), .IN2(n7939), .IN3(n7938), .IN4(n7937), .QN(
        n7941) );
  NOR2X0 U9529 ( .IN1(n8058), .IN2(n7941), .QN(n7942) );
  OA221X1 U9530 ( .IN1(n9435), .IN2(n7944), .IN3(n9435), .IN4(n7943), .IN5(
        n7942), .Q(n7949) );
  NAND4X0 U9531 ( .IN1(n8186), .IN2(n9436), .IN3(n7945), .IN4(n8026), .QN(
        n7948) );
  NAND2X0 U9532 ( .IN1(n7946), .IN2(n8938), .QN(n7947) );
  NAND4X0 U9533 ( .IN1(n7950), .IN2(n7949), .IN3(n7948), .IN4(n7947), .QN(
        \a2/N467 ) );
  INVX0 U9534 ( .INP(n7951), .ZN(n7963) );
  AO22X1 U9535 ( .IN1(n9435), .IN2(n7952), .IN3(n7973), .IN4(n8822), .Q(n7962)
         );
  AND2X1 U9536 ( .IN1(n7954), .IN2(n7953), .Q(n7955) );
  OA22X1 U9537 ( .IN1(n7955), .IN2(n8073), .IN3(n8171), .IN4(n8705), .Q(n7959)
         );
  NAND3X0 U9538 ( .IN1(degrees_tmp2[2]), .IN2(n7957), .IN3(n7956), .QN(n7958)
         );
  NAND4X0 U9539 ( .IN1(n7960), .IN2(n7959), .IN3(n8056), .IN4(n7958), .QN(
        n7961) );
  NOR4X0 U9540 ( .IN1(n7964), .IN2(n7963), .IN3(n7962), .IN4(n7961), .QN(n7966) );
  NAND4X0 U9541 ( .IN1(n7967), .IN2(n7966), .IN3(n8776), .IN4(n7965), .QN(
        \a2/N468 ) );
  INVX0 U9542 ( .INP(n7968), .ZN(n7980) );
  NOR2X0 U9543 ( .IN1(n8139), .IN2(n7969), .QN(n7979) );
  AO22X1 U9544 ( .IN1(n7971), .IN2(n8710), .IN3(n7970), .IN4(n8004), .Q(n7978)
         );
  INVX0 U9545 ( .INP(n7972), .ZN(n7976) );
  NAND2X0 U9546 ( .IN1(n8890), .IN2(n7973), .QN(n7974) );
  NAND4X0 U9547 ( .IN1(n8193), .IN2(n7976), .IN3(n7975), .IN4(n7974), .QN(
        n7977) );
  NOR4X0 U9548 ( .IN1(n7980), .IN2(n7979), .IN3(n7978), .IN4(n7977), .QN(n7982) );
  NAND4X0 U9549 ( .IN1(n7983), .IN2(n7982), .IN3(n7981), .IN4(n8845), .QN(
        \a2/N469 ) );
  NOR2X0 U9550 ( .IN1(n7984), .IN2(n8429), .QN(n9081) );
  NAND4X0 U9551 ( .IN1(n9081), .IN2(n8029), .IN3(n8448), .IN4(n8248), .QN(
        n7996) );
  OA21X1 U9552 ( .IN1(n8728), .IN2(n8882), .IN3(n7985), .Q(n8313) );
  NAND4X0 U9553 ( .IN1(n8313), .IN2(n8437), .IN3(n7987), .IN4(n7986), .QN(
        n7995) );
  OA22X1 U9554 ( .IN1(n8122), .IN2(n7989), .IN3(n9445), .IN4(n7988), .Q(n7993)
         );
  NAND4X0 U9555 ( .IN1(n7993), .IN2(n7992), .IN3(n7991), .IN4(n7990), .QN(
        n7994) );
  OR4X1 U9556 ( .IN1(n7997), .IN2(n7996), .IN3(n7995), .IN4(n7994), .Q(
        \a2/N470 ) );
  INVX0 U9557 ( .INP(n7998), .ZN(n8019) );
  OA221X1 U9558 ( .IN1(n9124), .IN2(n8000), .IN3(n9124), .IN4(n7999), .IN5(
        n9445), .Q(n8018) );
  NOR2X0 U9559 ( .IN1(n8922), .IN2(n8001), .QN(n8015) );
  OR2X1 U9560 ( .IN1(n8592), .IN2(n8511), .Q(n8002) );
  NAND4X0 U9561 ( .IN1(n8226), .IN2(n8003), .IN3(n8263), .IN4(n8002), .QN(
        n8014) );
  AOI22X1 U9562 ( .IN1(degrees_tmp2[5]), .IN2(n8006), .IN3(n8005), .IN4(n8004), 
        .QN(n8010) );
  NAND2X0 U9563 ( .IN1(n8624), .IN2(n8007), .QN(n8008) );
  NAND2X0 U9564 ( .IN1(n8171), .IN2(n8008), .QN(n8009) );
  NAND4X0 U9565 ( .IN1(n8012), .IN2(n8011), .IN3(n8010), .IN4(n8009), .QN(
        n8013) );
  OR4X1 U9566 ( .IN1(n8016), .IN2(n8015), .IN3(n8014), .IN4(n8013), .Q(n8017)
         );
  AO221X1 U9567 ( .IN1(n9435), .IN2(n8019), .IN3(n9435), .IN4(n8018), .IN5(
        n8017), .Q(\a2/N471 ) );
  OA22X1 U9568 ( .IN1(n8022), .IN2(n8021), .IN3(degrees_tmp2[0]), .IN4(n8020), 
        .Q(n8036) );
  INVX0 U9569 ( .INP(n8023), .ZN(n8032) );
  NAND4X0 U9570 ( .IN1(n8025), .IN2(n8689), .IN3(n8024), .IN4(n8367), .QN(
        n8031) );
  NAND2X0 U9571 ( .IN1(n8186), .IN2(n8026), .QN(n8027) );
  NAND4X0 U9572 ( .IN1(n8624), .IN2(n8029), .IN3(n8028), .IN4(n8027), .QN(
        n8030) );
  NOR4X0 U9573 ( .IN1(n8786), .IN2(n8032), .IN3(n8031), .IN4(n8030), .QN(n8035) );
  NAND2X0 U9574 ( .IN1(n8034), .IN2(n8033), .QN(n8325) );
  NAND4X0 U9575 ( .IN1(n8037), .IN2(n8036), .IN3(n8035), .IN4(n8325), .QN(
        \a2/N472 ) );
  OA21X1 U9576 ( .IN1(n8494), .IN2(n8979), .IN3(n8038), .Q(n8051) );
  OAI221X1 U9577 ( .IN1(n8041), .IN2(n8040), .IN3(n8041), .IN4(n8039), .IN5(
        n8060), .QN(n8047) );
  NAND4X0 U9578 ( .IN1(n8043), .IN2(n8042), .IN3(n8609), .IN4(n8732), .QN(
        n8046) );
  OAI22X1 U9579 ( .IN1(n9054), .IN2(n8044), .IN3(n9082), .IN4(n8779), .QN(
        n8045) );
  NOR4X0 U9580 ( .IN1(n8048), .IN2(n8047), .IN3(n8046), .IN4(n8045), .QN(n8050) );
  NAND4X0 U9581 ( .IN1(n8051), .IN2(n8050), .IN3(n8156), .IN4(n8049), .QN(
        \a2/N474 ) );
  NAND2X0 U9582 ( .IN1(n8875), .IN2(n8467), .QN(n8052) );
  NAND4X0 U9583 ( .IN1(n8167), .IN2(n8053), .IN3(n8747), .IN4(n8052), .QN(
        n8065) );
  NAND4X0 U9584 ( .IN1(n8055), .IN2(n8452), .IN3(n8054), .IN4(n8961), .QN(
        n8064) );
  OA21X1 U9585 ( .IN1(n8057), .IN2(n9122), .IN3(n8056), .Q(n8062) );
  INVX0 U9586 ( .INP(n8058), .ZN(n8061) );
  NAND4X0 U9587 ( .IN1(n8062), .IN2(n8061), .IN3(n8060), .IN4(n8059), .QN(
        n8063) );
  OR4X1 U9588 ( .IN1(n8066), .IN2(n8065), .IN3(n8064), .IN4(n8063), .Q(
        \a2/N475 ) );
  AND3X1 U9589 ( .IN1(n8067), .IN2(n8817), .IN3(n8941), .Q(n8080) );
  NAND4X0 U9590 ( .IN1(n8070), .IN2(n8069), .IN3(n8068), .IN4(n8838), .QN(
        n8076) );
  NAND2X0 U9591 ( .IN1(n8071), .IN2(n8977), .QN(n8072) );
  AO22X1 U9592 ( .IN1(n8074), .IN2(n8531), .IN3(n8073), .IN4(n8072), .Q(n8075)
         );
  NOR4X0 U9593 ( .IN1(n8078), .IN2(n8077), .IN3(n8076), .IN4(n8075), .QN(n8079) );
  NAND4X0 U9594 ( .IN1(n8082), .IN2(n8081), .IN3(n8080), .IN4(n8079), .QN(
        \a2/N476 ) );
  OA22X1 U9595 ( .IN1(n8883), .IN2(n8748), .IN3(n8859), .IN4(n8083), .Q(n8096)
         );
  NOR2X0 U9596 ( .IN1(n8249), .IN2(n8084), .QN(n8093) );
  NOR2X0 U9597 ( .IN1(n9013), .IN2(n8085), .QN(n8088) );
  NAND2X0 U9598 ( .IN1(n8731), .IN2(n8086), .QN(n8087) );
  NAND2X0 U9599 ( .IN1(n8088), .IN2(n8087), .QN(n8092) );
  NOR2X0 U9600 ( .IN1(n8742), .IN2(n8089), .QN(n8090) );
  NAND4X0 U9601 ( .IN1(n8090), .IN2(n8200), .IN3(n8913), .IN4(n9126), .QN(
        n8091) );
  NOR4X0 U9602 ( .IN1(n8094), .IN2(n8093), .IN3(n8092), .IN4(n8091), .QN(n8095) );
  NAND2X0 U9603 ( .IN1(n8898), .IN2(n8240), .QN(n8798) );
  NAND4X0 U9604 ( .IN1(n8096), .IN2(n8095), .IN3(n8522), .IN4(n8798), .QN(
        \a2/N477 ) );
  OA21X1 U9605 ( .IN1(n8097), .IN2(n9176), .IN3(n9436), .Q(n8110) );
  INVX0 U9606 ( .INP(n8098), .ZN(n8498) );
  NAND4X0 U9607 ( .IN1(n8100), .IN2(n8099), .IN3(n8498), .IN4(n8672), .QN(
        n8109) );
  NAND2X0 U9608 ( .IN1(n8188), .IN2(n8101), .QN(n8102) );
  OA22X1 U9609 ( .IN1(n8511), .IN2(n8104), .IN3(n8103), .IN4(n8102), .Q(n8107)
         );
  INVX0 U9610 ( .INP(n8105), .ZN(n8908) );
  NAND4X0 U9611 ( .IN1(n8107), .IN2(n8908), .IN3(n8499), .IN4(n8106), .QN(
        n8108) );
  NOR4X0 U9612 ( .IN1(n8111), .IN2(n8110), .IN3(n8109), .IN4(n8108), .QN(n8115) );
  NAND2X0 U9613 ( .IN1(n8112), .IN2(n9438), .QN(n8113) );
  NAND4X0 U9614 ( .IN1(n8115), .IN2(n8720), .IN3(n8114), .IN4(n8113), .QN(
        \a2/N478 ) );
  OA21X1 U9615 ( .IN1(degrees_tmp2[2]), .IN2(n8117), .IN3(n8116), .Q(n8134) );
  NAND3X0 U9616 ( .IN1(degrees_tmp2[2]), .IN2(n8119), .IN3(n8118), .QN(n8121)
         );
  OA22X1 U9617 ( .IN1(n8630), .IN2(n8591), .IN3(n8121), .IN4(n8120), .Q(n8133)
         );
  NOR2X0 U9618 ( .IN1(n8122), .IN2(n8968), .QN(n8129) );
  OAI22X1 U9619 ( .IN1(n8424), .IN2(n8281), .IN3(n8124), .IN4(n8123), .QN(
        n8128) );
  OAI21X1 U9620 ( .IN1(n8995), .IN2(n8126), .IN3(n8125), .QN(n8127) );
  NOR4X0 U9621 ( .IN1(n8130), .IN2(n8129), .IN3(n8128), .IN4(n8127), .QN(n8132) );
  NAND4X0 U9622 ( .IN1(n8134), .IN2(n8133), .IN3(n8132), .IN4(n8131), .QN(
        \a2/N479 ) );
  OA21X1 U9623 ( .IN1(degrees_tmp2[5]), .IN2(n8136), .IN3(n8135), .Q(n8151) );
  OA21X1 U9624 ( .IN1(n8139), .IN2(n8138), .IN3(n8137), .Q(n8150) );
  NOR2X0 U9625 ( .IN1(n8140), .IN2(n8495), .QN(n8141) );
  NOR4X0 U9626 ( .IN1(n8144), .IN2(n8143), .IN3(n8142), .IN4(n8141), .QN(n8149) );
  NAND2X0 U9627 ( .IN1(n9182), .IN2(n8145), .QN(n8146) );
  AND4X1 U9628 ( .IN1(n8720), .IN2(n8147), .IN3(n8339), .IN4(n8146), .Q(n8148)
         );
  NAND4X0 U9629 ( .IN1(n8151), .IN2(n8150), .IN3(n8149), .IN4(n8148), .QN(
        \a2/N481 ) );
  NAND2X0 U9630 ( .IN1(n8153), .IN2(n8152), .QN(n8154) );
  AO22X1 U9631 ( .IN1(n8155), .IN2(n9438), .IN3(n9166), .IN4(n8154), .Q(n8161)
         );
  NAND3X0 U9632 ( .IN1(n8193), .IN2(n8157), .IN3(n8156), .QN(n8160) );
  NAND4X0 U9633 ( .IN1(n8964), .IN2(n8158), .IN3(n8382), .IN4(n8347), .QN(
        n8159) );
  NOR4X0 U9634 ( .IN1(n8162), .IN2(n8161), .IN3(n8160), .IN4(n8159), .QN(n8166) );
  NAND2X0 U9635 ( .IN1(n8188), .IN2(n8163), .QN(n8165) );
  NAND4X0 U9636 ( .IN1(n8166), .IN2(n8165), .IN3(n8164), .IN4(n8403), .QN(
        \a2/N482 ) );
  NAND2X0 U9637 ( .IN1(n8592), .IN2(n8167), .QN(n8177) );
  OA22X1 U9638 ( .IN1(n8568), .IN2(n8170), .IN3(n8169), .IN4(n8168), .Q(n8174)
         );
  NAND2X0 U9639 ( .IN1(n8640), .IN2(n8171), .QN(n8173) );
  NAND4X0 U9640 ( .IN1(n8175), .IN2(n8174), .IN3(n8173), .IN4(n8172), .QN(
        n8176) );
  NOR4X0 U9641 ( .IN1(n8179), .IN2(n8178), .IN3(n8177), .IN4(n8176), .QN(n8184) );
  NAND2X0 U9642 ( .IN1(n8180), .IN2(n8639), .QN(n8409) );
  NAND2X0 U9643 ( .IN1(n8181), .IN2(n8947), .QN(n8182) );
  NAND4X0 U9644 ( .IN1(n8184), .IN2(n8183), .IN3(n8409), .IN4(n8182), .QN(
        \a2/N483 ) );
  NAND2X0 U9645 ( .IN1(n8186), .IN2(n8185), .QN(n8187) );
  NAND4X0 U9646 ( .IN1(n8349), .IN2(n8187), .IN3(n8477), .IN4(n8504), .QN(
        n8196) );
  NAND2X0 U9647 ( .IN1(n8188), .IN2(n8431), .QN(n8191) );
  OA21X1 U9648 ( .IN1(n8191), .IN2(n8190), .IN3(n8189), .Q(n8194) );
  NAND4X0 U9649 ( .IN1(n8194), .IN2(n8193), .IN3(n9102), .IN4(n8192), .QN(
        n8195) );
  NOR2X0 U9650 ( .IN1(n8196), .IN2(n8195), .QN(n8201) );
  NAND2X0 U9651 ( .IN1(n8198), .IN2(n8197), .QN(n8199) );
  NAND4X0 U9652 ( .IN1(n8201), .IN2(n8602), .IN3(n8200), .IN4(n8199), .QN(
        \a2/N484 ) );
  NAND4X0 U9653 ( .IN1(n8927), .IN2(n8204), .IN3(n8203), .IN4(n8202), .QN(
        n8205) );
  NOR3X0 U9654 ( .IN1(n8207), .IN2(n8206), .IN3(n8205), .QN(n8210) );
  NAND4X0 U9655 ( .IN1(n8211), .IN2(n8210), .IN3(n8209), .IN4(n8208), .QN(
        \a2/N486 ) );
  OA22X1 U9656 ( .IN1(n8699), .IN2(n8268), .IN3(n8213), .IN4(n8212), .Q(n8215)
         );
  NAND3X0 U9657 ( .IN1(n8216), .IN2(n8215), .IN3(n8214), .QN(\a2/N487 ) );
  NAND3X0 U9658 ( .IN1(n8219), .IN2(n8218), .IN3(n8217), .QN(\a2/N488 ) );
  NAND2X0 U9659 ( .IN1(n9212), .IN2(n8422), .QN(n9186) );
  OR2X1 U9660 ( .IN1(n9186), .IN2(n8220), .Q(\a2/N490 ) );
  OA21X1 U9661 ( .IN1(n8220), .IN2(\a3/N492 ), .IN3(quad[1]), .Q(\a1/N491 ) );
  NAND2X0 U9662 ( .IN1(quad[0]), .IN2(quad[1]), .QN(n8221) );
  OA21X1 U9663 ( .IN1(\a1/N491 ), .IN2(\a3/N493 ), .IN3(n8221), .Q(\a2/N491 )
         );
  NAND2X0 U9664 ( .IN1(n8223), .IN2(n8222), .QN(n9056) );
  NAND4X0 U9665 ( .IN1(n8226), .IN2(n8225), .IN3(n8224), .IN4(n9056), .QN(
        n8234) );
  OA22X1 U9666 ( .IN1(n8229), .IN2(n8228), .IN3(n9083), .IN4(n8227), .Q(n8232)
         );
  NAND4X0 U9667 ( .IN1(n8232), .IN2(n8231), .IN3(n8230), .IN4(n8263), .QN(
        n8233) );
  NOR2X0 U9668 ( .IN1(n8234), .IN2(n8233), .QN(n8237) );
  NAND4X0 U9669 ( .IN1(n8238), .IN2(n8237), .IN3(n8236), .IN4(n8235), .QN(
        \a1/N435 ) );
  NAND2X0 U9670 ( .IN1(n8240), .IN2(n8239), .QN(n9151) );
  NAND2X0 U9671 ( .IN1(n8242), .IN2(n8241), .QN(n8243) );
  AND3X1 U9672 ( .IN1(n8244), .IN2(n9151), .IN3(n8243), .Q(n8260) );
  OA22X1 U9673 ( .IN1(n8247), .IN2(n8246), .IN3(n9440), .IN4(n8245), .Q(n8259)
         );
  NOR2X0 U9674 ( .IN1(n8249), .IN2(n8248), .QN(n8255) );
  NAND2X0 U9675 ( .IN1(n9023), .IN2(n9075), .QN(n8250) );
  NAND4X0 U9676 ( .IN1(n8253), .IN2(n8252), .IN3(n8251), .IN4(n8250), .QN(
        n8254) );
  NOR4X0 U9677 ( .IN1(n8257), .IN2(n8256), .IN3(n8255), .IN4(n8254), .QN(n8258) );
  NAND4X0 U9678 ( .IN1(n8260), .IN2(n8259), .IN3(n8258), .IN4(n8913), .QN(
        \a1/N436 ) );
  OA22X1 U9679 ( .IN1(n8978), .IN2(n8262), .IN3(n8984), .IN4(n8261), .Q(n8266)
         );
  NAND4X0 U9680 ( .IN1(n8266), .IN2(n8265), .IN3(n8264), .IN4(n8263), .QN(
        n8271) );
  NAND4X0 U9681 ( .IN1(n8268), .IN2(n8726), .IN3(n8267), .IN4(n8294), .QN(
        n8269) );
  AO22X1 U9682 ( .IN1(n8424), .IN2(n8305), .IN3(n8575), .IN4(n8269), .Q(n8270)
         );
  NOR2X0 U9683 ( .IN1(n8271), .IN2(n8270), .QN(n8275) );
  INVX0 U9684 ( .INP(n8272), .ZN(n8493) );
  NAND2X0 U9685 ( .IN1(n9080), .IN2(n8273), .QN(n8274) );
  NAND4X0 U9686 ( .IN1(n8275), .IN2(n8493), .IN3(n8388), .IN4(n8274), .QN(
        \a1/N437 ) );
  NAND3X0 U9687 ( .IN1(n8276), .IN2(n8445), .IN3(n8960), .QN(n8277) );
  NAND2X0 U9688 ( .IN1(n8277), .IN2(n9031), .QN(n8278) );
  NAND3X0 U9689 ( .IN1(n8280), .IN2(n8279), .IN3(n8278), .QN(n8285) );
  OA22X1 U9690 ( .IN1(n9434), .IN2(n8281), .IN3(n8431), .IN4(n9212), .Q(n8283)
         );
  NAND3X0 U9691 ( .IN1(degrees_tmp2[3]), .IN2(n8468), .IN3(n8282), .QN(n8712)
         );
  NAND4X0 U9692 ( .IN1(n8283), .IN2(n8712), .IN3(n8554), .IN4(n8492), .QN(
        n8284) );
  NOR4X0 U9693 ( .IN1(n8287), .IN2(n8286), .IN3(n8285), .IN4(n8284), .QN(n8293) );
  NAND2X0 U9694 ( .IN1(n8289), .IN2(n8288), .QN(n8290) );
  NAND4X0 U9695 ( .IN1(n8293), .IN2(n8292), .IN3(n8291), .IN4(n8290), .QN(
        \a1/N438 ) );
  NOR2X0 U9696 ( .IN1(n8294), .IN2(n9082), .QN(n8298) );
  NAND2X0 U9697 ( .IN1(n8296), .IN2(n8295), .QN(n8297) );
  NOR2X0 U9698 ( .IN1(n8298), .IN2(n8297), .QN(n8312) );
  NOR2X0 U9699 ( .IN1(n9440), .IN2(n8299), .QN(n8309) );
  OA221X1 U9700 ( .IN1(n8302), .IN2(n8301), .IN3(n8302), .IN4(n8300), .IN5(
        n9189), .Q(n8308) );
  NAND3X0 U9701 ( .IN1(n8707), .IN2(n8304), .IN3(n8303), .QN(n8306) );
  AO22X1 U9702 ( .IN1(n9031), .IN2(n8306), .IN3(n8305), .IN4(n8467), .Q(n8307)
         );
  NOR4X0 U9703 ( .IN1(n8310), .IN2(n8309), .IN3(n8308), .IN4(n8307), .QN(n8311) );
  NAND4X0 U9704 ( .IN1(n8313), .IN2(n8312), .IN3(n8311), .IN4(n8817), .QN(
        \a1/N439 ) );
  AND3X1 U9705 ( .IN1(n8316), .IN2(n8315), .IN3(n8314), .Q(n8318) );
  OA22X1 U9706 ( .IN1(n9071), .IN2(n8318), .IN3(n8317), .IN4(n8904), .Q(n8329)
         );
  OA21X1 U9707 ( .IN1(n8320), .IN2(n8319), .IN3(n9001), .Q(n8323) );
  NOR2X0 U9708 ( .IN1(n8321), .IN2(n8685), .QN(n8322) );
  NOR4X0 U9709 ( .IN1(n8324), .IN2(n8323), .IN3(n8628), .IN4(n8322), .QN(n8328) );
  AO21X1 U9710 ( .IN1(n8326), .IN2(n8325), .IN3(degrees_tmp2[3]), .Q(n8327) );
  NAND4X0 U9711 ( .IN1(n8329), .IN2(n8328), .IN3(n8327), .IN4(n8403), .QN(
        \a1/N440 ) );
  NAND2X0 U9712 ( .IN1(n8330), .IN2(n9099), .QN(n8335) );
  AO21X1 U9713 ( .IN1(n8333), .IN2(n8332), .IN3(n8331), .Q(n8334) );
  NAND4X0 U9714 ( .IN1(n8336), .IN2(n8551), .IN3(n8335), .IN4(n8334), .QN(
        n8342) );
  NAND2X0 U9715 ( .IN1(n8337), .IN2(n9445), .QN(n8340) );
  NAND3X0 U9716 ( .IN1(n8340), .IN2(n8339), .IN3(n8338), .QN(n8341) );
  NOR4X0 U9717 ( .IN1(n8344), .IN2(n8343), .IN3(n8342), .IN4(n8341), .QN(n8348) );
  INVX0 U9718 ( .INP(n9187), .ZN(n8346) );
  NAND2X0 U9719 ( .IN1(n9183), .IN2(n8655), .QN(n8345) );
  NAND4X0 U9720 ( .IN1(n8348), .IN2(n8347), .IN3(n8346), .IN4(n8345), .QN(
        \a1/N441 ) );
  OA21X1 U9721 ( .IN1(n8824), .IN2(n8350), .IN3(n8349), .Q(n8351) );
  OA22X1 U9722 ( .IN1(n8351), .IN2(n8649), .IN3(n8489), .IN4(n8406), .Q(n8362)
         );
  NAND2X0 U9723 ( .IN1(n8352), .IN2(n9032), .QN(n8814) );
  OA22X1 U9724 ( .IN1(n9125), .IN2(n8814), .IN3(degrees_tmp2[2]), .IN4(n8353), 
        .Q(n8361) );
  OA221X1 U9725 ( .IN1(n8898), .IN2(n9037), .IN3(n8898), .IN4(n8354), .IN5(
        n8796), .Q(n8357) );
  NAND2X0 U9726 ( .IN1(n8355), .IN2(n8900), .QN(n8356) );
  NOR4X0 U9727 ( .IN1(n8359), .IN2(n8358), .IN3(n8357), .IN4(n8356), .QN(n8360) );
  NAND4X0 U9728 ( .IN1(n8363), .IN2(n8362), .IN3(n8361), .IN4(n8360), .QN(
        \a1/N442 ) );
  OA22X1 U9729 ( .IN1(n9001), .IN2(n9079), .IN3(n8431), .IN4(n8507), .Q(n8377)
         );
  INVX0 U9730 ( .INP(n8364), .ZN(n8370) );
  NOR2X0 U9731 ( .IN1(n9440), .IN2(n9109), .QN(n9138) );
  INVX0 U9732 ( .INP(n9138), .ZN(n8365) );
  NAND4X0 U9733 ( .IN1(n8564), .IN2(n8367), .IN3(n8366), .IN4(n8365), .QN(
        n8368) );
  NOR4X0 U9734 ( .IN1(n8371), .IN2(n8370), .IN3(n8369), .IN4(n8368), .QN(n8372) );
  OA21X1 U9735 ( .IN1(n8710), .IN2(n8373), .IN3(n8372), .Q(n8376) );
  NAND4X0 U9736 ( .IN1(n8377), .IN2(n8376), .IN3(n8375), .IN4(n8374), .QN(
        \a1/N445 ) );
  NOR2X0 U9737 ( .IN1(n8379), .IN2(n8378), .QN(n8398) );
  INVX0 U9738 ( .INP(n8380), .ZN(n8394) );
  NOR2X0 U9739 ( .IN1(n9440), .IN2(n8381), .QN(n8392) );
  OA22X1 U9740 ( .IN1(n8598), .IN2(n8383), .IN3(n9080), .IN4(n8382), .Q(n8390)
         );
  INVX0 U9741 ( .INP(n8384), .ZN(n8805) );
  NOR2X0 U9742 ( .IN1(n8898), .IN2(n8805), .QN(n8387) );
  OA22X1 U9743 ( .IN1(n8387), .IN2(n8568), .IN3(n8386), .IN4(n8385), .Q(n8389)
         );
  NAND4X0 U9744 ( .IN1(n8390), .IN2(n8389), .IN3(n9098), .IN4(n8388), .QN(
        n8391) );
  NOR4X0 U9745 ( .IN1(n8394), .IN2(n8393), .IN3(n8392), .IN4(n8391), .QN(n8397) );
  NAND2X0 U9746 ( .IN1(degrees_tmp2[5]), .IN2(n8395), .QN(n8648) );
  NAND4X0 U9747 ( .IN1(n8398), .IN2(n8397), .IN3(n8396), .IN4(n8648), .QN(
        \a1/N446 ) );
  OA221X1 U9748 ( .IN1(n9149), .IN2(n8960), .IN3(n9149), .IN4(n8400), .IN5(
        n8399), .Q(n8420) );
  NOR2X0 U9749 ( .IN1(n8401), .IN2(n8727), .QN(n8405) );
  NAND2X0 U9750 ( .IN1(n8403), .IN2(n8402), .QN(n8404) );
  NOR2X0 U9751 ( .IN1(n8405), .IN2(n8404), .QN(n8419) );
  INVX0 U9752 ( .INP(n8406), .ZN(n8416) );
  OA21X1 U9753 ( .IN1(n8408), .IN2(n8407), .IN3(n8816), .Q(n8414) );
  NAND4X0 U9754 ( .IN1(n8412), .IN2(n8411), .IN3(n8410), .IN4(n8409), .QN(
        n8413) );
  NOR4X0 U9755 ( .IN1(n8416), .IN2(n8415), .IN3(n8414), .IN4(n8413), .QN(n8418) );
  NAND4X0 U9756 ( .IN1(n8420), .IN2(n8419), .IN3(n8418), .IN4(n8417), .QN(
        \a1/N447 ) );
  NOR2X0 U9757 ( .IN1(n9438), .IN2(n8421), .QN(n8428) );
  OA22X1 U9758 ( .IN1(n8424), .IN2(n8423), .IN3(n9166), .IN4(n8422), .Q(n8425)
         );
  NAND2X0 U9759 ( .IN1(n8426), .IN2(n8425), .QN(n8427) );
  NOR2X0 U9760 ( .IN1(n8428), .IN2(n8427), .QN(n8443) );
  OA21X1 U9761 ( .IN1(n8430), .IN2(n8429), .IN3(n9433), .Q(n8435) );
  NOR2X0 U9762 ( .IN1(n8752), .IN2(n8685), .QN(n8434) );
  NAND2X0 U9763 ( .IN1(n8432), .IN2(n8431), .QN(n8544) );
  NAND4X0 U9764 ( .IN1(n8962), .IN2(n8743), .IN3(n8776), .IN4(n8544), .QN(
        n8433) );
  NOR4X0 U9765 ( .IN1(n8436), .IN2(n8435), .IN3(n8434), .IN4(n8433), .QN(n8442) );
  NAND3X0 U9766 ( .IN1(n8845), .IN2(n8438), .IN3(n8437), .QN(n8439) );
  NAND2X0 U9767 ( .IN1(n8439), .IN2(n8575), .QN(n8440) );
  NAND4X0 U9768 ( .IN1(n8443), .IN2(n8442), .IN3(n8441), .IN4(n8440), .QN(
        \a1/N448 ) );
  OA22X1 U9769 ( .IN1(n8446), .IN2(n8445), .IN3(n9166), .IN4(n8444), .Q(n8466)
         );
  AND3X1 U9770 ( .IN1(n8447), .IN2(n9442), .IN3(n8645), .Q(n8457) );
  NOR2X0 U9771 ( .IN1(n8523), .IN2(n8494), .QN(n8451) );
  NAND2X0 U9772 ( .IN1(n8449), .IN2(n8448), .QN(n8450) );
  NOR2X0 U9773 ( .IN1(n8451), .IN2(n8450), .QN(n8455) );
  NAND4X0 U9774 ( .IN1(n8455), .IN2(n8454), .IN3(n8453), .IN4(n8452), .QN(
        n8456) );
  NOR4X0 U9775 ( .IN1(n8459), .IN2(n8458), .IN3(n8457), .IN4(n8456), .QN(n8465) );
  NAND2X0 U9776 ( .IN1(n8461), .IN2(n8460), .QN(n8464) );
  NAND2X0 U9777 ( .IN1(n8710), .IN2(n8462), .QN(n8463) );
  NAND4X0 U9778 ( .IN1(n8466), .IN2(n8465), .IN3(n8464), .IN4(n8463), .QN(
        \a1/N450 ) );
  NOR2X0 U9779 ( .IN1(n8467), .IN2(n9212), .QN(n8481) );
  NAND3X0 U9780 ( .IN1(n8468), .IN2(n9438), .IN3(n9001), .QN(n8469) );
  OA221X1 U9781 ( .IN1(n8489), .IN2(n8471), .IN3(n8489), .IN4(n8470), .IN5(
        n8469), .Q(n8479) );
  NOR2X0 U9782 ( .IN1(n8473), .IN2(n8472), .QN(n8478) );
  NAND2X0 U9783 ( .IN1(n8475), .IN2(n8474), .QN(n8476) );
  NAND4X0 U9784 ( .IN1(n8479), .IN2(n8478), .IN3(n8477), .IN4(n8476), .QN(
        n8480) );
  NOR4X0 U9785 ( .IN1(n8483), .IN2(n8482), .IN3(n8481), .IN4(n8480), .QN(n8488) );
  NAND2X0 U9786 ( .IN1(n8485), .IN2(n8484), .QN(n8486) );
  NAND4X0 U9787 ( .IN1(n8488), .IN2(n8487), .IN3(n8486), .IN4(n8672), .QN(
        \a1/N451 ) );
  NOR2X0 U9788 ( .IN1(n8489), .IN2(n8527), .QN(n8682) );
  INVX0 U9789 ( .INP(n8682), .ZN(n8490) );
  OA21X1 U9790 ( .IN1(n8491), .IN2(n9122), .IN3(n8490), .Q(n8506) );
  NAND4X0 U9791 ( .IN1(n8493), .IN2(n9067), .IN3(n8834), .IN4(n8492), .QN(
        n8502) );
  OA22X1 U9792 ( .IN1(n9071), .IN2(n8495), .IN3(n8801), .IN4(n8494), .Q(n8500)
         );
  NAND2X0 U9793 ( .IN1(n8496), .IN2(n9001), .QN(n8497) );
  NAND4X0 U9794 ( .IN1(n8500), .IN2(n8499), .IN3(n8498), .IN4(n8497), .QN(
        n8501) );
  NOR4X0 U9795 ( .IN1(n8888), .IN2(n8637), .IN3(n8502), .IN4(n8501), .QN(n8505) );
  NAND4X0 U9796 ( .IN1(n8506), .IN2(n8505), .IN3(n8504), .IN4(n8503), .QN(
        \a1/N452 ) );
  OA22X1 U9797 ( .IN1(n9183), .IN2(n8508), .IN3(n9061), .IN4(n8507), .Q(n8521)
         );
  NOR2X0 U9798 ( .IN1(n8510), .IN2(n8509), .QN(n8517) );
  NAND2X0 U9799 ( .IN1(n8512), .IN2(n8511), .QN(n8513) );
  NAND4X0 U9800 ( .IN1(n8515), .IN2(n8908), .IN3(n8514), .IN4(n8513), .QN(
        n8516) );
  NOR4X0 U9801 ( .IN1(n8519), .IN2(n8518), .IN3(n8517), .IN4(n8516), .QN(n8520) );
  AND4X1 U9802 ( .IN1(n8521), .IN2(n8520), .IN3(n8821), .IN4(n8668), .Q(n8525)
         );
  NAND4X0 U9803 ( .IN1(n8525), .IN2(n8524), .IN3(n8523), .IN4(n8522), .QN(
        \a1/N453 ) );
  OA22X1 U9804 ( .IN1(n8528), .IN2(n8527), .IN3(n9207), .IN4(n8526), .Q(n8543)
         );
  OA21X1 U9805 ( .IN1(n8529), .IN2(n9013), .IN3(n8598), .Q(n8539) );
  NOR2X0 U9806 ( .IN1(n8531), .IN2(n8530), .QN(n8538) );
  NAND4X0 U9807 ( .IN1(n9127), .IN2(n8532), .IN3(n8609), .IN4(n8695), .QN(
        n8537) );
  NAND2X0 U9808 ( .IN1(n8534), .IN2(n8533), .QN(n8957) );
  NAND3X0 U9809 ( .IN1(n8535), .IN2(n8850), .IN3(n8957), .QN(n8536) );
  NOR4X0 U9810 ( .IN1(n8539), .IN2(n8538), .IN3(n8537), .IN4(n8536), .QN(n8542) );
  NAND4X0 U9811 ( .IN1(n8543), .IN2(n8542), .IN3(n8541), .IN4(n8540), .QN(
        \a1/N454 ) );
  NAND2X0 U9812 ( .IN1(n8720), .IN2(n8544), .QN(n8558) );
  NOR2X0 U9813 ( .IN1(n8545), .IN2(n9147), .QN(n8549) );
  NAND2X0 U9814 ( .IN1(n8547), .IN2(n8546), .QN(n8548) );
  NOR2X0 U9815 ( .IN1(n8549), .IN2(n8548), .QN(n8556) );
  NAND3X0 U9816 ( .IN1(n8591), .IN2(n8551), .IN3(n8550), .QN(n8552) );
  NAND2X0 U9817 ( .IN1(n8552), .IN2(n9445), .QN(n8553) );
  NAND4X0 U9818 ( .IN1(n8556), .IN2(n8555), .IN3(n8554), .IN4(n8553), .QN(
        n8557) );
  NOR4X0 U9819 ( .IN1(n8560), .IN2(n8559), .IN3(n8558), .IN4(n8557), .QN(n8565) );
  NAND2X0 U9820 ( .IN1(n8760), .IN2(n8561), .QN(n8562) );
  NAND4X0 U9821 ( .IN1(n8565), .IN2(n8564), .IN3(n8563), .IN4(n8562), .QN(
        \a1/N456 ) );
  NOR2X0 U9822 ( .IN1(n8567), .IN2(n8566), .QN(n8569) );
  OA22X1 U9823 ( .IN1(n8883), .IN2(n8570), .IN3(n8569), .IN4(n8568), .Q(n8586)
         );
  NOR2X0 U9824 ( .IN1(n8572), .IN2(n8571), .QN(n8581) );
  OA22X1 U9825 ( .IN1(n8575), .IN2(n8574), .IN3(n8573), .IN4(n9053), .Q(n8579)
         );
  NAND4X0 U9826 ( .IN1(n8579), .IN2(n8578), .IN3(n8577), .IN4(n8576), .QN(
        n8580) );
  NOR4X0 U9827 ( .IN1(n9171), .IN2(n8682), .IN3(n8581), .IN4(n8580), .QN(n8585) );
  NAND2X0 U9828 ( .IN1(degrees_tmp2[3]), .IN2(n8582), .QN(n8583) );
  NAND4X0 U9829 ( .IN1(n8586), .IN2(n8585), .IN3(n8584), .IN4(n8583), .QN(
        \a1/N457 ) );
  NOR2X0 U9830 ( .IN1(n8754), .IN2(n8587), .QN(n8605) );
  NAND3X0 U9831 ( .IN1(n8898), .IN2(n8588), .IN3(n9099), .QN(n8589) );
  OA21X1 U9832 ( .IN1(degrees_tmp2[3]), .IN2(n8590), .IN3(n8589), .Q(n8603) );
  NAND3X0 U9833 ( .IN1(n8593), .IN2(n8592), .IN3(n8591), .QN(n8594) );
  NAND3X0 U9834 ( .IN1(n8978), .IN2(n8595), .IN3(n8594), .QN(n8601) );
  NAND3X0 U9835 ( .IN1(n8880), .IN2(n8597), .IN3(n8596), .QN(n8599) );
  NAND2X0 U9836 ( .IN1(n8599), .IN2(n8598), .QN(n8600) );
  NAND4X0 U9837 ( .IN1(n8603), .IN2(n8602), .IN3(n8601), .IN4(n8600), .QN(
        n8604) );
  NOR4X0 U9838 ( .IN1(n9066), .IN2(n8606), .IN3(n8605), .IN4(n8604), .QN(n8611) );
  OR2X1 U9839 ( .IN1(n8787), .IN2(n8607), .Q(n8608) );
  NAND4X0 U9840 ( .IN1(n8611), .IN2(n8610), .IN3(n8609), .IN4(n8608), .QN(
        \a1/N458 ) );
  OA22X1 U9841 ( .IN1(n9433), .IN2(n8612), .IN3(n9155), .IN4(n9192), .Q(n8627)
         );
  AO21X1 U9842 ( .IN1(n9072), .IN2(n8613), .IN3(n9031), .Q(n8616) );
  NAND2X0 U9843 ( .IN1(n8932), .IN2(n9436), .QN(n8614) );
  AND3X1 U9844 ( .IN1(n8616), .IN2(n8615), .IN3(n8614), .Q(n8619) );
  NAND4X0 U9845 ( .IN1(n8620), .IN2(n8619), .IN3(n8618), .IN4(n8617), .QN(
        n8621) );
  NOR4X0 U9846 ( .IN1(n8718), .IN2(n8623), .IN3(n8622), .IN4(n8621), .QN(n8626) );
  NAND4X0 U9847 ( .IN1(n8627), .IN2(n8626), .IN3(n8625), .IN4(n8624), .QN(
        \a1/N459 ) );
  NOR2X0 U9848 ( .IN1(n8883), .IN2(n9029), .QN(n8636) );
  INVX0 U9849 ( .INP(n8628), .ZN(n8634) );
  INVX0 U9850 ( .INP(n8629), .ZN(n8632) );
  NAND2X0 U9851 ( .IN1(n8943), .IN2(n8630), .QN(n8631) );
  NAND4X0 U9852 ( .IN1(n8634), .IN2(n8633), .IN3(n8632), .IN4(n8631), .QN(
        n8635) );
  NOR4X0 U9853 ( .IN1(n8638), .IN2(n8637), .IN3(n8636), .IN4(n8635), .QN(n8643) );
  NAND2X0 U9854 ( .IN1(n8640), .IN2(n8639), .QN(n8642) );
  NAND4X0 U9855 ( .IN1(n8644), .IN2(n8643), .IN3(n8642), .IN4(n8641), .QN(
        \a1/N460 ) );
  NAND2X0 U9856 ( .IN1(n8948), .IN2(n8645), .QN(n8652) );
  INVX0 U9857 ( .INP(n8646), .ZN(n8647) );
  OA22X1 U9858 ( .IN1(n8649), .IN2(n8648), .IN3(n9019), .IN4(n8647), .Q(n8650)
         );
  NAND3X0 U9859 ( .IN1(n8652), .IN2(n8651), .IN3(n8650), .QN(n8653) );
  NOR4X0 U9860 ( .IN1(n8656), .IN2(n8655), .IN3(n8654), .IN4(n8653), .QN(n8666) );
  INVX0 U9861 ( .INP(n8657), .ZN(n8661) );
  NOR4X0 U9862 ( .IN1(n8661), .IN2(n8660), .IN3(n8659), .IN4(n8658), .QN(n8665) );
  NAND2X0 U9863 ( .IN1(n8995), .IN2(n8662), .QN(n8663) );
  NAND4X0 U9864 ( .IN1(n8666), .IN2(n8665), .IN3(n8664), .IN4(n8663), .QN(
        \a1/N461 ) );
  NOR2X0 U9865 ( .IN1(n9020), .IN2(n8667), .QN(n8671) );
  NAND2X0 U9866 ( .IN1(n8669), .IN2(n8668), .QN(n8670) );
  NOR2X0 U9867 ( .IN1(n8671), .IN2(n8670), .QN(n8691) );
  NAND2X0 U9868 ( .IN1(n8673), .IN2(n8672), .QN(n8681) );
  AOI22X1 U9869 ( .IN1(n9437), .IN2(n8676), .IN3(n8675), .IN4(n8674), .QN(
        n8679) );
  NAND4X0 U9870 ( .IN1(n8679), .IN2(n8678), .IN3(n8677), .IN4(n9057), .QN(
        n8680) );
  NOR4X0 U9871 ( .IN1(n8683), .IN2(n8682), .IN3(n8681), .IN4(n8680), .QN(n8690) );
  NAND4X0 U9872 ( .IN1(n8686), .IN2(n8685), .IN3(n8684), .IN4(n9100), .QN(
        n8687) );
  NAND2X0 U9873 ( .IN1(n9080), .IN2(n8687), .QN(n8688) );
  NAND4X0 U9874 ( .IN1(n8691), .IN2(n8690), .IN3(n8689), .IN4(n8688), .QN(
        \a1/N462 ) );
  OA22X1 U9875 ( .IN1(n9437), .IN2(n8694), .IN3(n8693), .IN4(n8692), .Q(n8722)
         );
  INVX0 U9876 ( .INP(n8695), .ZN(n8717) );
  AO22X1 U9877 ( .IN1(n8699), .IN2(n8698), .IN3(n8697), .IN4(n8696), .Q(n8716)
         );
  NOR2X0 U9878 ( .IN1(n8700), .IN2(n9205), .QN(n8704) );
  NAND2X0 U9879 ( .IN1(n8702), .IN2(n8701), .QN(n8703) );
  NOR2X0 U9880 ( .IN1(n8704), .IN2(n8703), .QN(n8714) );
  NAND4X0 U9881 ( .IN1(n8708), .IN2(n8707), .IN3(n8706), .IN4(n8705), .QN(
        n8709) );
  NAND2X0 U9882 ( .IN1(n8710), .IN2(n8709), .QN(n8711) );
  NAND4X0 U9883 ( .IN1(n8714), .IN2(n8713), .IN3(n8712), .IN4(n8711), .QN(
        n8715) );
  NOR4X0 U9884 ( .IN1(n8718), .IN2(n8717), .IN3(n8716), .IN4(n8715), .QN(n8721) );
  NAND4X0 U9885 ( .IN1(n8722), .IN2(n8721), .IN3(n8720), .IN4(n8719), .QN(
        \a1/N463 ) );
  NOR2X0 U9886 ( .IN1(n8723), .IN2(n9010), .QN(n8725) );
  OA22X1 U9887 ( .IN1(n8727), .IN2(n8726), .IN3(n8725), .IN4(n8724), .Q(n8750)
         );
  NOR2X0 U9888 ( .IN1(n8968), .IN2(n8728), .QN(n8746) );
  INVX0 U9889 ( .INP(n8729), .ZN(n9148) );
  OA21X1 U9890 ( .IN1(n8731), .IN2(n9148), .IN3(n8730), .Q(n8741) );
  NAND2X0 U9891 ( .IN1(n8733), .IN2(n8732), .QN(n8740) );
  NAND2X0 U9892 ( .IN1(n9037), .IN2(n8734), .QN(n8735) );
  NAND4X0 U9893 ( .IN1(n8738), .IN2(n8737), .IN3(n8736), .IN4(n8735), .QN(
        n8739) );
  NOR4X0 U9894 ( .IN1(n8742), .IN2(n8741), .IN3(n8740), .IN4(n8739), .QN(n8744) );
  NAND2X0 U9895 ( .IN1(n8744), .IN2(n8743), .QN(n8745) );
  NOR2X0 U9896 ( .IN1(n8746), .IN2(n8745), .QN(n8749) );
  NAND4X0 U9897 ( .IN1(n8750), .IN2(n8749), .IN3(n8748), .IN4(n8747), .QN(
        \a1/N464 ) );
  NOR2X0 U9898 ( .IN1(n8752), .IN2(n8751), .QN(n8771) );
  NAND2X0 U9899 ( .IN1(n8754), .IN2(n8753), .QN(n8758) );
  INVX0 U9900 ( .INP(n8755), .ZN(n8757) );
  NAND4X0 U9901 ( .IN1(n8758), .IN2(n9103), .IN3(n8757), .IN4(n8756), .QN(
        n8769) );
  OA22X1 U9902 ( .IN1(n9183), .IN2(n8761), .IN3(n8760), .IN4(n8759), .Q(n8767)
         );
  OA22X1 U9903 ( .IN1(n8764), .IN2(n8763), .IN3(degrees_tmp2[3]), .IN4(n8762), 
        .Q(n8766) );
  NAND4X0 U9904 ( .IN1(n8767), .IN2(n8766), .IN3(n8868), .IN4(n8765), .QN(
        n8768) );
  OR4X1 U9905 ( .IN1(n8771), .IN2(n8770), .IN3(n8769), .IN4(n8768), .Q(
        \a1/N465 ) );
  NOR2X0 U9906 ( .IN1(degrees_tmp2[0]), .IN2(n8772), .QN(n8794) );
  OA21X1 U9907 ( .IN1(n8774), .IN2(n8773), .IN3(n9445), .Q(n8785) );
  NAND4X0 U9908 ( .IN1(n8778), .IN2(n8777), .IN3(n8776), .IN4(n8775), .QN(
        n8784) );
  OAI22X1 U9909 ( .IN1(n8782), .IN2(n8781), .IN3(n8780), .IN4(n8779), .QN(
        n8783) );
  NOR4X0 U9910 ( .IN1(n8786), .IN2(n8785), .IN3(n8784), .IN4(n8783), .QN(n8791) );
  NAND2X0 U9911 ( .IN1(n8788), .IN2(n8787), .QN(n8789) );
  NAND4X0 U9912 ( .IN1(n8792), .IN2(n8791), .IN3(n8790), .IN4(n8789), .QN(
        n8793) );
  AO221X1 U9913 ( .IN1(n8796), .IN2(n8795), .IN3(n8796), .IN4(n8794), .IN5(
        n8793), .Q(\a1/N466 ) );
  NOR2X0 U9914 ( .IN1(degrees_tmp2[3]), .IN2(n8797), .QN(n8813) );
  NAND4X0 U9915 ( .IN1(n8801), .IN2(n8800), .IN3(n8799), .IN4(n8798), .QN(
        n8812) );
  NAND4X0 U9916 ( .IN1(n8804), .IN2(n8892), .IN3(n8803), .IN4(n8802), .QN(
        n8811) );
  NAND2X0 U9917 ( .IN1(n8805), .IN2(n8822), .QN(n8806) );
  NAND4X0 U9918 ( .IN1(n8809), .IN2(n8808), .IN3(n8807), .IN4(n8806), .QN(
        n8810) );
  OR4X1 U9919 ( .IN1(n8813), .IN2(n8812), .IN3(n8811), .IN4(n8810), .Q(
        \a1/N467 ) );
  OA21X1 U9920 ( .IN1(n8816), .IN2(n8815), .IN3(n8814), .Q(n8837) );
  INVX0 U9921 ( .INP(n8817), .ZN(n8833) );
  NAND4X0 U9922 ( .IN1(n8821), .IN2(n8820), .IN3(n8819), .IN4(n8818), .QN(
        n8831) );
  NAND2X0 U9923 ( .IN1(n8823), .IN2(n8822), .QN(n8828) );
  NAND3X0 U9924 ( .IN1(n8826), .IN2(n8825), .IN3(n8824), .QN(n8827) );
  NAND4X0 U9925 ( .IN1(n8829), .IN2(n9110), .IN3(n8828), .IN4(n8827), .QN(
        n8830) );
  NOR4X0 U9926 ( .IN1(n8833), .IN2(n8832), .IN3(n8831), .IN4(n8830), .QN(n8836) );
  NAND4X0 U9927 ( .IN1(n8837), .IN2(n8836), .IN3(n8835), .IN4(n8834), .QN(
        \a1/N468 ) );
  NAND4X0 U9928 ( .IN1(n8840), .IN2(n8839), .IN3(n8838), .IN4(n8925), .QN(
        n8854) );
  AO21X1 U9929 ( .IN1(n8842), .IN2(n8841), .IN3(n9048), .Q(n8843) );
  NAND4X0 U9930 ( .IN1(n8846), .IN2(n8845), .IN3(n8844), .IN4(n8843), .QN(
        n8853) );
  NAND2X0 U9931 ( .IN1(n8848), .IN2(n8847), .QN(n8849) );
  NAND4X0 U9932 ( .IN1(n8851), .IN2(n8868), .IN3(n8850), .IN4(n8849), .QN(
        n8852) );
  NOR4X0 U9933 ( .IN1(n8855), .IN2(n8854), .IN3(n8853), .IN4(n8852), .QN(n8858) );
  NAND4X0 U9934 ( .IN1(n8858), .IN2(n9118), .IN3(n8857), .IN4(n8856), .QN(
        \a1/N469 ) );
  NOR2X0 U9935 ( .IN1(n8728), .IN2(n8859), .QN(n8874) );
  NAND2X0 U9936 ( .IN1(n8962), .IN2(n8860), .QN(n8873) );
  NAND2X0 U9937 ( .IN1(n8862), .IN2(n8861), .QN(n8863) );
  NAND4X0 U9938 ( .IN1(n8866), .IN2(n8865), .IN3(n8864), .IN4(n8863), .QN(
        n8872) );
  NAND4X0 U9939 ( .IN1(n8870), .IN2(n8869), .IN3(n8868), .IN4(n8867), .QN(
        n8871) );
  NOR4X0 U9940 ( .IN1(n8874), .IN2(n8873), .IN3(n8872), .IN4(n8871), .QN(n8879) );
  NAND2X0 U9941 ( .IN1(n8876), .IN2(n8875), .QN(n8877) );
  NAND4X0 U9942 ( .IN1(n8879), .IN2(n8878), .IN3(n9101), .IN4(n8877), .QN(
        \a1/N470 ) );
  OA22X1 U9943 ( .IN1(n9125), .IN2(n8882), .IN3(n8881), .IN4(n8880), .Q(n8902)
         );
  OA221X1 U9944 ( .IN1(n8884), .IN2(n9131), .IN3(n8884), .IN4(n9190), .IN5(
        n8883), .Q(n8897) );
  INVX0 U9945 ( .INP(n8885), .ZN(n8887) );
  OA21X1 U9946 ( .IN1(n8888), .IN2(n8887), .IN3(n8886), .Q(n8896) );
  OA22X1 U9947 ( .IN1(n8890), .IN2(n9192), .IN3(n9031), .IN4(n8889), .Q(n8894)
         );
  NAND4X0 U9948 ( .IN1(n8894), .IN2(n8893), .IN3(n8892), .IN4(n8891), .QN(
        n8895) );
  NOR3X0 U9949 ( .IN1(n8897), .IN2(n8896), .IN3(n8895), .QN(n8901) );
  NAND2X0 U9950 ( .IN1(n8898), .IN2(n9131), .QN(n8899) );
  NAND4X0 U9951 ( .IN1(n8902), .IN2(n8901), .IN3(n8900), .IN4(n8899), .QN(
        \a1/N471 ) );
  OA22X1 U9952 ( .IN1(n9071), .IN2(n8905), .IN3(n8904), .IN4(n8903), .Q(n8907)
         );
  NAND2X0 U9953 ( .IN1(n8907), .IN2(n8906), .QN(n8919) );
  OA221X1 U9954 ( .IN1(n8909), .IN2(n9119), .IN3(n8909), .IN4(n9085), .IN5(
        n8908), .Q(n8912) );
  NAND4X0 U9955 ( .IN1(n8912), .IN2(n8911), .IN3(n8910), .IN4(n9146), .QN(
        n8918) );
  NAND4X0 U9956 ( .IN1(n8916), .IN2(n8915), .IN3(n8914), .IN4(n8913), .QN(
        n8917) );
  OR4X1 U9957 ( .IN1(n8920), .IN2(n8919), .IN3(n8918), .IN4(n8917), .Q(
        \a1/N472 ) );
  OA22X1 U9958 ( .IN1(n8728), .IN2(n8922), .IN3(n9125), .IN4(n8921), .Q(n8936)
         );
  NOR2X0 U9959 ( .IN1(n8924), .IN2(n8923), .QN(n8935) );
  NAND4X0 U9960 ( .IN1(n8928), .IN2(n8927), .IN3(n8926), .IN4(n8925), .QN(
        n8929) );
  NOR4X0 U9961 ( .IN1(n8932), .IN2(n8931), .IN3(n8930), .IN4(n8929), .QN(n8934) );
  NAND4X0 U9962 ( .IN1(n8936), .IN2(n8935), .IN3(n8934), .IN4(n8933), .QN(
        \a1/N473 ) );
  OA22X1 U9963 ( .IN1(n8940), .IN2(n8939), .IN3(n8938), .IN4(n8937), .Q(n8959)
         );
  NOR2X0 U9964 ( .IN1(n9001), .IN2(n8941), .QN(n8952) );
  NOR2X0 U9965 ( .IN1(n8943), .IN2(n8942), .QN(n8946) );
  NAND2X0 U9966 ( .IN1(n8944), .IN2(n9445), .QN(n8945) );
  NAND2X0 U9967 ( .IN1(n8946), .IN2(n8945), .QN(n8951) );
  AO22X1 U9968 ( .IN1(degrees_tmp2[3]), .IN2(n8949), .IN3(n8948), .IN4(n8947), 
        .Q(n8950) );
  NOR4X0 U9969 ( .IN1(n8953), .IN2(n8952), .IN3(n8951), .IN4(n8950), .QN(n8958) );
  NAND2X0 U9970 ( .IN1(n8955), .IN2(n8954), .QN(n8956) );
  NAND4X0 U9971 ( .IN1(n8959), .IN2(n8958), .IN3(n8957), .IN4(n8956), .QN(
        \a1/N474 ) );
  OA22X1 U9972 ( .IN1(n8995), .IN2(n8996), .IN3(n8960), .IN4(n9166), .Q(n8976)
         );
  NOR2X0 U9973 ( .IN1(n8978), .IN2(n8961), .QN(n8971) );
  INVX0 U9974 ( .INP(n9171), .ZN(n8963) );
  NAND3X0 U9975 ( .IN1(n8964), .IN2(n8963), .IN3(n8962), .QN(n8970) );
  NAND4X0 U9976 ( .IN1(n8968), .IN2(n8967), .IN3(n8966), .IN4(n8965), .QN(
        n8969) );
  NOR4X0 U9977 ( .IN1(n8972), .IN2(n8971), .IN3(n8970), .IN4(n8969), .QN(n8975) );
  NAND4X0 U9978 ( .IN1(n8976), .IN2(n8975), .IN3(n8974), .IN4(n8973), .QN(
        \a1/N475 ) );
  NOR2X0 U9979 ( .IN1(n8978), .IN2(n8977), .QN(n8981) );
  NOR2X0 U9980 ( .IN1(n9433), .IN2(n8979), .QN(n8980) );
  NOR4X0 U9981 ( .IN1(n8983), .IN2(n8982), .IN3(n8981), .IN4(n8980), .QN(n9000) );
  NOR2X0 U9982 ( .IN1(n8984), .IN2(n9083), .QN(n8992) );
  NOR2X0 U9983 ( .IN1(n8986), .IN2(n8985), .QN(n8990) );
  NAND2X0 U9984 ( .IN1(n8988), .IN2(n8987), .QN(n8989) );
  NAND2X0 U9985 ( .IN1(n8990), .IN2(n8989), .QN(n8991) );
  NOR4X0 U9986 ( .IN1(n8994), .IN2(n8993), .IN3(n8992), .IN4(n8991), .QN(n8999) );
  OR2X1 U9987 ( .IN1(n8996), .IN2(n8995), .Q(n8997) );
  NAND4X0 U9988 ( .IN1(n9000), .IN2(n8999), .IN3(n8998), .IN4(n8997), .QN(
        \a1/N476 ) );
  OA22X1 U9989 ( .IN1(n9004), .IN2(n9003), .IN3(n9002), .IN4(n9001), .Q(n9018)
         );
  OA21X1 U9990 ( .IN1(n9435), .IN2(n9183), .IN3(n9005), .Q(n9012) );
  NOR2X0 U9991 ( .IN1(n9436), .IN2(n9006), .QN(n9007) );
  OR4X1 U9992 ( .IN1(n9010), .IN2(n9009), .IN3(n9008), .IN4(n9007), .Q(n9011)
         );
  NOR4X0 U9993 ( .IN1(n9014), .IN2(n9013), .IN3(n9012), .IN4(n9011), .QN(n9017) );
  NAND4X0 U9994 ( .IN1(n9018), .IN2(n9017), .IN3(n9016), .IN4(n9015), .QN(
        \a1/N478 ) );
  OA22X1 U9995 ( .IN1(n9054), .IN2(n9020), .IN3(n9019), .IN4(n9079), .Q(n9021)
         );
  OA221X1 U9996 ( .IN1(n9023), .IN2(n9102), .IN3(n9023), .IN4(n9022), .IN5(
        n9021), .Q(n9044) );
  AOI21X1 U9997 ( .IN1(n9026), .IN2(n9025), .IN3(n9024), .QN(n9043) );
  NAND4X0 U9998 ( .IN1(n9030), .IN2(n9029), .IN3(n9028), .IN4(n9027), .QN(
        n9034) );
  OA221X1 U9999 ( .IN1(n9034), .IN2(n9033), .IN3(n9034), .IN4(n9032), .IN5(
        n9031), .Q(n9040) );
  AO22X1 U10000 ( .IN1(n9037), .IN2(n9036), .IN3(n9035), .IN4(n9155), .Q(n9038) );
  NOR4X0 U10001 ( .IN1(n9040), .IN2(n9062), .IN3(n9039), .IN4(n9038), .QN(
        n9042) );
  NAND4X0 U10002 ( .IN1(n9044), .IN2(n9043), .IN3(n9042), .IN4(n9041), .QN(
        \a1/N479 ) );
  NAND3X0 U10003 ( .IN1(n9047), .IN2(n9046), .IN3(n9045), .QN(n9049) );
  AO21X1 U10004 ( .IN1(n9050), .IN2(n9049), .IN3(n9048), .Q(n9051) );
  OA221X1 U10005 ( .IN1(n9054), .IN2(n9053), .IN3(n9054), .IN4(n9052), .IN5(
        n9051), .Q(n9070) );
  OA21X1 U10006 ( .IN1(n9442), .IN2(n9056), .IN3(n9055), .Q(n9069) );
  NAND2X0 U10007 ( .IN1(n9058), .IN2(n9057), .QN(n9059) );
  AO22X1 U10008 ( .IN1(n9062), .IN2(n9061), .IN3(n9060), .IN4(n9059), .Q(n9063) );
  NOR4X0 U10009 ( .IN1(n9066), .IN2(n9065), .IN3(n9064), .IN4(n9063), .QN(
        n9068) );
  NAND4X0 U10010 ( .IN1(n9070), .IN2(n9069), .IN3(n9068), .IN4(n9067), .QN(
        \a1/N480 ) );
  OA22X1 U10011 ( .IN1(n9073), .IN2(n9072), .IN3(n9071), .IN4(n9098), .Q(n9097) );
  NOR3X0 U10012 ( .IN1(n9076), .IN2(n9075), .IN3(n9074), .QN(n9078) );
  OA221X1 U10013 ( .IN1(n9080), .IN2(n9079), .IN3(n9181), .IN4(n9078), .IN5(
        n9077), .Q(n9096) );
  NOR2X0 U10014 ( .IN1(n9081), .IN2(n9433), .QN(n9090) );
  AO221X1 U10015 ( .IN1(n9085), .IN2(n9084), .IN3(n9085), .IN4(n9083), .IN5(
        n9082), .Q(n9086) );
  NAND3X0 U10016 ( .IN1(n9088), .IN2(n9087), .IN3(n9086), .QN(n9089) );
  NOR4X0 U10017 ( .IN1(n9092), .IN2(n9091), .IN3(n9090), .IN4(n9089), .QN(
        n9095) );
  NAND2X0 U10018 ( .IN1(n9435), .IN2(n9093), .QN(n9094) );
  NAND4X0 U10019 ( .IN1(n9097), .IN2(n9096), .IN3(n9095), .IN4(n9094), .QN(
        \a1/N481 ) );
  OA22X1 U10020 ( .IN1(n8728), .IN2(n9100), .IN3(n9099), .IN4(n9098), .Q(n9121) );
  NAND2X0 U10021 ( .IN1(n9102), .IN2(n9101), .QN(n9116) );
  INVX0 U10022 ( .INP(n9103), .ZN(n9106) );
  AO22X1 U10023 ( .IN1(n9437), .IN2(n9106), .IN3(n9105), .IN4(n9104), .Q(n9115) );
  OA22X1 U10024 ( .IN1(n9440), .IN2(n9109), .IN3(n9108), .IN4(n9107), .Q(n9113) );
  NAND4X0 U10025 ( .IN1(n9113), .IN2(n9112), .IN3(n9111), .IN4(n9110), .QN(
        n9114) );
  NOR4X0 U10026 ( .IN1(n9117), .IN2(n9116), .IN3(n9115), .IN4(n9114), .QN(
        n9120) );
  NAND4X0 U10027 ( .IN1(n9121), .IN2(n9120), .IN3(n9119), .IN4(n9118), .QN(
        \a1/N482 ) );
  AOI22X1 U10028 ( .IN1(n9125), .IN2(n9124), .IN3(n9123), .IN4(n9122), .QN(
        n9142) );
  NAND2X0 U10029 ( .IN1(n9127), .IN2(n9126), .QN(n9137) );
  OAI22X1 U10030 ( .IN1(n9131), .IN2(n9130), .IN3(n9129), .IN4(n9128), .QN(
        n9136) );
  AO22X1 U10031 ( .IN1(degrees_tmp2[0]), .IN2(n9134), .IN3(n9133), .IN4(n9132), 
        .Q(n9135) );
  NOR4X0 U10032 ( .IN1(n9138), .IN2(n9137), .IN3(n9136), .IN4(n9135), .QN(
        n9141) );
  NAND4X0 U10033 ( .IN1(n9142), .IN2(n9141), .IN3(n9140), .IN4(n9139), .QN(
        n9143) );
  AO221X1 U10034 ( .IN1(n9435), .IN2(n9145), .IN3(n9435), .IN4(n9144), .IN5(
        n9143), .Q(\a1/N483 ) );
  INVX0 U10035 ( .INP(n9146), .ZN(n9163) );
  NAND2X0 U10036 ( .IN1(n9148), .IN2(n9147), .QN(n9153) );
  NAND2X0 U10037 ( .IN1(n9150), .IN2(n9149), .QN(n9152) );
  NAND3X0 U10038 ( .IN1(n9153), .IN2(n9152), .IN3(n9151), .QN(n9162) );
  INVX0 U10039 ( .INP(n9154), .ZN(n9158) );
  NAND2X0 U10040 ( .IN1(n9156), .IN2(n9155), .QN(n9157) );
  NAND4X0 U10041 ( .IN1(n9160), .IN2(n9159), .IN3(n9158), .IN4(n9157), .QN(
        n9161) );
  NOR4X0 U10042 ( .IN1(n9164), .IN2(n9163), .IN3(n9162), .IN4(n9161), .QN(
        n9170) );
  OR2X1 U10043 ( .IN1(n9166), .IN2(n9165), .Q(n9167) );
  NAND4X0 U10044 ( .IN1(n9170), .IN2(n9169), .IN3(n9168), .IN4(n9167), .QN(
        \a1/N484 ) );
  AOI21X1 U10045 ( .IN1(n9173), .IN2(n9172), .IN3(n9171), .QN(n9180) );
  NOR4X0 U10046 ( .IN1(n9176), .IN2(n9175), .IN3(n9174), .IN4(n9186), .QN(
        n9179) );
  NAND4X0 U10047 ( .IN1(n9180), .IN2(n9179), .IN3(n9178), .IN4(n9177), .QN(
        \a1/N485 ) );
  AO22X1 U10048 ( .IN1(n9184), .IN2(n9183), .IN3(n9182), .IN4(n9181), .Q(n9185) );
  NOR4X0 U10049 ( .IN1(n9188), .IN2(n9187), .IN3(n9186), .IN4(n9185), .QN(
        n9194) );
  NAND2X0 U10050 ( .IN1(n9190), .IN2(n9189), .QN(n9191) );
  NAND4X0 U10051 ( .IN1(n9194), .IN2(n9193), .IN3(n9192), .IN4(n9191), .QN(
        \a1/N486 ) );
  NAND2X0 U10052 ( .IN1(n9195), .IN2(n9166), .QN(n9199) );
  AO21X1 U10053 ( .IN1(n9437), .IN2(n9197), .IN3(n9196), .Q(n9198) );
  NAND4X0 U10054 ( .IN1(n9201), .IN2(n9200), .IN3(n9199), .IN4(n9198), .QN(
        \a1/N487 ) );
  NOR2X0 U10055 ( .IN1(n9203), .IN2(n9202), .QN(n9206) );
  NAND3X0 U10056 ( .IN1(n9205), .IN2(n9206), .IN3(n9204), .QN(\a1/N489 ) );
  OA21X1 U10057 ( .IN1(n9208), .IN2(n9207), .IN3(n9206), .Q(n9214) );
  NAND2X0 U10058 ( .IN1(n9210), .IN2(n9209), .QN(n9211) );
  NAND4X0 U10059 ( .IN1(n9214), .IN2(n9213), .IN3(n9212), .IN4(n9211), .QN(
        \a1/N490 ) );
  NOR2X0 U10060 ( .IN1(n9216), .IN2(n9215), .QN(n9222) );
  NOR2X0 U10061 ( .IN1(n9218), .IN2(n9217), .QN(n9221) );
  NAND2X0 U10062 ( .IN1(degrees[7]), .IN2(n9219), .QN(n9220) );
  NAND3X0 U10063 ( .IN1(n9222), .IN2(n9221), .IN3(n9220), .QN(N356) );
  INVX0 U10064 ( .INP(actv[2]), .ZN(n9224) );
  NAND2X0 U10065 ( .IN1(actv[0]), .IN2(n9224), .QN(n9223) );
  OR2X1 U10066 ( .IN1(actv[1]), .IN2(n9223), .Q(n9239) );
  INVX0 U10067 ( .INP(n9239), .ZN(n9426) );
  INVX0 U10068 ( .INP(actv[1]), .ZN(n9225) );
  NAND3X0 U10069 ( .IN1(actv[2]), .IN2(actv[0]), .IN3(n9225), .QN(n9235) );
  INVX0 U10070 ( .INP(n9235), .ZN(n9419) );
  AO22X1 U10071 ( .IN1(n9426), .IN2(data_cos[63]), .IN3(n9419), .IN4(
        data_cot[63]), .Q(n9229) );
  NOR3X0 U10072 ( .IN1(actv[1]), .IN2(actv[2]), .IN3(actv[0]), .QN(n9428) );
  NAND3X0 U10073 ( .IN1(actv[1]), .IN2(actv[0]), .IN3(n9224), .QN(n9230) );
  INVX0 U10074 ( .INP(n9230), .ZN(n9427) );
  AO22X1 U10075 ( .IN1(n9428), .IN2(data_sin[63]), .IN3(n9427), .IN4(
        data_csc[63]), .Q(n9228) );
  NAND2X0 U10076 ( .IN1(actv[2]), .IN2(n9225), .QN(n9226) );
  NOR2X0 U10077 ( .IN1(actv[0]), .IN2(n9226), .QN(n9429) );
  AO22X1 U10078 ( .IN1(n4561), .IN2(data_tan[63]), .IN3(n9429), .IN4(
        data_sec[63]), .Q(n9227) );
  OR3X1 U10079 ( .IN1(n9229), .IN2(n9228), .IN3(n9227), .Q(N449) );
  NAND2X0 U10080 ( .IN1(n4559), .IN2(data_tan[62]), .QN(n9234) );
  NAND2X0 U10081 ( .IN1(n9429), .IN2(data_sec[62]), .QN(n9233) );
  NAND2X0 U10082 ( .IN1(n9419), .IN2(data_cot[62]), .QN(n9232) );
  INVX0 U10083 ( .INP(n9230), .ZN(n9420) );
  NAND2X0 U10084 ( .IN1(n9420), .IN2(data_csc[62]), .QN(n9231) );
  NAND4X0 U10085 ( .IN1(n9234), .IN2(n9233), .IN3(n9232), .IN4(n9231), .QN(
        N448) );
  AO22X1 U10086 ( .IN1(n9426), .IN2(data_cos[61]), .IN3(n9420), .IN4(
        data_csc[61]), .Q(n9238) );
  AO22X1 U10087 ( .IN1(n9429), .IN2(data_sec[61]), .IN3(n9428), .IN4(
        data_sin[61]), .Q(n9237) );
  INVX0 U10088 ( .INP(n9235), .ZN(n9425) );
  AO22X1 U10089 ( .IN1(n4558), .IN2(data_tan[61]), .IN3(n9425), .IN4(
        data_cot[61]), .Q(n9236) );
  OR3X1 U10090 ( .IN1(n9238), .IN2(n9237), .IN3(n9236), .Q(N447) );
  AO22X1 U10091 ( .IN1(n9419), .IN2(data_cot[60]), .IN3(n9427), .IN4(
        data_csc[60]), .Q(n9242) );
  INVX0 U10092 ( .INP(n9239), .ZN(n9421) );
  AO22X1 U10093 ( .IN1(n4558), .IN2(data_tan[60]), .IN3(n9421), .IN4(
        data_cos[60]), .Q(n9241) );
  AO22X1 U10094 ( .IN1(n9429), .IN2(data_sec[60]), .IN3(n9428), .IN4(
        data_sin[60]), .Q(n9240) );
  OR3X1 U10095 ( .IN1(n9242), .IN2(n9241), .IN3(n9240), .Q(N446) );
  AO22X1 U10096 ( .IN1(n9429), .IN2(data_sec[59]), .IN3(n9426), .IN4(
        data_cos[59]), .Q(n9245) );
  AO22X1 U10097 ( .IN1(n9428), .IN2(data_sin[59]), .IN3(n9420), .IN4(
        data_csc[59]), .Q(n9244) );
  AO22X1 U10098 ( .IN1(n4558), .IN2(data_tan[59]), .IN3(n9425), .IN4(
        data_cot[59]), .Q(n9243) );
  OR3X1 U10099 ( .IN1(n9245), .IN2(n9244), .IN3(n9243), .Q(N445) );
  AO22X1 U10100 ( .IN1(n4560), .IN2(data_tan[58]), .IN3(n9427), .IN4(
        data_csc[58]), .Q(n9248) );
  AO22X1 U10101 ( .IN1(n9429), .IN2(data_sec[58]), .IN3(n9426), .IN4(
        data_cos[58]), .Q(n9247) );
  AO22X1 U10102 ( .IN1(n9425), .IN2(data_cot[58]), .IN3(n9428), .IN4(
        data_sin[58]), .Q(n9246) );
  OR3X1 U10103 ( .IN1(n9248), .IN2(n9247), .IN3(n9246), .Q(N444) );
  AO22X1 U10104 ( .IN1(n9429), .IN2(data_sec[57]), .IN3(n9425), .IN4(
        data_cot[57]), .Q(n9251) );
  AO22X1 U10105 ( .IN1(n4561), .IN2(data_tan[57]), .IN3(n9420), .IN4(
        data_csc[57]), .Q(n9250) );
  AO22X1 U10106 ( .IN1(n9426), .IN2(data_cos[57]), .IN3(n9428), .IN4(
        data_sin[57]), .Q(n9249) );
  OR3X1 U10107 ( .IN1(n9251), .IN2(n9250), .IN3(n9249), .Q(N443) );
  AO22X1 U10108 ( .IN1(n9419), .IN2(data_cot[56]), .IN3(n9428), .IN4(
        data_sin[56]), .Q(n9254) );
  AO22X1 U10109 ( .IN1(n9429), .IN2(data_sec[56]), .IN3(n9427), .IN4(
        data_csc[56]), .Q(n9253) );
  AO22X1 U10110 ( .IN1(n4560), .IN2(data_tan[56]), .IN3(n9421), .IN4(
        data_cos[56]), .Q(n9252) );
  OR3X1 U10111 ( .IN1(n9254), .IN2(n9253), .IN3(n9252), .Q(N442) );
  AO22X1 U10112 ( .IN1(n4559), .IN2(data_tan[55]), .IN3(n9421), .IN4(
        data_cos[55]), .Q(n9257) );
  AO22X1 U10113 ( .IN1(n9428), .IN2(data_sin[55]), .IN3(n9420), .IN4(
        data_csc[55]), .Q(n9256) );
  AO22X1 U10114 ( .IN1(n9429), .IN2(data_sec[55]), .IN3(n9425), .IN4(
        data_cot[55]), .Q(n9255) );
  OR3X1 U10115 ( .IN1(n9257), .IN2(n9256), .IN3(n9255), .Q(N441) );
  AO22X1 U10116 ( .IN1(n4559), .IN2(data_tan[54]), .IN3(n9426), .IN4(
        data_cos[54]), .Q(n9260) );
  AO22X1 U10117 ( .IN1(n9428), .IN2(data_sin[54]), .IN3(n9427), .IN4(
        data_csc[54]), .Q(n9259) );
  AO22X1 U10118 ( .IN1(n9429), .IN2(data_sec[54]), .IN3(n9425), .IN4(
        data_cot[54]), .Q(n9258) );
  OR3X1 U10119 ( .IN1(n9260), .IN2(n9259), .IN3(n9258), .Q(N440) );
  AO22X1 U10120 ( .IN1(n9429), .IN2(data_sec[53]), .IN3(n9420), .IN4(
        data_csc[53]), .Q(n9263) );
  AO22X1 U10121 ( .IN1(n4559), .IN2(data_tan[53]), .IN3(n9421), .IN4(
        data_cos[53]), .Q(n9262) );
  AO22X1 U10122 ( .IN1(n9425), .IN2(data_cot[53]), .IN3(n9428), .IN4(
        data_sin[53]), .Q(n9261) );
  OR3X1 U10123 ( .IN1(n9263), .IN2(n9262), .IN3(n9261), .Q(N439) );
  AO22X1 U10124 ( .IN1(n9426), .IN2(data_cos[52]), .IN3(n9427), .IN4(
        data_csc[52]), .Q(n9266) );
  AO22X1 U10125 ( .IN1(n9429), .IN2(data_sec[52]), .IN3(n9419), .IN4(
        data_cot[52]), .Q(n9265) );
  AO22X1 U10126 ( .IN1(n4561), .IN2(data_tan[52]), .IN3(n9428), .IN4(
        data_sin[52]), .Q(n9264) );
  OR3X1 U10127 ( .IN1(n9266), .IN2(n9265), .IN3(n9264), .Q(N438) );
  AO22X1 U10128 ( .IN1(n9426), .IN2(data_cos[51]), .IN3(n9420), .IN4(
        data_csc[51]), .Q(n9269) );
  AO22X1 U10129 ( .IN1(n9429), .IN2(data_sec[51]), .IN3(n9419), .IN4(
        data_cot[51]), .Q(n9268) );
  AO22X1 U10130 ( .IN1(n4560), .IN2(data_tan[51]), .IN3(n9428), .IN4(
        data_sin[51]), .Q(n9267) );
  OR3X1 U10131 ( .IN1(n9269), .IN2(n9268), .IN3(n9267), .Q(N437) );
  AO22X1 U10132 ( .IN1(n4561), .IN2(data_tan[50]), .IN3(n9421), .IN4(
        data_cos[50]), .Q(n9272) );
  AO22X1 U10133 ( .IN1(n9429), .IN2(data_sec[50]), .IN3(n9427), .IN4(
        data_csc[50]), .Q(n9271) );
  AO22X1 U10134 ( .IN1(n9419), .IN2(data_cot[50]), .IN3(n9428), .IN4(
        data_sin[50]), .Q(n9270) );
  OR3X1 U10135 ( .IN1(n9272), .IN2(n9271), .IN3(n9270), .Q(N436) );
  AO22X1 U10136 ( .IN1(n4560), .IN2(data_tan[49]), .IN3(n9429), .IN4(
        data_sec[49]), .Q(n9275) );
  AO22X1 U10137 ( .IN1(n9428), .IN2(data_sin[49]), .IN3(n9427), .IN4(
        data_csc[49]), .Q(n9274) );
  AO22X1 U10138 ( .IN1(n9426), .IN2(data_cos[49]), .IN3(n9419), .IN4(
        data_cot[49]), .Q(n9273) );
  OR3X1 U10139 ( .IN1(n9275), .IN2(n9274), .IN3(n9273), .Q(N435) );
  AO22X1 U10140 ( .IN1(n9428), .IN2(data_sin[48]), .IN3(n9427), .IN4(
        data_csc[48]), .Q(n9278) );
  AO22X1 U10141 ( .IN1(n9429), .IN2(data_sec[48]), .IN3(n9426), .IN4(
        data_cos[48]), .Q(n9277) );
  AO22X1 U10142 ( .IN1(n4561), .IN2(data_tan[48]), .IN3(n9425), .IN4(
        data_cot[48]), .Q(n9276) );
  OR3X1 U10143 ( .IN1(n9278), .IN2(n9277), .IN3(n9276), .Q(N434) );
  AO22X1 U10144 ( .IN1(n9421), .IN2(data_cos[47]), .IN3(n9427), .IN4(
        data_csc[47]), .Q(n9281) );
  AO22X1 U10145 ( .IN1(n9429), .IN2(data_sec[47]), .IN3(n9419), .IN4(
        data_cot[47]), .Q(n9280) );
  AO22X1 U10146 ( .IN1(n4560), .IN2(data_tan[47]), .IN3(n9428), .IN4(
        data_sin[47]), .Q(n9279) );
  OR3X1 U10147 ( .IN1(n9281), .IN2(n9280), .IN3(n9279), .Q(N433) );
  AO22X1 U10148 ( .IN1(n9421), .IN2(data_cos[46]), .IN3(n9419), .IN4(
        data_cot[46]), .Q(n9284) );
  AO22X1 U10149 ( .IN1(n9429), .IN2(data_sec[46]), .IN3(n9427), .IN4(
        data_csc[46]), .Q(n9283) );
  AO22X1 U10150 ( .IN1(n4559), .IN2(data_tan[46]), .IN3(n9428), .IN4(
        data_sin[46]), .Q(n9282) );
  OR3X1 U10151 ( .IN1(n9284), .IN2(n9283), .IN3(n9282), .Q(N432) );
  AO22X1 U10152 ( .IN1(n9425), .IN2(data_cot[45]), .IN3(n9428), .IN4(
        data_sin[45]), .Q(n9287) );
  AO22X1 U10153 ( .IN1(n9429), .IN2(data_sec[45]), .IN3(n9427), .IN4(
        data_csc[45]), .Q(n9286) );
  AO22X1 U10154 ( .IN1(n4559), .IN2(data_tan[45]), .IN3(n9426), .IN4(
        data_cos[45]), .Q(n9285) );
  OR3X1 U10155 ( .IN1(n9287), .IN2(n9286), .IN3(n9285), .Q(N431) );
  AO22X1 U10156 ( .IN1(n9421), .IN2(data_cos[44]), .IN3(n9427), .IN4(
        data_csc[44]), .Q(n9290) );
  AO22X1 U10157 ( .IN1(n9429), .IN2(data_sec[44]), .IN3(n9419), .IN4(
        data_cot[44]), .Q(n9289) );
  AO22X1 U10158 ( .IN1(n4559), .IN2(data_tan[44]), .IN3(n9428), .IN4(
        data_sin[44]), .Q(n9288) );
  OR3X1 U10159 ( .IN1(n9290), .IN2(n9289), .IN3(n9288), .Q(N430) );
  AO22X1 U10160 ( .IN1(n9426), .IN2(data_cos[43]), .IN3(n9428), .IN4(
        data_sin[43]), .Q(n9293) );
  AO22X1 U10161 ( .IN1(n9429), .IN2(data_sec[43]), .IN3(n9427), .IN4(
        data_csc[43]), .Q(n9292) );
  AO22X1 U10162 ( .IN1(n4561), .IN2(data_tan[43]), .IN3(n9419), .IN4(
        data_cot[43]), .Q(n9291) );
  OR3X1 U10163 ( .IN1(n9293), .IN2(n9292), .IN3(n9291), .Q(N429) );
  AO22X1 U10164 ( .IN1(n9421), .IN2(data_cos[42]), .IN3(n9419), .IN4(
        data_cot[42]), .Q(n9296) );
  AO22X1 U10165 ( .IN1(n9429), .IN2(data_sec[42]), .IN3(n9427), .IN4(
        data_csc[42]), .Q(n9295) );
  AO22X1 U10166 ( .IN1(n4560), .IN2(data_tan[42]), .IN3(n9428), .IN4(
        data_sin[42]), .Q(n9294) );
  OR3X1 U10167 ( .IN1(n9296), .IN2(n9295), .IN3(n9294), .Q(N428) );
  AO22X1 U10168 ( .IN1(n9425), .IN2(data_cot[41]), .IN3(n9428), .IN4(
        data_sin[41]), .Q(n9299) );
  AO22X1 U10169 ( .IN1(n4561), .IN2(data_tan[41]), .IN3(n9427), .IN4(
        data_csc[41]), .Q(n9298) );
  AO22X1 U10170 ( .IN1(n9429), .IN2(data_sec[41]), .IN3(n9426), .IN4(
        data_cos[41]), .Q(n9297) );
  OR3X1 U10171 ( .IN1(n9299), .IN2(n9298), .IN3(n9297), .Q(N427) );
  AO22X1 U10172 ( .IN1(n4560), .IN2(data_tan[40]), .IN3(n9429), .IN4(
        data_sec[40]), .Q(n9302) );
  AO22X1 U10173 ( .IN1(n9425), .IN2(data_cot[40]), .IN3(n9427), .IN4(
        data_csc[40]), .Q(n9301) );
  AO22X1 U10174 ( .IN1(n9426), .IN2(data_cos[40]), .IN3(n9428), .IN4(
        data_sin[40]), .Q(n9300) );
  OR3X1 U10175 ( .IN1(n9302), .IN2(n9301), .IN3(n9300), .Q(N426) );
  AO22X1 U10176 ( .IN1(n9421), .IN2(data_cos[39]), .IN3(n9427), .IN4(
        data_csc[39]), .Q(n9306) );
  INVX0 U10177 ( .INP(n9428), .ZN(n9303) );
  INVX0 U10178 ( .INP(n9303), .ZN(n9418) );
  AO22X1 U10179 ( .IN1(n9419), .IN2(data_cot[39]), .IN3(n9418), .IN4(
        data_sin[39]), .Q(n9305) );
  AO22X1 U10180 ( .IN1(n4561), .IN2(data_tan[39]), .IN3(n9429), .IN4(
        data_sec[39]), .Q(n9304) );
  OR3X1 U10181 ( .IN1(n9306), .IN2(n9305), .IN3(n9304), .Q(N425) );
  AO22X1 U10182 ( .IN1(n9419), .IN2(data_cot[38]), .IN3(n9428), .IN4(
        data_sin[38]), .Q(n9309) );
  AO22X1 U10183 ( .IN1(n9429), .IN2(data_sec[38]), .IN3(n9420), .IN4(
        data_csc[38]), .Q(n9308) );
  AO22X1 U10184 ( .IN1(n4560), .IN2(data_tan[38]), .IN3(n9421), .IN4(
        data_cos[38]), .Q(n9307) );
  OR3X1 U10185 ( .IN1(n9309), .IN2(n9308), .IN3(n9307), .Q(N424) );
  AO22X1 U10186 ( .IN1(n9426), .IN2(data_cos[37]), .IN3(n9425), .IN4(
        data_cot[37]), .Q(n9312) );
  AO22X1 U10187 ( .IN1(n4559), .IN2(data_tan[37]), .IN3(n9420), .IN4(
        data_csc[37]), .Q(n9311) );
  AO22X1 U10188 ( .IN1(n9429), .IN2(data_sec[37]), .IN3(n9418), .IN4(
        data_sin[37]), .Q(n9310) );
  OR3X1 U10189 ( .IN1(n9312), .IN2(n9311), .IN3(n9310), .Q(N423) );
  AO22X1 U10190 ( .IN1(n9421), .IN2(data_cos[36]), .IN3(n9425), .IN4(
        data_cot[36]), .Q(n9315) );
  AO22X1 U10191 ( .IN1(n4559), .IN2(data_tan[36]), .IN3(n9427), .IN4(
        data_csc[36]), .Q(n9314) );
  AO22X1 U10192 ( .IN1(n9429), .IN2(data_sec[36]), .IN3(n9418), .IN4(
        data_sin[36]), .Q(n9313) );
  OR3X1 U10193 ( .IN1(n9315), .IN2(n9314), .IN3(n9313), .Q(N422) );
  AO22X1 U10194 ( .IN1(n9429), .IN2(data_sec[35]), .IN3(n9427), .IN4(
        data_csc[35]), .Q(n9318) );
  AO22X1 U10195 ( .IN1(n9421), .IN2(data_cos[35]), .IN3(n9418), .IN4(
        data_sin[35]), .Q(n9317) );
  AO22X1 U10196 ( .IN1(n4559), .IN2(data_tan[35]), .IN3(n9419), .IN4(
        data_cot[35]), .Q(n9316) );
  OR3X1 U10197 ( .IN1(n9318), .IN2(n9317), .IN3(n9316), .Q(N421) );
  AO22X1 U10198 ( .IN1(n9429), .IN2(data_sec[34]), .IN3(n9426), .IN4(
        data_cos[34]), .Q(n9321) );
  AO22X1 U10199 ( .IN1(n4561), .IN2(data_tan[34]), .IN3(n9420), .IN4(
        data_csc[34]), .Q(n9320) );
  AO22X1 U10200 ( .IN1(n9419), .IN2(data_cot[34]), .IN3(n9418), .IN4(
        data_sin[34]), .Q(n9319) );
  OR3X1 U10201 ( .IN1(n9321), .IN2(n9320), .IN3(n9319), .Q(N420) );
  AO22X1 U10202 ( .IN1(n9426), .IN2(data_cos[33]), .IN3(n9419), .IN4(
        data_cot[33]), .Q(n9324) );
  AO22X1 U10203 ( .IN1(n9429), .IN2(data_sec[33]), .IN3(n9427), .IN4(
        data_csc[33]), .Q(n9323) );
  AO22X1 U10204 ( .IN1(n4560), .IN2(data_tan[33]), .IN3(n9418), .IN4(
        data_sin[33]), .Q(n9322) );
  OR3X1 U10205 ( .IN1(n9324), .IN2(n9323), .IN3(n9322), .Q(N419) );
  AO22X1 U10206 ( .IN1(n9426), .IN2(data_cos[32]), .IN3(n9418), .IN4(
        data_sin[32]), .Q(n9327) );
  AO22X1 U10207 ( .IN1(n9429), .IN2(data_sec[32]), .IN3(n9420), .IN4(
        data_csc[32]), .Q(n9326) );
  AO22X1 U10208 ( .IN1(n4561), .IN2(data_tan[32]), .IN3(n9425), .IN4(
        data_cot[32]), .Q(n9325) );
  OR3X1 U10209 ( .IN1(n9327), .IN2(n9326), .IN3(n9325), .Q(N418) );
  AO22X1 U10210 ( .IN1(n9425), .IN2(data_cot[31]), .IN3(n9420), .IN4(
        data_csc[31]), .Q(n9330) );
  AO22X1 U10211 ( .IN1(n9429), .IN2(data_sec[31]), .IN3(n9421), .IN4(
        data_cos[31]), .Q(n9329) );
  AO22X1 U10212 ( .IN1(n4560), .IN2(data_tan[31]), .IN3(n9418), .IN4(
        data_sin[31]), .Q(n9328) );
  OR3X1 U10213 ( .IN1(n9330), .IN2(n9329), .IN3(n9328), .Q(N417) );
  AO22X1 U10214 ( .IN1(n9419), .IN2(data_cot[30]), .IN3(n9427), .IN4(
        data_csc[30]), .Q(n9333) );
  AO22X1 U10215 ( .IN1(n9429), .IN2(data_sec[30]), .IN3(n9426), .IN4(
        data_cos[30]), .Q(n9332) );
  AO22X1 U10216 ( .IN1(n4561), .IN2(data_tan[30]), .IN3(n9418), .IN4(
        data_sin[30]), .Q(n9331) );
  OR3X1 U10217 ( .IN1(n9333), .IN2(n9332), .IN3(n9331), .Q(N416) );
  AO22X1 U10218 ( .IN1(n9425), .IN2(data_cot[29]), .IN3(n9427), .IN4(
        data_csc[29]), .Q(n9336) );
  AO22X1 U10219 ( .IN1(n9429), .IN2(data_sec[29]), .IN3(n9421), .IN4(
        data_cos[29]), .Q(n9335) );
  AO22X1 U10220 ( .IN1(n4560), .IN2(data_tan[29]), .IN3(n9418), .IN4(
        data_sin[29]), .Q(n9334) );
  OR3X1 U10221 ( .IN1(n9336), .IN2(n9335), .IN3(n9334), .Q(N415) );
  AO22X1 U10222 ( .IN1(n9429), .IN2(data_sec[28]), .IN3(n9420), .IN4(
        data_csc[28]), .Q(n9339) );
  AO22X1 U10223 ( .IN1(n4559), .IN2(data_tan[28]), .IN3(n9426), .IN4(
        data_cos[28]), .Q(n9338) );
  AO22X1 U10224 ( .IN1(n9419), .IN2(data_cot[28]), .IN3(n9428), .IN4(
        data_sin[28]), .Q(n9337) );
  OR3X1 U10225 ( .IN1(n9339), .IN2(n9338), .IN3(n9337), .Q(N414) );
  AO22X1 U10226 ( .IN1(n9429), .IN2(data_sec[27]), .IN3(n9421), .IN4(
        data_cos[27]), .Q(n9342) );
  AO22X1 U10227 ( .IN1(n4559), .IN2(data_tan[27]), .IN3(n9420), .IN4(
        data_csc[27]), .Q(n9341) );
  AO22X1 U10228 ( .IN1(n9425), .IN2(data_cot[27]), .IN3(n9418), .IN4(
        data_sin[27]), .Q(n9340) );
  OR3X1 U10229 ( .IN1(n9342), .IN2(n9341), .IN3(n9340), .Q(N413) );
  AO22X1 U10230 ( .IN1(n4559), .IN2(data_tan[26]), .IN3(n9419), .IN4(
        data_cot[26]), .Q(n9345) );
  AO22X1 U10231 ( .IN1(n9428), .IN2(data_sin[26]), .IN3(n9427), .IN4(
        data_csc[26]), .Q(n9344) );
  AO22X1 U10232 ( .IN1(n9429), .IN2(data_sec[26]), .IN3(n9426), .IN4(
        data_cos[26]), .Q(n9343) );
  OR3X1 U10233 ( .IN1(n9345), .IN2(n9344), .IN3(n9343), .Q(N412) );
  AO22X1 U10234 ( .IN1(n9419), .IN2(data_cot[25]), .IN3(n9420), .IN4(
        data_csc[25]), .Q(n9348) );
  AO22X1 U10235 ( .IN1(n9429), .IN2(data_sec[25]), .IN3(n9421), .IN4(
        data_cos[25]), .Q(n9347) );
  AO22X1 U10236 ( .IN1(n4561), .IN2(data_tan[25]), .IN3(n9418), .IN4(
        data_sin[25]), .Q(n9346) );
  OR3X1 U10237 ( .IN1(n9348), .IN2(n9347), .IN3(n9346), .Q(N411) );
  AO22X1 U10238 ( .IN1(n4560), .IN2(data_tan[24]), .IN3(n9426), .IN4(
        data_cos[24]), .Q(n9351) );
  AO22X1 U10239 ( .IN1(n9429), .IN2(data_sec[24]), .IN3(n9427), .IN4(
        data_csc[24]), .Q(n9350) );
  AO22X1 U10240 ( .IN1(n9425), .IN2(data_cot[24]), .IN3(n9428), .IN4(
        data_sin[24]), .Q(n9349) );
  OR3X1 U10241 ( .IN1(n9351), .IN2(n9350), .IN3(n9349), .Q(N410) );
  AO22X1 U10242 ( .IN1(n9429), .IN2(data_sec[23]), .IN3(n9419), .IN4(
        data_cot[23]), .Q(n9354) );
  AO22X1 U10243 ( .IN1(n4558), .IN2(data_tan[23]), .IN3(n9420), .IN4(
        data_csc[23]), .Q(n9353) );
  AO22X1 U10244 ( .IN1(n9421), .IN2(data_cos[23]), .IN3(n9418), .IN4(
        data_sin[23]), .Q(n9352) );
  OR3X1 U10245 ( .IN1(n9354), .IN2(n9353), .IN3(n9352), .Q(N409) );
  AO22X1 U10246 ( .IN1(n4558), .IN2(data_tan[22]), .IN3(n9421), .IN4(
        data_cos[22]), .Q(n9357) );
  AO22X1 U10247 ( .IN1(n9425), .IN2(data_cot[22]), .IN3(n9427), .IN4(
        data_csc[22]), .Q(n9356) );
  AO22X1 U10248 ( .IN1(n9429), .IN2(data_sec[22]), .IN3(n9418), .IN4(
        data_sin[22]), .Q(n9355) );
  OR3X1 U10249 ( .IN1(n9357), .IN2(n9356), .IN3(n9355), .Q(N408) );
  AO22X1 U10250 ( .IN1(n9426), .IN2(data_cos[21]), .IN3(n9418), .IN4(
        data_sin[21]), .Q(n9360) );
  AO22X1 U10251 ( .IN1(n9419), .IN2(data_cot[21]), .IN3(n9427), .IN4(
        data_csc[21]), .Q(n9359) );
  AO22X1 U10252 ( .IN1(n4558), .IN2(data_tan[21]), .IN3(n9429), .IN4(
        data_sec[21]), .Q(n9358) );
  OR3X1 U10253 ( .IN1(n9360), .IN2(n9359), .IN3(n9358), .Q(N407) );
  AO22X1 U10254 ( .IN1(n9429), .IN2(data_sec[20]), .IN3(n9428), .IN4(
        data_sin[20]), .Q(n9363) );
  AO22X1 U10255 ( .IN1(n4558), .IN2(data_tan[20]), .IN3(n9420), .IN4(
        data_csc[20]), .Q(n9362) );
  AO22X1 U10256 ( .IN1(n9421), .IN2(data_cos[20]), .IN3(n9419), .IN4(
        data_cot[20]), .Q(n9361) );
  OR3X1 U10257 ( .IN1(n9363), .IN2(n9362), .IN3(n9361), .Q(N406) );
  AO22X1 U10258 ( .IN1(n9425), .IN2(data_cot[19]), .IN3(n9418), .IN4(
        data_sin[19]), .Q(n9366) );
  AO22X1 U10259 ( .IN1(n4558), .IN2(data_tan[19]), .IN3(n9420), .IN4(
        data_csc[19]), .Q(n9365) );
  AO22X1 U10260 ( .IN1(n9429), .IN2(data_sec[19]), .IN3(n9421), .IN4(
        data_cos[19]), .Q(n9364) );
  OR3X1 U10261 ( .IN1(n9366), .IN2(n9365), .IN3(n9364), .Q(N405) );
  AO22X1 U10262 ( .IN1(n9426), .IN2(data_cos[18]), .IN3(n9419), .IN4(
        data_cot[18]), .Q(n9369) );
  AO22X1 U10263 ( .IN1(n9428), .IN2(data_sin[18]), .IN3(n9427), .IN4(
        data_csc[18]), .Q(n9368) );
  AO22X1 U10264 ( .IN1(n4558), .IN2(data_tan[18]), .IN3(n9429), .IN4(
        data_sec[18]), .Q(n9367) );
  OR3X1 U10265 ( .IN1(n9369), .IN2(n9368), .IN3(n9367), .Q(N404) );
  AO22X1 U10266 ( .IN1(n4558), .IN2(data_tan[17]), .IN3(n9427), .IN4(
        data_csc[17]), .Q(n9372) );
  AO22X1 U10267 ( .IN1(n9426), .IN2(data_cos[17]), .IN3(n9425), .IN4(
        data_cot[17]), .Q(n9371) );
  AO22X1 U10268 ( .IN1(n9429), .IN2(data_sec[17]), .IN3(n9418), .IN4(
        data_sin[17]), .Q(n9370) );
  OR3X1 U10269 ( .IN1(n9372), .IN2(n9371), .IN3(n9370), .Q(N403) );
  AO22X1 U10270 ( .IN1(n9429), .IN2(data_sec[16]), .IN3(n9421), .IN4(
        data_cos[16]), .Q(n9375) );
  AO22X1 U10271 ( .IN1(n4558), .IN2(data_tan[16]), .IN3(n9420), .IN4(
        data_csc[16]), .Q(n9374) );
  AO22X1 U10272 ( .IN1(n9425), .IN2(data_cot[16]), .IN3(n9418), .IN4(
        data_sin[16]), .Q(n9373) );
  OR3X1 U10273 ( .IN1(n9375), .IN2(n9374), .IN3(n9373), .Q(N402) );
  AO22X1 U10274 ( .IN1(n9429), .IN2(data_sec[15]), .IN3(n9428), .IN4(
        data_sin[15]), .Q(n9378) );
  AO22X1 U10275 ( .IN1(n9419), .IN2(data_cot[15]), .IN3(n9420), .IN4(
        data_csc[15]), .Q(n9377) );
  AO22X1 U10276 ( .IN1(n4558), .IN2(data_tan[15]), .IN3(n9421), .IN4(
        data_cos[15]), .Q(n9376) );
  OR3X1 U10277 ( .IN1(n9378), .IN2(n9377), .IN3(n9376), .Q(N401) );
  AO22X1 U10278 ( .IN1(n4558), .IN2(data_tan[14]), .IN3(n9420), .IN4(
        data_csc[14]), .Q(n9381) );
  AO22X1 U10279 ( .IN1(n9426), .IN2(data_cos[14]), .IN3(n9418), .IN4(
        data_sin[14]), .Q(n9380) );
  AO22X1 U10280 ( .IN1(n9429), .IN2(data_sec[14]), .IN3(n9425), .IN4(
        data_cot[14]), .Q(n9379) );
  OR3X1 U10281 ( .IN1(n9381), .IN2(n9380), .IN3(n9379), .Q(N400) );
  AO22X1 U10282 ( .IN1(n9425), .IN2(data_cot[13]), .IN3(n9418), .IN4(
        data_sin[13]), .Q(n9384) );
  AO22X1 U10283 ( .IN1(n9429), .IN2(data_sec[13]), .IN3(n9420), .IN4(
        data_csc[13]), .Q(n9383) );
  AO22X1 U10284 ( .IN1(n4558), .IN2(data_tan[13]), .IN3(n9421), .IN4(
        data_cos[13]), .Q(n9382) );
  OR3X1 U10285 ( .IN1(n9384), .IN2(n9383), .IN3(n9382), .Q(N399) );
  AO22X1 U10286 ( .IN1(n4558), .IN2(data_tan[12]), .IN3(n9421), .IN4(
        data_cos[12]), .Q(n9387) );
  AO22X1 U10287 ( .IN1(n9429), .IN2(data_sec[12]), .IN3(n9420), .IN4(
        data_csc[12]), .Q(n9386) );
  AO22X1 U10288 ( .IN1(n9419), .IN2(data_cot[12]), .IN3(n9418), .IN4(
        data_sin[12]), .Q(n9385) );
  OR3X1 U10289 ( .IN1(n9387), .IN2(n9386), .IN3(n9385), .Q(N398) );
  AO22X1 U10290 ( .IN1(n9426), .IN2(data_cos[11]), .IN3(n9418), .IN4(
        data_sin[11]), .Q(n9390) );
  AO22X1 U10291 ( .IN1(n9429), .IN2(data_sec[11]), .IN3(n9420), .IN4(
        data_csc[11]), .Q(n9389) );
  AO22X1 U10292 ( .IN1(n4561), .IN2(data_tan[11]), .IN3(n9425), .IN4(
        data_cot[11]), .Q(n9388) );
  OR3X1 U10293 ( .IN1(n9390), .IN2(n9389), .IN3(n9388), .Q(N397) );
  AO22X1 U10294 ( .IN1(n9426), .IN2(data_cos[10]), .IN3(n9425), .IN4(
        data_cot[10]), .Q(n9393) );
  AO22X1 U10295 ( .IN1(n4560), .IN2(data_tan[10]), .IN3(n9420), .IN4(
        data_csc[10]), .Q(n9392) );
  AO22X1 U10296 ( .IN1(n9429), .IN2(data_sec[10]), .IN3(n9418), .IN4(
        data_sin[10]), .Q(n9391) );
  OR3X1 U10297 ( .IN1(n9393), .IN2(n9392), .IN3(n9391), .Q(N396) );
  AO22X1 U10298 ( .IN1(n9429), .IN2(data_sec[9]), .IN3(n9420), .IN4(
        data_csc[9]), .Q(n9396) );
  AO22X1 U10299 ( .IN1(n9426), .IN2(data_cos[9]), .IN3(n9425), .IN4(
        data_cot[9]), .Q(n9395) );
  AO22X1 U10300 ( .IN1(n4561), .IN2(data_tan[9]), .IN3(n9418), .IN4(
        data_sin[9]), .Q(n9394) );
  OR3X1 U10301 ( .IN1(n9396), .IN2(n9395), .IN3(n9394), .Q(N395) );
  AO22X1 U10302 ( .IN1(n4559), .IN2(data_tan[8]), .IN3(n9421), .IN4(
        data_cos[8]), .Q(n9399) );
  AO22X1 U10303 ( .IN1(n9425), .IN2(data_cot[8]), .IN3(n9420), .IN4(
        data_csc[8]), .Q(n9398) );
  AO22X1 U10304 ( .IN1(n9429), .IN2(data_sec[8]), .IN3(n9418), .IN4(
        data_sin[8]), .Q(n9397) );
  OR3X1 U10305 ( .IN1(n9399), .IN2(n9398), .IN3(n9397), .Q(N394) );
  AO22X1 U10306 ( .IN1(n9419), .IN2(data_cot[7]), .IN3(n9420), .IN4(
        data_csc[7]), .Q(n9402) );
  AO22X1 U10307 ( .IN1(n9426), .IN2(data_cos[7]), .IN3(n9418), .IN4(
        data_sin[7]), .Q(n9401) );
  AO22X1 U10308 ( .IN1(n4559), .IN2(data_tan[7]), .IN3(n9429), .IN4(
        data_sec[7]), .Q(n9400) );
  OR3X1 U10309 ( .IN1(n9402), .IN2(n9401), .IN3(n9400), .Q(N393) );
  AO22X1 U10310 ( .IN1(n9429), .IN2(data_sec[6]), .IN3(n9421), .IN4(
        data_cos[6]), .Q(n9405) );
  AO22X1 U10311 ( .IN1(n9425), .IN2(data_cot[6]), .IN3(n9427), .IN4(
        data_csc[6]), .Q(n9404) );
  AO22X1 U10312 ( .IN1(n4560), .IN2(data_tan[6]), .IN3(n9418), .IN4(
        data_sin[6]), .Q(n9403) );
  OR3X1 U10313 ( .IN1(n9405), .IN2(n9404), .IN3(n9403), .Q(N392) );
  AO22X1 U10314 ( .IN1(n4560), .IN2(data_tan[5]), .IN3(n9429), .IN4(
        data_sec[5]), .Q(n9408) );
  AO22X1 U10315 ( .IN1(n9419), .IN2(data_cot[5]), .IN3(n9427), .IN4(
        data_csc[5]), .Q(n9407) );
  AO22X1 U10316 ( .IN1(n9426), .IN2(data_cos[5]), .IN3(n9418), .IN4(
        data_sin[5]), .Q(n9406) );
  OR3X1 U10317 ( .IN1(n9408), .IN2(n9407), .IN3(n9406), .Q(N391) );
  AO22X1 U10318 ( .IN1(n9429), .IN2(data_sec[4]), .IN3(n9420), .IN4(
        data_csc[4]), .Q(n9411) );
  AO22X1 U10319 ( .IN1(n4561), .IN2(data_tan[4]), .IN3(n9421), .IN4(
        data_cos[4]), .Q(n9410) );
  AO22X1 U10320 ( .IN1(n9425), .IN2(data_cot[4]), .IN3(n9418), .IN4(
        data_sin[4]), .Q(n9409) );
  OR3X1 U10321 ( .IN1(n9411), .IN2(n9410), .IN3(n9409), .Q(N390) );
  AO22X1 U10322 ( .IN1(n9429), .IN2(data_sec[3]), .IN3(n9421), .IN4(
        data_cos[3]), .Q(n9414) );
  AO22X1 U10323 ( .IN1(n9419), .IN2(data_cot[3]), .IN3(n9420), .IN4(
        data_csc[3]), .Q(n9413) );
  AO22X1 U10324 ( .IN1(n4559), .IN2(data_tan[3]), .IN3(n9418), .IN4(
        data_sin[3]), .Q(n9412) );
  OR3X1 U10325 ( .IN1(n9414), .IN2(n9413), .IN3(n9412), .Q(N389) );
  AO22X1 U10326 ( .IN1(n9429), .IN2(data_sec[2]), .IN3(n9421), .IN4(
        data_cos[2]), .Q(n9417) );
  AO22X1 U10327 ( .IN1(n9425), .IN2(data_cot[2]), .IN3(n9420), .IN4(
        data_csc[2]), .Q(n9416) );
  AO22X1 U10328 ( .IN1(n4561), .IN2(data_tan[2]), .IN3(n9418), .IN4(
        data_sin[2]), .Q(n9415) );
  OR3X1 U10329 ( .IN1(n9417), .IN2(n9416), .IN3(n9415), .Q(N388) );
  AO22X1 U10330 ( .IN1(n9419), .IN2(data_cot[1]), .IN3(n9418), .IN4(
        data_sin[1]), .Q(n9424) );
  AO22X1 U10331 ( .IN1(n9429), .IN2(data_sec[1]), .IN3(n9420), .IN4(
        data_csc[1]), .Q(n9423) );
  AO22X1 U10332 ( .IN1(n4560), .IN2(data_tan[1]), .IN3(n9421), .IN4(
        data_cos[1]), .Q(n9422) );
  OR3X1 U10333 ( .IN1(n9424), .IN2(n9423), .IN3(n9422), .Q(N387) );
  AO22X1 U10334 ( .IN1(n9426), .IN2(data_cos[0]), .IN3(n9425), .IN4(
        data_cot[0]), .Q(n9432) );
  AO22X1 U10335 ( .IN1(n9428), .IN2(data_sin[0]), .IN3(n9427), .IN4(
        data_csc[0]), .Q(n9431) );
  AO22X1 U10336 ( .IN1(n4558), .IN2(data_tan[0]), .IN3(n9429), .IN4(
        data_sec[0]), .Q(n9430) );
  OR3X1 U10337 ( .IN1(n9432), .IN2(n9431), .IN3(n9430), .Q(N386) );
endmodule

